// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FoSIlx5jZhFipTAXw6vMVOScXArP2NI+yndFRHVdnKwFYj4q6ofDcocelUAtdbwU
krXpSzwkI7+H6YRfQptPSgvBZ8nsaxgOXcgytCIZA72CHRdxMeB0m32ArfukUCcq
swDRqdTNKfurw8dLo5re872rzgD6O5HrxkwRJZvbEt0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20368)
PC8jIxgnj3mK/NG/LY1xQZgomOUILqm30vu3fDIX3Ry3KHyhprO/U8rK0aV7k1Rh
Y8ARfglXhIg1XxVWZR4KqC2nIoBlek00Ny4uV04sRGfMsgDSzpRbqjZ9pBwRcz2z
ycnStM3P31lIXQIE4v7YpQFAaxYNYUWI71z3ZqRECxrlzuVZRjGoftla6vO3MEWX
wui1k/dsX2no3LQETTh8p0H2k3Rd9sgX2lUdkjk34ySTncRwvnpjJrvaHrLgPGf2
vZyD2ov64gZP8Or31G4LbvFL+Vlz6XR41eEfb3oqUwkwp6eD8+x/RYivRzXZz0/y
KqpB24Qerb2H/S6g+ZBbPl5EfTeN2aFgEeDz+ARabGmb39XnCARE/vM0RUuIRAug
jRJu6u8F/lUR09xdOrq0XLvwLGmQV5b6Ic+HoHuT6lhRu/RX/O46jojkX5Z2+fqG
5sF4C6LPY7zrXEOWrrotnhR5ZiJsyjYCNaIEEcxZB03hcMu//mqLGAkEOGxyVXz0
fIyMJass8VgOGY8zcUNdhMrJqq6JF2VQUMrtYeZeFHYQ62UPCOaUN7lJR2kuCnDs
90VUW2tMyBDYjXqbuVMX9N+9qD4PNmZXrOXJ+HakT/imcg7ytDHLkSwIL5R59Lfp
GLYX5FgWYDshSqglip2Nv5ZqnhO2nNJcg2IID4qI2QtMRzz/WH3ob6ZtFvNcj4xC
pOBnEli35WcYfRLNidY0R2i9KiOIWfNZDfXY5Kve+heEFOcGCBTVRj4AxU+JqPy2
UAyoTfWRTvEn175QUn4EJapbdvI9q95RWaOCGTcTWgT+TOMpUJw/mDBANzRyTk+Z
fl1saPbG540DCkM4cP3Qy3qmWGX+2WDUbRtaIvh6TB1uhESH8MprhG1Hd/P7gwgb
M7aHAXQvnpOUd5hIiGS+O7AD75UHoLhSfW4m972Sbx/R9p5et5RvuMpEzIg8frOH
4SwydHcrPLVgBX2uRBQ+EnobfMaMIJbUS4fsimMO6alkZ07cWfyTG8D62QTmErpN
UGATnhJi4LAgKKniLpO1TcM5uV5A+WbRTpT3SgkELTqYio3W2fgScEueivkHK4Ha
b76jOgPMhNiKRHDGgIysy73jPJ21Ob+LFyJ3BASwqOeVpyfuwj25rPBCKGIgVIx2
EVyDHc8B0TKZ4nBWKhFn238ujKDs1RN3cmrVtopnjm/E0wCy/1KMzSvl9IhHIA1z
M1Hi0EV+ciOwbt+wiYTw8vV3ZA1OElZDb/920qZFFjWoyAoRFGIlvrqKuLAqU54Q
rybfB8zQ3nS8GYn3LcoEI7tEzTlF3/l8sGLR/8dzugHFfvTchXXpA6HYeKKhbA2O
JXEeJgL/5z6IrusDTQN2iahd0lv7TB5UvOXa+1nro9jlZh8kX3i/bnuvoX5yro+N
Kg9Yzw+9iv2iDwpvZu9hvrVIX/VK0dzv03IRhWbIsI+mQv4J8HoTdvHnafcxa5oo
eq/46wJI8mZYgFDXDQKrHWqHzJ8R2pcvWLdEvFLTpfTF8bDznwBhvub9Pg9COnkD
eOmQhBDNWhYmj10HO6/RUqS8MfAbEILvETlAo7qmkJsw7G7XNaAStsY2DCD9TsJ4
uc8dqfLtaNqwngaBXrZLA8rQhfGZiqgvqsZkrwvVy9itppjiKb2nMlNcHbU1zJvy
KczgRzLC06KwJU5cn/XY019otPrenUcupatXMI8VvdwHMfdSCxRYNvW/2pk6AGkk
Lq8rZfdhH3UYHq/ISdDVoF4AhmuC4beY109psYqVf742QdFjmb2AbcapO/GVxVuw
SawwJUyc2pbA5rHdh+KMUdYr/xiFcDIoeXpEA14RyyvevcDlav/QqWhQ7dlgIZXW
eOOsfMQX56mmzOH2m7qUc6jWyb7jqpgJ7bU1+3Qvb+87sN3WqQSunSTkizJ0qfgN
Xp08Z3/t+IZU/1Stl9AZh/3+5Jin3R81N2oDeDaCe3GBe9dQnDjOJyXdmxmpT7R6
R5NaZgLO05ZbOk3+jFtcBcpGaZ/qQZxI1BLoE1w3diPedBAXWzCasuYoNm//byj/
pMnsQHIHAUOtzy1EucUzSBgKblW5caDzeJrhKcT4QzKOOz1uV9mmNLTQB9XjwcYy
iLCXv2OWntR2olDtVMgFuWdzNuDnlWwljwH6+GDcYymnSBWsXHj0eaSwps6vCpmQ
HCYKiS7CNm2qUR3isvkAovlEE+O9IX49GIwgPtffk/cAMKlUeNVmJ36RAf8/eRgL
jM3D5PQS65eIB8bMo3cZOMU/b2EA2emtaPJVUdAZrUOp+uEm1BUE0IAtffHwEfLy
okz6iKPfqU/MVD+PFaIq5l5t7qaHpcrfyykfdJGeeVNtqP17nOvQpsNMDXSp26sE
Puv0lrIb6hf3Z3uVzxe9gxvXlvc9FTuVJIOQy8JmYpmuZCXKrNpa4zUTQD3ivYWB
HXyNV74UbaZoM/35hxyh09GqYdX17R5PC3Bd0BYNe+Kb3oRVbujvVj8FSG8hJC+A
qnJ2IvGs7xP2znj8lCMCrA73+ZOO+vt8NTAJ2uOa6JDRl3Nw4hPfDiBkd68OdZre
sDU6+k+yltQ5sqYHyJdUpkeucw9I6dvU/9zMLH2CCgALD8+gkPqkPIpEK1cY2ejt
hS8YKrsNf+rPS1+laVI28I9K0rigJfBBmQfEVW79nqQdKFGOg5TCxBp1r/nuOKYF
yZQ5WP1YrQxOe6OFa9s5fbNZX4S6m7gVy1Axec37w5vCAPHc1kDa7Mu3k7ilkZIX
2J/Ziyv6HaNlOvtBNkDaZCiMNeFmcN0GBDudYiH9hmqMC0e+57kLXhVlM5VwpyVu
d5o2rBZySmWAvJZjdpQ/pCrZH7ZcqTr+XH1orxpil6J1NYNPEV9SIhEX1y2JPfwL
Ki2CURrzvFOdFB6M1vE3gWpEmT1uzYvLzxbPX630ui2gl4Q6MixPrFrh/zoHAylT
JoZcfjWzacVVvQxtfG1DZEZ3y27A462dFNw3qbaYXu2YIjbIYaf/Qn0Hb2O2nHZ1
uA9OK10wdtZlj4pcDbrWQnrdHBnR71wQZ1RPm/nAbBXU1Qmc5jNKnUsjTDYn8Mx0
fA83UHOKYRqusZUFy4JQI6IKBKEkoDBEq3/GE/NQSWk/xv3SMgs5K58xyBWgpjiu
Rt7HTNufCD5Feoa4XWvkzbB/OViXfRPPfn/WdQmaHrNUq2QUPu5axFFMOgn0OmFV
UxmrgCJe5egQ2p/dlppPHrOmF8TymssPAqLPjoLUlG4a57xH0qBFOEBn9oBYBQ//
kdaAppUImXz1KX20Rvg/loH2lRfB2J4zbuqR6HNCUU0t7Jr0H/FfIBsehHvzeHZJ
F3dL0G2qgr1Bti759vfTJliGWZfkQS//G7OtpKId0dXbd5Ch13KZx/TLDQNB1UfW
eclP/DwOx9acj/crxX/ibYitB4BY9Hq6bC/j8F+ueA71TRVnrUY+6FTJ2KlPfwsv
B13Hbp0hYsK190x0d6ldAZzW1tIABC6WYtl2j8OdOZnJTixjicIR8mp7s8coN14C
vYkazszUA3KWtCFmPKGay+CNBgbBM1/H7rkoA0i7lpCNrqHkhYXrOg/lq0/Rf0j2
bzvdqDd0q/LVsGjMgieeMZEoShj0Ttnt8XhcVxMFKefQMjJX2M0U1udfMndkq3xw
AAkz6IeDvo9lh2f/ZECctzQoRvRzgzvdgBAWMz7TYh/sY71PHdLctFCZ/34p9lnF
MrBh6oFV1qthx6xCLFblmEvtm5IFBUEbw0A3D6+4KAjHuGHRQtOfTCJI52y4Ymv3
wQkL5KVR5Bez864CP/ReaRt3Ajz+gJp7TgRf1tH2Rm+E3G6JJ9xQWbNFJkG7TWZb
+DkTTkSs/6RLhChG/kmat5KBDpXS5r52JQAEh7MeeiItbyDITdt2+HxIdPFc+RFW
zhO+G8ypfw6aVWm2Ga2zHv/ka+jNml69S8xc4SjYylktV/KvHvNfCtLxMeFSNDLQ
lVOhVidZWrPe3JGzGHQVtFCesO23RdBV6CLwDeuFE1Rl43M7S/Ymfe1zu1KbmKLu
FX6Ll5poKJy31UPDhoCbud+G/tKg8X3CdfteI5zgGTsTDDYIyYt80/PdGgrGWGDK
BsbuVW17VAW1DNzxTF2rWVv/o36bKpT+BVhEGOWB44n8/D3g6bSKdaM1wzPBa5Wk
czlnrEwsryrpLj2XNeSJkZvYyO9+vrSd6r0qqBOCvJ/B3YN11cvDpYgwK1aBTZsN
YH8DrOiQATGa891Ej4nTgvVhMvc9n0fWM10i/NeDgfZx7yO+1zuqwpGJwEYvSYk/
uBle/DDN/K8X7HAC7xRowhf+wvj+nQeFaHg9sXkShHoeaEWctvrMM2v2YryG3W/M
yIGErsIH/MgED9YXM+/XmH8DIu0qMRO8o+eCTylqmhtNwEqLhZV1+KBwAch25KF5
sVa9t6l7GegrN0iROneTGwE4/Pa30kIeUAFD+lVsKPdCRwqmcMezNydIXlQTQDOq
szcII+I1Red7BqH6MmYvDnkv4itu5e5jz7VEvB1H+qtySBu+6wIS1OrzWm+NwWml
uw39AtpgKMg00kEKjqS4qp3i163M0FPcYKwFPW2/QMJSrDIYfc7bLDPHcgLpaC1t
Y6Dwu/9qX+seqNZo6LovQaJ/XyuST5CM4UGjioDQ7+hfMGgPW6OvfPw1P81j1WWq
OmtFjN+yoxSKTAJaIIZ54sQNid93sgrrFJ/VSD/P7lVbFDShSvrROOzc+mR1Xbhw
UiOnZ3JPg8TJS4JGVIgtHR4o3GIQGnAjAhduqtMon5LHtCf3kfXcVRP0rOotYnr1
NcvqWJkspZc6TR971kgpYSEIYrG+3ewOvIvLJDA6HRJ+CSINatMT5FSUSFvljkka
aWJArgIRk7+NK9xVu/uTWCJ/IGSaV6H5hwN6TceKTX1SprKK6epOI50Fuky564pY
+L36TkMJbX9C27IvvIv8sUxry3uQ/+8ga55e/oP4gb7tfOJfruOP23ICWgH6cv+W
kkrxE49GcepctqlbX+vskGSwQGnqqfaGF5CtgUvE4NWt1BN/IeVstCVO7D7LaskA
n4gebdTs4Pi3qF1sSOYbOko3MBin1Dl2qrswlNeWka5/pgstwPnXut2iyQvz1Mss
LutpeMI/qsdkMHF8zOCVm8xptblbZpEEfowxiB/MNAE3BPsQyg8wgQ4IAcUQIXGk
vYXOK1RqMtIurYhjMT5dFJd8uq9JzSLm+bAQsqBepcQ8RndVEB+H0kgCwNPHFb33
9CUoTgGbuA9h6VtnYE8D5zHKOzwDAxKO7wLs3Ihnt/96qW1eiQayOEv4UqtQbzmj
4pRV3lp8SeZLpwu7uIGaF6qcmEWVdMMdaTUPfyX0pte2pFEigQOMwRV8xbWv/TeS
OfKnogtCvJUY9qzhNRoso6gTcdm1lzcEawsmtie/K17V+i0yWP+HbFznVgRUNMoM
WCF8V7ZbtK1knyu+iMrBw/L5BqIsaiN0sBeeKaYcLae/sc8xyHrUFGB3+kzfvz+n
aHg0CTy2qGVDAIDHk+EeRrLY/9scFjj+pxJeg/ZZ6nzKkYvNkuN3AQBxJBQMrL2g
cktTkPjSrqJI+9meakmf2qqkNvqTEq0SOO7Fn8QDPosh2031kLZpHXDPqHMgSG5A
fcrgNviDkLEizmiKuhu5xKQs/b1IOj2Jf8NBG1HG8mRTuAW+4SSuttsS87u3pIeJ
xh96VKd689l+TEFBUmqhi3fFaj3vI/sVHAuZPUZ1JuNQB4SHk0XFhpicaAWzWlsd
60einKoX0rljMV1iRfu0jsdVR/Kjs93nMwcEwKjwSavQU97WfQObVC4XKfbxj7s7
7UjGI5CwqZt89cAZNMy1oFNlQK77KJoGohkmlMS0sNWz3ybRma74p+KJR7pun3/f
+KCFFaX4flV4Dj/e4XSc2ynAOO0QFRJAxpcK3jLtJMGcfmU0hWz1/4ynScK0+TD/
0/unBPf39KbtzE6hRjN/Vv8qPVPkRftjAp+ZQtU3RxeiDts4qeEWJdignTjgNZeS
X0QYFU6z7MpSXVG+ZC13QT23hBa//SmGKI4Iwz35M4gmbOowThqN8JjuyMu96EiT
aSJpZAANsgLcsHgqQJqmdGs2xaWhecngYac4/bUtcZKWrhTSMEJogZOj56FnUeHB
PwB8X5TQPIxPFWoZxIraW4iSGBzLbNhvf4WLPD8diosIm/rLYGoQbnDsEe2rPz19
ALX4wUMx3/fULYLGjxIhziyT/vPDQF5BemNoEByjfG53oA7Dhw9ZdoMcdJuzqS4m
on6o55FEBVDTLEGL10WBbJH5A3z1ANgFO+8r/pINV1pbAmSzS/G+IN7NQ9afb7U1
i5e3sxxUtbpTKN/36whygW5O4wCt16RKAM0Nyb5IsJKF0zJ+3/9yo0B2bI9LG/gr
YQrUCHSGkSPBMDm6ABM3pO2KdzD9fwvmhX56Lskf5TrxmkEewyODca7xdaUrCAsa
M48NjermhQtMZAcsr0X8ROJw6l898L95D0KKmg2s0rtauRJF0IrjVBdH5zjE+MlX
uzVV9ZwxCGDahP4EVsrmsbnDHwGqhQ2dvROQgu/Os036XZIsI6nmGWN2OWvvF2nV
Ah6oI1SsfIi91bRyYNbZxsXor9F+LtCYWhWKtMsCezpJksFZgLXkgEzTSIv2jSX8
VcDepfRfxZGqkRFCvKkcGCKhEMQj8pdZi9MhOWlHnYM1zjR5QNBoNXOPoAn8Qnmz
N5Xi4eJ70iLOoOwrf+9Evd7yAMVjcpZC6037mD6mGjX5EAhpZf0dwmVbLUBNoHXm
wxx0TY7YPwOolh6udYIsc2aQqXNGm/TZ3VNwhl8n8apBEysHjma16YQqBNFncHFM
BbX9dKnbfAxMdcHQljCd0vqzJ3HMQIVPPLN7QP7dTkzZxwpFRBvPxCK305yQ3nL4
VrWEE4QgPdMIohUXI9yxG17rN0ONtlstYNd/d4yj55mYva2GrrPECki5Sr40YFj5
tbetR0RIQm+wxfN1F29YzvAUe8z45r3LGIUgk/mfbXKKTVWN8Dj6GiCE5Ynwhxpm
SopczuCbNwJClb/ZWLBc6HRC4xDOm8gWUylhB60zsoADgfcvSTELguRZnLqVOFkF
IH8ycx8K9vt1SJHNWBrU+iSGM1fwEqk9n34+0lgGHBn7A5cW4UHFoTWv8WfI9bF0
oujC+Wwg6jGqZQaHnzogHINbbKWNOSu87hQALTos3M4fnefHrptoLPc1M46+1Zw+
aorTeI1ZT9p0CwcvqUEj6IEmfRvdy4rNJBoJnpe/xjHi+Zn/OwT/HYXi+e+shRd6
jzMbsrtETXuqh+Yhd20/aflh7dzyQP1abQiu/snC0pp0dpeGMIlgXJHizjqetydl
/4Y1Ok7pxFVwojp8nEjtUly+0ujqTVZjyrsmdYpDutvSdve0/+IFROVa5GI45S6T
+bdr7wq461qjnWhHaAb0FSdc4ZfJ7wVSwqXzPqOttV2xWiXwYdgpiH5N9ZmU2Me5
VC7fZ3ciJDV5Epmcd/T09xnIpZ0pvrcaulgHmfrcKv7gPOz3sAJvlBOZ3fhbSP++
2bJgUrSER/B6j0TFCFDhEWHcZrKCOBx0ozA6yyqkB6LimZFOd6s4NKH7XP3IJOQd
G52wo0VhBXgT4CW9wqa0vf0zd9Y5wJ2ASbHl/zcxGWNgIpXlQB7PVjVErOjD5ZyN
iUap9PRb680PSBIdOtojUSuuQ+iPpy0oaT1KM14WhjvzsYZb1aP8wwnoCgFNpFee
VeLf6TFolg4aHAcRYyCSjk6/h6HmPKosBarXmCkbXCiy2JhatBSlbjIJHH/dgW/o
/STEdfbXEhWWE4wdTm7XV+5/ciu3DfkGIcb9yo7zgQ92KJiREz6nDrGNt+B43ajj
QDqBo6qJeSFQ1ANYrnX8pmKKGmzQnEjlPn/gVvaeKajo0871SZhC7eXiBLiT+KeO
X5uPMgpNM6yUibK89b+sveu0aRQdSRl0xLa2SV4zUD/aRAKZI7/WXFZCw1OxSasH
OP1lQ8ffKqBI2/911VEMjQ4yxHee3/5moq5J4kGPhD2XNEYqDi51dmZmJIDs+GSF
jG8eoP1GhUwQJM5bS10x53ytEX/oi0zLGw4LXP1eA4hCiZtzr0azUO7/t1jyzigt
SaIAfL4/XZSyeVdiCjzQJWt94R/zHuTRy0xbOoq9mZKZpgWGuD/NvSAZYmwhf7NQ
eptQpNW4ssOYRHFDw348mH+WXXlEuEo/PTKiknB3b4RVnXsYnuswxIQPeRJ57d77
V4XK4OYe14Sc1GdWdeV24HdxF065UrzaZ+xSab3BkoUUnpqd0Vk3bXiSjLdHSxQc
tKPL5huQ6y2Yh/uR3tNX2fhFvsmxpGCS5XvoRZ5U5k20+K54eYOq4fw9V/cNAeYL
X9R/xMYsNPhzI8Le9NBON8ECemN4Xu5ogFSYVUE2LYvDSjJmz5lAcSrXh1FF9LIL
3YiHqJD7YCOTfCCif1uTJVsELcZhVzm8gGtfxAWkQOXTa9rahU7FE31eYRIoGm9n
t/W3jtqmHf4DJ+qnT3kj+1hKizu6w8p+Z2mCtnSknPQHEP61PefopQq8A2335okz
OgQAREBSZktxNp93+QgLFsD/VS1Z4jc/Upv4drJeTCN0DldH/9I6on5nMWlhx3ya
DnFp1mxarlnywE2MDi0QZNEv0eUfwrCjDn03cbYTgaS3GsofeGd7JEf5pFZ/l3el
vfz4UH3VX912cr2p9kuMcPMGS9rgMNzyIbKl3Iw7xd1gi/h/qu+vXPVKJCEES1wa
Hggvrpg8JZiBfBURMJGJSOrU9DsKGCh1PdnnYZGhyJmX6cXWqCBx/M9xFug8QGKL
pC3SWE+07OOa2Cpf5lWPtZrE/x1eig+TB3aLHx0UFpf2/czt26bqKY5WmY0oMSFS
edj2OPCgDxuPToZwfsQYSWglhyvToTarT1JbsfV+3ZZRpdz0eDp/Jy40oMicEk/b
Ieyp3lGl+6T6YVfkrXH4sKIhplC1Z084c6hbNOQ/CRq66cv379hGNuk3Mo3uN8JM
jD+lLN4OiJz7iSokjnLmZrs7iVIwk2CN0WrGtHxWysCD/fSpQCKIJHkQIPdSJ9Rf
qu20DLg1umzNvJEzKQe34FnmhtuLervi16tagRZC8d4xPukIww9wzlYCr6urXvG6
pdTuXmlOR5UW2R8lW9hFvbOkv3OFV3PQWKWq65nrxiT8wo6m7+UP5PHtHM+pGx1C
ll3qk00be024vOPzSFOow5d538uDxQi8HUJ2uymCvRIxsfNC7ZkK1yMUgw/YYjIq
FUEomptharWvfK/Fevpz/XjNc/1t/b7I2KxyBYT/kBQbT1okPz7oFgCkuQR9KoP4
3ycyNRgStwsgT8PnJW3cNqTQ1PjG+gi3Vcbejc5JfdYNCE3JZ3pbZaXNnZdosqMf
zIH+WnBcvY0VbpZqP8q8jndLLn3f71ZdLDk+TyOWORW0oUOFLAhhnweteEBaAesq
dLbbXLqWuFUIVAJdFEtTjYZJDv5DuP++0ZBYHUaA7jOMqtBQ+0mHG49Qq8AEI4ck
hX5dN6aYmAidZmv1SyKGfz3wNgXMuF0sJEPjbcKRzg4X4mTqa4a3UXEZnb/vVKre
Bg7i8RGi1YuDU8A9DvvtLTw0i72tGSzEB8/JNRnuY4Tyz3UxiFLKMJict59uThhu
/PKggXPb1gfGNu8XdVv/PdGXeW/nKFgGszjlAE7+TGY/D7Nx/U54CiL7Ro2Re8zC
U0cfdTI8dZpIH/hoUnAs5ctURtlWtcu2j69PB0/CGRQXNfT1nfFgIO9AoOhAidji
LHs4Cm4IeYtx55lgVYnxu7nk0MaHshXPg20qsBGZLEnea8REs0D50Mwe1V7eGQrC
4Fi1P4b3VmsqLYaAI2cAZX4AG8ORB9QEh9Q765V+cd6W0zPStg5tiW2JKh7flsCo
+jOQdJE75PKGESlDXjcdOHnKbtLEBd13R86jtB3VyAS5pTLeweie52ohu/RrVJZM
hHwu2+YvAN+DYFAR0W+Ia7M1BUMqhis3B6bOuSTR5PsXTar0Xwvslfv5GBw5wOuQ
8FEXmY6/LuXtCmYsO8NYnpWrKj1B6v0yAhcfEVlaJzlG+IWD0R6YPNia9HPX2oXc
zaFoPOvtoTS3uCSxAba0XbVYAULtIoNBuaXXDzcG1bfyfOzv/miiaw9cgpOop3Oe
FLjTh88lW0jDvrzMHx1EFi3WZJGdpzBeB889kADbvzv8zlUDuUoG1UhXh+C0xWJD
7WZMO01eWd7tozrHb51ic3jDsq6PszSMPxUpC92K0m6Iry6sW05k5NWEyZlyhb3a
kIijBQtpmT/WC6moj0/KJhsjMSnDBMjWthg8aGXf/F7kBPKX9Ikh0cVsVqz5om1B
bP5yDYmSVRH026hucm8Ydf40DGj9NF8n1A8KAX51Tgf9QPtKJo2dnu9jSznGj2K4
EfhhpnR42xr2XqDADWPjtDTODpUKgSU7sCKLFBMnazqlS0tTN+GGLrMtqHzYOw3i
ars6rsvLs8j7/vL+w3pUYfUaNf+c5zMH9lHYOK2D/alJ1xb8ELqHJ6og9XPS6MQG
M8lw6TMhqaePtRzIVz5/pXGieMKAAmvPP36GdBwL2XRhgvcSAj6Qx5AggwuPTVa+
skHGsvWgBMZeNqlKb1IB9yGeJgy/Cpq7A6i+K6J1FF6yMy/5RFZ1THyzVplYif+N
VbE3lVQsapA0i9bvo2yaeK7PaQXXM+8Sh9d2jraaJJ5I7GidpVfZjp0NHjVViJnS
cF7ET8DCK+c0mQn4MY1tFB9Xc57O+LYIfghaChWa2hzcRNI/8DjlR6H5zwHclTdq
4NjUdxGeqMNX7OhzHJ1U5OBiS/AzQ3sAEzICqtdIutcLZXur1NfTmSr7fLL3P/58
DeJ1mXAupkMXV5UOFmVTnfTOut0LR09lJGNC7eWZU+gHXvv4SITZa+c33ohYlecM
6SiiE8SzjujeYCAY4AAQWyPsdHj43wENb3cRjm1sLV9OanDEZAFwox4j6NpTsi4E
qWH6fLHqyl15fJwUaJgnohbSzEjH9Mb9jL2nJJP9TgmvaV/57d+/3xE5Uy2RVx8S
DuDCcfec+UXtDtIp4wxGYNu6C2YWS0LYymvDeKWcaqQqEzdsJaK02b7MsxQ8Kw+f
da+q87O3nr6wiY1lzB1mODDdeVeX5Wh+GclZVG/WxGwd4ip6ApqctwjnMguGALNz
WheamwfVePimkslkS4qgmUh5rbuqtpu9TcIJ9TnM9zerMeJsXeCUw/px9LH1gA9K
ZIp7urWxVL9jlo6esPy9oMOcozBmpOy6Nm6Saz+LZu+HWX2wHJntEO2/o/prG/aN
E37U4BZC7iUAaHdE0rKy4S1Q6BvfIhNEcbXXvaQESMCDx9FrBqvYIfsr3naw3BaS
bpvLFQzo2+p4RVLrxBZaXdmulRv4XHBT/zfHW+ESFGMr4TIlA6ihKVprpEeUKqds
zXroaMdv1pjYwqBRDH6BxmS/dF9HulPEMmOyC9QJ4IDQnGMC6mp2CagB6kQzbGyG
aiZUfuoM1zfVYnsrnJEgOSRXb7DrGRYUAM4l2Fn1+Px05gtbXx1/IW0YdPuC8Kbz
41BJ1TpQwhWYgmTgwP3y8KUWRwEnwoAVAzslD4LEPnlqv2Dl6WjqjRa4qlYk6QJ3
mpwMnm1D5EXRgikOht8Xj3dza/FJ2iLvYg5PhL/6wJyX+tnFYpb17uuX0rNGE3Er
jI9H+JV58TF/2OqKx4FPoFVI7P8Ug5jXEi3gfsWFACKD8H7i0AoPoMDYsR6JItSw
r8CriZqkDdZOMYg42jjbnOfsK973sSqW33fRg9f7HnVq0Ot6WJJwT6FFtEoX3mtH
Sh/aMZOumz8puL2KZg5qIyF2UkCLFE0xHljL5brGpwUJ6NiDy6PsgLZZAmSlw2cZ
BmWsORKxIAXQYRVE8aMiOmIFH8yXcMCo80zKMCmBYp2Ln5OuzEEBvS5IDZsUiS6D
y+jSRr+GTHNkeOEcP7BGaJJcU8UexjiVpUN2tY7r2M4uxi0FG3GAljZslsHHMGKa
zrUkzViZ2nwa33johDRKUisyQvnaBtQcwUZYLhzI/5gNCBS4DiuSXw9KOlurSmPI
5e8rJp8UUkeg/SkyG8pJdH3ZJ49irSVs7oVJOCjiu5WR6USaM/lH+hxgslp3lH2Y
7uUCJLBA4kIFFa0Q5cn1EBY6mLO+SGLSHEwq49STrMCP123iyLmE4W8dkdLJjZFp
QxllwzE1lPKC3LcxhF72k8iaordXsLkSoFZJ6xe2tT6rphDUtHIQEwwvRLWwVp+P
lcuzzGyO+MapdSR8p/ZP/kV80J2Xos9vQRs1dYhP24xUuhQW0Vh4sB8TUvBwC1mG
YJa0m0IvMkSnYdyaYEe3cDVqloBrTgg2J3mA8PvTgJgw3j4twhkCxPQWz7s6NUOQ
QzDnWJHqMtMhy9VdhezTM/wjzvQHB+xiaRQtJg5q/Lsn+l4IpyryxJ/k1fUY5Ik0
sftxxy1gsw+TBuZYgnFAiU0TAFxYLw+VfXe6dJ041R+F08NynRwN7ppgjrxoQP2A
LcnxRxP+3HZvIQK/tpe90PaJnwHTHFMw2YbM8Ar9J7dcpMlB2ghyPn7eh16Sp7nM
FzRdwADQnvwqDvWtSljJe0VWs2E5tO/ok9w17NdRR1ubEa+qPjy8D9LSHWkIqphW
AYXYiUMiWZUaC26pizUR8T+xgGEari8aeOq3ryDEHwkaT2+PiS7vqHVbB6Vrr6KX
4vbedeMgkhs+l2zjF9ubuDncRCYEA6puM3SryJ4CKK34q6vFES/X52MldzJ8VbzE
85o8jvHqOl8sZYxvoOJ13r64Q36FsUbYxGog127NONPj0F2aLb0FMefrJqLHfH1A
nloB1JlDhkr7a8yiTcpvMWwtoeB97z6KIKXKUtDV+u9y3MHkJoHBM6ghiDYXuSbv
+f5Zn1vF1CdCMYvYacuajYN6dT3gkuu5mw+QbbLCMsM/Uo3SExbEA130nwD8B/iD
ZD64VmfuCubM6c27oh8MUw29jE4U6/cxFNAB2wPUmfaigO0sKwbyOh215Wle7HGG
pMCqAqD1vR6v4kteiexwmovy5L4xa+ll3Wlru0XeQI390G96pzB221zMGWEqJHiq
KeHzyjRtywu4i7WBki5vTHvSW4pCv6pBNIF7TB6l/lxIjjoE8fT+9fcTT7AlfmjQ
acI3EZIZLSUdbct0IiKl13pVJwDGiafxV4daL+e7JZyqzBwU6lWkA2n3eD+M0zhD
ewKUAnEi3Y39Zul884lKXZqNsauTsCEHLIn92O55JQrTwD6VtkVyWG+yJGlHlnuq
6vUxswaYAIeGfUv9NAG4eHy883zsslfeqAURfUHnujgGqKoQQRawx65rGxiWxUAF
HUf68TgqgaAUH+4HgwxPnksqTe2tmhfhEVXYJzEIoZ7bfa/EqYIkLuhwEiwD2vEt
G+QMBEDhiOhXrHy7WSFM7LXWEN2hzzCM8fPbLfQ4IXepXjxgkr0wOj8XJw7CUrCR
RcAouucO0Cy4EYbubBeh+HNi7LNWp88czlLOPiapEyXvC4UUkj0x2dMHzmOAjtNf
HrZn2nc4mTJy0DBUL40otW/3496xYuKa/A8P83v5thtcTQj2E2VV0LETXoQyRkeJ
eMhhX8ip1lbw1+8cJmt1BLjyzPA25kbdNyEoca3resSZYJEuS/dFFBVSv/MktnQp
f3rd1KKIp1/tynKGk0MQaAZ+Q1KQGgW12T+lpk/k/6dMjxLVbD15rYDP/q9sagpq
3F/V7vakHUX3dE00hVQQaug0uMSB/WH4Bmqh20kfa4IQAVrBEavGgPh2AbH8Q64e
D8A7nffthDBt+T8xvxbjBP5BCdrG/rJjl6i/zeZCFK1Mm0txff6r3hriYKN2ASHu
rtdwYNKQd5EnXwhT8dU9+adAykFXMrKpis7+HcGrcxAOggxqEUMjZtocFKdwTp6p
wjNEzITwFffedt5wCagR2md1LsG9U31qhVgS062TYh/lqPaBMQeWQtjKk8/BxaYm
c90Q4Q2mPmvr+zBsOYIAYCwdHYCJoZZgFTJ5hQmrc43ygixQe7cb4n2gAKdINBfI
VJtBCPGdZrm5t1r9VXXPbIadHGeoagZXPDC7gDY3J4/7RyDPA7p8udazm8wPsMdX
dPYfol8se6+kkNK8tGrVhJRmkT7IEMyhTyB1HiH6CuvnJzmURFLKokoW0C87okzV
fjhAP8TCYUdmoi/Z3f2WBG+4PQAZkGNDfwYUXM3o9bh6hF7XgD/7hzH1Ntf8hMN1
1aFSPI1EEH1voSJcFBbMhLMgxPYkmFVvvLs1IJ8e0UTLN3V2QDTRyQcVuU1RlVri
Ndb3FvIWiEt248jLDk1edP3bymAtRTUsX5EpzbBWkADVf87h+9qxEBt+pLp6hBYe
CvjGkN1XsFxtqyOnwtFtZR1MEtlM56CCbY7eIIdtjWBmt2CmBB5YDnc1T0q9oSHS
8eK8sOgqdpzJAaTSz6her0ThBGehfo8knwjWiz0m2VuP25IP1lnJ1XbI6XE8OBnj
AnggKVCFT7k8KbA47ceWRVoIz7kxTv6zhgbrfjGLXZKE5eFEFpuG8Gh8oeN4Kkgw
tsloF8OKenT52ShHoI3EXjofvy80F8TQQoD1KPiQXQWSgAD4PuHjQkIHI3tXEddb
PNACZEwJI73qc9xRzW4+3HU+xXt11S4G+mAOzJjTtlwsWJ4wcqd7DpTgWwaEtWB5
bb/Fwig0/fwEhP/lBLFZfsz2Ts1bG5shmIYSWTPkfzDCltiQQvDn3LCyZrC4jlTz
bR8Xuhxa5CGp2fvBavO0Jr8luuHlkuCx5HCUbwQreYzBm5XUoJ4BQcxdlCgkDRPN
rZxUrtT1GKWSYvSEfzwoHa88u8ZxLr4YW8kc4VTAmFCCx84SC7Y0TEY3gjg6+hCI
ppMhptCCFW2R8sXzB+eDUUexa6mifAs/1WzpB0OFogpj4pYa9qqT8GC1lrkYq/AB
3um5ctjjaW2mpjEW5pqNZ8bAHYqAOHtqoopPhAeHVyuyOdEH1weN/I6NPfrmVQAc
q7RyIHK9lewntEcbzvNKyG/GXCsUFSP3KEoi67YLKKaqXUrDs5AaZp1W2ZN4MOcQ
7UbllmR8lI7Pennw2hG0RNn0bFGpSwgwb3IrKzK/cDzpoIKmdtqrS6fqqpCYt2Ah
9wOPcOYPhjn2dEN54TKxfCZm3N4KNEhsttFf7fzRbOZpswaV5VW3KQYq+kQ3m6LA
hStPCxSKH+WBLQKHY3wC5rETLkE4H093K8iBHpOJngwGPxEYNyOocicOZt1dfEDd
H5wBxNkMcP2X5KFBwZsVGb3USW1KWjhbgwP5wnFPa45/RjMiBjRNeOME2bAZlA9Y
x44p0nj+aGmXUcHVd0f43ugIeLRJeUSx3PXbBAJr5iJRqcxqC/QE2QMvOSXhwsa1
Dl9B+w8gGBhUaMduFJ424W5KAIwYQzA96pPvMS5SPLdaS5mJt0OYhUFGLjtVdbXP
i+wH8977AeTs1s8J3NXNq7EDOhX7G3bK1hbY4htmlqLss3KsQ6WYX4IlnDyhopEV
pvDIPCaZ2Q5zFYZvjgXjttURdXZicd/4CDuQzyEg/UGQZZ1SX0ws5qYJel7Vs2Bd
PbWXkFV5c2/q9p7qKzAF/6IawCzQrHMsqRIRdjPVJTNe/MYpkYPMzJuNfc1PPGvf
vy6dxSouQGJy2RVktrMQqJumvkJQ99XP6txxhDCoyse7A96Lkmfox9Nf2zcrFq9T
agoT3oPvdFDM++GtzsxIzKue6Z7Bo/h6fP0FXqhm+wBgz2xX/ZKMB2ntti6SgS0r
v3B9vVvRP9MmRUPMKa6T8o7nQtEUoa2BYhecm16vj5VAYdA3JKu5R+v0zpL08ReU
R/L2rJbaetccJwXLCeHaiJbjAi0l88SbmjP/6AbLHyhbfknDOjE6Oig0x83L9Eqr
s564826uy3BEstBYOOPQMJm0JF/YwBBot05gibTedgs3L88HpBqgxkI7A3NejB4h
61pWi7pPq4ViAEc2FEe8mQ/JR+lHjGzy8iTojlbJDGOO7LZnVa7oPnTIUfhWOAM7
O1groMKk7mtwVeLRjluIo0xlZn63PG3B/BmNkg3rOZSMSTgGkq7wOy6mwc8RaLRG
chuNhniQr/C4kB8mzQEjKvMjQMD8vd+9Glfv/iORgt9J4xy5idkHQAIlf9QlTlVb
aH2wzIPhSkiTnx6cguJgK3CvRBEDZ0w6HBwkQrw4pjOXkKRNMA6tAbT37XiP5O43
9D/CcU892QOy6n6BW+l+H+uloexSRx0iG21TgPEbrhMUzrJvf9MHa7e670cjJzGI
EJ1vrWMo4FufLzSeotL9lSqMnZ/92zyv4tTzgp1pcXAwu25mWcQHjm77wN6t0nI0
1ZN12u0YAZSA8+4In9Z/Baf7oewLAWW6RnfynmzAHC9avbAB/sKnDA6OGko0sDbi
AkhWTmY/i5R7D7pJAONX6dUH6C9M3tVeRQlUp7OZ4KRbfvNgVRlqaUV799eyG78L
y9C9jDy9FsQ5c9mWr20MthNe+sig/+ZutbYmTfQPONbh8iOa0y+P24qKMQCaeo77
7yjioaeYD2b0GI+sNzYXvZLz2QAu4JVnvazFBc9MKGx9W5hHV7GCR2O1NEW5dZzo
fkeOOXVDyHc9uFlhSF8PLD7dJxL4ck8eeJNQ7erNN/YA2VWX1RMBx2itNNkjYYTi
KfwJcZTpzCnHts1l2tZ97EFWZLRuq7ssZXn/2nBU6W4DqMW3d53kAz2zsZwbPjXs
5oaSBOt1JGU81vtBE4NFEhSjg/Ubc7So3EaRlOz4GR+Te4cj3mDFWzmuDJiitJ5U
vHovheUxmi/1KmOx/f9TtI0Km0z58cOepKeCVOGUAc5HtckK20suJwHj+L7Q5WNb
2rS7AeyuBh0K+BPyp1UvwcSaZ0qobhLeFPHUA+0gyDOwxCpLxV/Ib8ud68UZznkv
Ud8E/rninCdkbBEPr6e6MVfYWBMPWyOPjOpqll0IESsuf6lug2F0Qv3slSJrAwRw
0sjhaPJ7bFL+yTtoOxOIFzJEyoRrsz4UM3GW3yIPeeOr6hFe8aWYhVW3LFeoFDAt
rAP6Wj4jv2ff/XtgJuLPjt9S7YC6z5CUdJbD2ghyplyquYUS+b5zYnc2r//4p3WC
F72EnSu+Ec7lJsxs3TxR5wyM0qknVnrupngWbA6/8hvGnxgsq4NTqN53G2cS0CN+
DzyZnc3uZy47rS7iuNvk+yq+3EPkFRkTCg9YhwuVwT+MPGTVw0o0MRjX9Jk+22KP
TjAzkXUgqCUD7QJ4JzaI5W1Qiqonffz4fl0wk3Ycq+b5iudtaJmdxiEJUCTUOPBk
59aIBlVPvEdKQjin+me08l442OwT3+bUP+9metej04DulQmbOa7AKdUnX9ApvhoA
F+yoapH7KT8wX/v3vke2hlrU0PqxMSlSI/97BmIlLx5mHY4rOMQZls0dSlHkZSWB
+sC/lE+NIDRMjYQ4ikWxMCE/tMeqTUUX2A+X51nucABAD/Y8/iiov0oYorUYgkcm
Ko3FShySqNH0MvB3vt4SwIsivJy0nl8eGKd11lFRjbfc4U3PTPl4zFvHimN1ARhU
WbCch3sOC5UkfEfeGBogphxbCm69yFojD83ZYvzhcMzLOnSvf1wpb6/uOQ/puGgW
4cTsI2PS4fKbZvvtmZaq+bj47kld7qyJqhFL0PG6j+qkBjjCEtqd6sFr05k63yFe
BXi6CAZGY62eMdHKdyJFO9EZ2vz7V+9uQEKtF8qQYhKiOqRYXEAKjPNZ28bUfMMz
Slpqf6hYoiX993HcmEbWp/fs4LmTEEtWj9aXnCFGCe/gL8CGnd58Nui1oawUgQNy
x8xdTzHNoTSLuehRkHMt+8eaRWkhi0yrE1EgkNBJOQN4aPJ/8arA+AA8ukcRq/Jn
EJCrl2UKBJR0sTeECunqrl/DOdfo8q7oqxKWN3ZV7xoP5ASmrXeZAJrZHKhoQBEa
8vzU1VVqzbI/DnvX7DGXdXnmTz8MCvvdwe0jrqDJDxm/QcnwPo/fjVgGUC63w77y
xhEpjRLJQLdY7etqQ+XdXEGYWRZSNL3TRiuciGZ0phU/W1Q1iNRcjObvdSWnQQp0
3NK6u3Eh4a6n6e83yzunbzZH4jhK1kYni3DO6nT3CswJfToOIX0CAvfEMhc0XA10
FqvbI82lLZzWPCutuU5taVsrMFiYVD6Ym6mlp3/8EsaMEE9FfyU3yw4gtdBZh8SP
u4cBppWqEsAC0pVbRyYbEhpmlDQ9MqjhfnGoAgenZE4KHpCwJE06nP966TUvWeJK
uz+se2em0kB90KHERnWnboLZ4Ys0Mk+8u4KjaZVNoW0542NfDjLLxL21K5IlMGZW
3TOFHG1sdyacv6FVrSNuNST3tpEKZ8JZhUDqCyjupx0unAvCpJJe20Cm4aFhzHrn
ol/NXlEURea0ETDmlVMW86RVZoHEKPBNUsQxfIYI8BaPujxU6yDxF7GyhXAiB0H4
OXi7+1B7SZKp45Rh5X2wbYjvbxn/bjd/gM5qGaaJS3Zlf5toaMwZs1OtB3iqJP64
Uh1d1ZidO2wAQ61scNr07CK1mL+pgBe5Lav2iJ8r/mCuVcOXcidtYLo52AJhMdp4
xipvL016F/QB3MB4gWehr0po4IQBRGSPjIj6SyYbSMxRotpUhEOkHkpMrYaarTNo
VVSPbpE+dDSfssX+RR7ZzoLRKrNVtlbFxk8kCNaGxC6kvdIoNvJO296HeIKDYbKr
kkAVwCUg1waleF4bJfRdSrc8TDs5KxehikrsG1sW8s7KbKaxIBK2wk6qW2MQ2n58
imf8gXqk9AXKq2bqdJJbFsUnqfEqES5BT/35FPUm/gAQtotelnE8R33f/zAFDuVu
jxIPLg1wi0bz1Rh3ETPwRUolcql1Zzv28anTB8GpF37yTY8CxJWIeCWI4gXxEDDu
9MWGXlUqlyobRsnSdUiy8KjiJNqTY648DpLaBrKgIlOMANWCXnXmoyHfAYUF+yyW
1ow+sslnz4x9ynvnuoGBB5xT+LCxrL5t4ZD3TMC1Ua8q+3MPV93dWFMWK11TxcNt
WV7ErxLXlGPZ+SKHIooKYOJ6KyJewhf1D4W5YA7mdBWKbEFGEwwjGoEj9HQOxX8u
pFHj4+yIIJYwpeptrRKVdfOU+4uXV2W19tgsBiucfDnenbMGipBqBEz3ZGq+9Dgk
y7UcihaXsDyRgXjYz0FP7mOxZCuej4ywpM9c0n8wiTEVIXpOYC+HPP/+gZQKhj3F
p0BjHLOZCatEypNGYkgpRaLEIBm23wYRs/h+mMOJ9dklwYCMZJXLAVszn446DGGm
Mt7Cl9SGI2GS0EgEPv61MquGvCs3NYJoWzmQpp4VM1ypQk0EzUcXwCuEpDfl8/DV
jl+WC3WYgSRO6Pgv4VfSqIzTuAcpm4+h/ZLtJLsAwKvnz5HGaKk+0HFm7Y/zpAzr
Fw89J27QDyc2fOrm3QKemIdZkloP28tP8vzONV8TL/BgwvPP4pQ5OAIGnlXdNyid
Mh1yZk8fj4F2B5aJAbeDvX+Jget8dJtNnl1xrHK6zmCCDnts/BWoMKox2TphMiFG
Xf+MEHBTci+qv3iocTDhc2NJQrZ0cVvtkIE2PnFNMIYllkcEle9/hbwynDZIb/RW
vFoTosCv8IBJwLdo4Ava5vaWMIJnJLlcdnB/8iKdaRGNfBegix+ZM9i6rhrugzFR
YddAY7ujmCxXA5zA7gR0KZCLAkdDG0nxS4/EORSHXHocbeqWbIR7C7ly3osBsqQ2
+PerzsFmYHJggjiRCM4xSQyuo2EPcKiJ1gKwco9XETp1ufCJ6nFBulNAJkIjF7lr
abEQ8OB6DA9zz4nFGeII7JzUc3m2nOUYecKtvw3pTbJnmdTjxB29cGzLVITqUP8m
8Rn3UWl12pAR6SoYUbnBX3VbCT3ISvF64CNkSGvRt19atUBacH92owu+giETy3+H
1PGwGdDy4MjPZBxHPK9oCXcmaxn2N6ItfllRV+ohMCtsRwCpa0cO6lTJ0LAX4lT7
Y/LzHFK2TkA6YK8xmxLr3Rw98jmFaV/+cEopabESz/kifessvM0CDkBDirmEW6MY
XwWKCLXDGYB+wkna+ATmv79UgBraX3OPt9HlKTxDS0TC/ZMs4urk+K18Luemhagr
VcYZUPq4X6X5rARBIF8WX3FYn/YZJy+Ul1qDk2BLZoqU+ojagQFtPQ1lQsupi0XU
+jFXjh7brECkJdI4d7lg6s4FXAQr76XF6aiAlvNbtYSF7PrdlLE9hTq83L7IoGOR
jhZ8XP5dYkNM7AyNdJVrguOUVEgtvS1gbhUxhZzMYdGyT8CW/NpmCwVwCVpxV43D
zFFCeXxUylAjm7DLB9RDLkN8SyXbArFN3N6nqw83lNUYxK0U5EwjrmzO1tl9fZ5m
vrCwASbLWX6B9J+h0Ka7BJ0vVmza6+xTuaykSlwLRW3tJ1rq4Xp7XPhz2GzHNZSl
N0EHIGYTBxe/F4y26SSw+/iajVlVClH24YB6h5Pm7xJYvnlC2zfzXULd0mnhD4r8
iIraGgNeiZe0s8Z4iRB2/ONYhP6ZxiyPBc+lU54pwsM2vf9iVvwBl5j9jkEEnRzL
wrorHVqS4t2iHmh0B7C2MuSZRcUrY73zPgfea9J4QlpWB1e/Hm7XOJ5BjsbwoWpi
SznZavPT8nhIqpFhYvkcYdQ+XaahMTXHiwm3LCCr72jcvtsoUxFi6g2rZZJDZkcv
pknQbinlVwKWnDb22fUrxhtzSbhffpnAMV4B6j4dwXS6KlmW6u2IaPZ9BJMxjFVi
OWiPjRYsZc4rOBgIIIJn/HLoMT7fDKAKZBXzjz5Pyjzz5f0AjBa8c+iqQ+hUYVu9
Y1E39Xi1MFjeT9/7+pHxBAlscDtPEXTGLE92qViSIkBvPt53KwzpLX4coZ5IN34Q
aUjpVvK76M2rfJh+U7cPXOo4f4Z+662yTrBMsVrn0UDZcwEoOEomzGYETXCxAheD
QG2q6R7PJoHh4d8xzd6CWpNiJ5fp115FwVD48MXuPgF1CI1x0/3fy//werIN1Szd
wa6QJblT7NwWFxzTOSwBOzoFiV0ScYyrA/vLkm6Lm15UxX1zn+YqWyUA5wk7Wg1I
MB+3zsvxwzzK+phtjj1KUFOH4SzZmBN/QkKqw5Qy6/F/3VPPO1jrcH3Nne27gNNb
7L78QTlHrtNMWkAWwbGG2LwCHTahhgnS0cDkmrjSVQ4uOAPJBCFGO+aQ/dx6oNZM
wAXaQBn0QXTVOuAiT/deftWxfh+qiVbklovFoKWVEI1Zursr6gNHJp7Ms5mWYpL6
1WpsBbbsjLJBWyVLLlyAxn7lUjqQOnckwwxfwC5ZFYdF33NsdbZVQ3+rYrYm9ahz
yyUe8lWHUt+nUQpxBpFrBPEXvVhOlmqP4ROgfuQZK1uzLFy7xExQBFwU7KgccxKt
II+fUnoArU8IVP3H/ABjTq7GxLo2o32w9jCb850+xYM3OGVWiL4sBqpmwURLNEaB
pip6ZobzQEs3NCmJnQlkeBa8nEcQpR4RgYysbBfFQ1SEGAU+sqq9PBBbxeDLYkZg
HVaojCwwaiYWUNwlwXe6eNSkZDT1Uh+cTyodhMx2pTR3eVOu5B7F08ioltjlHozX
4Tlgg4T8mOeVKTmf1v6tw7eFwaJfBdWSXTU47GxkBImkF0IDYqiWGZECoD+pv3hE
00/AV1p/R7Y00pYefAUIeDSb/Lu/xnKCuiLqhhmhrumwfHuyRnC4x4prfrYuU9i4
Wt2jj+F+dv1VDAYzaVuHEkDJ+C/hlxhiDaMZK5dnfZRzyNClWH2jbziQE2Z/ZIrH
kHb6sU6ac3wuiveotVc3X2UYJv/sd9d8Ub7TCV5nTP9CC1aEVveyitjMOf2UjG+0
YOT+lrMLQ1gZCO5jdpNoaCmxXCJlbqfdMUi7rnxxU9c3dIFG1C1tjmRPqwAOVKTB
yRyuUzrSLRx7S+z94i4fPDbZsKFO2xECd6Joln23unoPrRSer2mcJgHyjTftgQi4
u9kHqlqT51/IJn7ltfvD4npO+c+6KVjW3tTUnMAcifEhKkHjd0emQyvhSoXDlJ0e
TuKCHis/M88gAvm2+0x3nJPpZ6q8IrmPwowBxJRdYZsGEZ5qR4PBcQtpeo0hfQz8
l4IL7bIze2G+lnoe6q8s/D2RXkZyx1j+KGa/FT/GAcHBE4omh8GHiDMhNyWHh6FC
aryLEEG/6+yaWlN0g+Hm36KOjWo7Zq30cyWiaerooEinZ+fHxa9xAkCSxjQQpFkE
uk4O6AEzuIJ1l4Y6UzZ+ro/nSwgglB7dNjm9HmWljkulycOSHOZbcGATTTpU4nCC
0vH3oIFwwwxVOgb+NiCDiv7lmLTprIJ35wAFACfgyudvPYvTfsQuo2cfUKQFaFKL
BNbDObLZmDHhP6neLYmBVLEuFmrsG2wyttP0cBUiJspbRUOMHfCpXLXlchFB2GdL
RhykYzulhPxklkd+tmpQ2k73qjLOSokxI7hkCJ64XZGsUGZROrGc3a3ZaIo0l5q6
ov6v1uem2y70tpolpavZIlOR7csBhosjplRDmivEIKRFAdl/miS4zcH91UbF/iEv
DfTSx3enbT2pgA8JUaOcZlzfAwp1ktWfUsI12FOs2xisUJ2XCd/UUO9RQ+WqL0/A
AMYzWTqWn24n+IkpZ9uTtG4FsZ7c8olxIhzgGeyyHYdoxUS/Emnwzn9lqnM6FgVs
NzRk5xgRjYI2MdHbNPeDn4U+4lK4RJiEPZMJFUscT/58BJbL3okYayjymHxjm1qd
BhBpl9te42Q+RY032iPitIwv7aZN5tJJ0i6SOpzV2/Km30znbM8Ekx9iCAi6bg+K
p+HgmqvfaHTOJWwoo/JCxBS3hMZOCOZLCF765e6FTCZV2uRDRa2Q3VMqbTYe8cVT
it/9oDVJ/tly5UydKmOF7NI7+CdHJtcvQlH8B9apKWlvY6B7EdUX3YYFHoz0W72G
Oj8vSsqTimt06LHXONXIOa6Jk/1hkQ5DFnqHvwGFdqL4gTWiOFXgqF0IhGMyJtoa
U3Jxb3zywrCVeFfTAx53ZX7t/xsshQbLWPuOAZm345GuMjIciLE9jTEHl+98pAuY
wkE2DGxEQKdSIzx0rl6eo8+OLhE1bZP7prbdmtRVdSbnIt/pXv6oP+HcuCREQihh
XPydNXV9d+moNqpb5h/MbL7rAZw9AP9ruYtmAG4S5aRZGKIsHJIFeq7ueNjczXxl
r5rZzMCNg19GfZQq6VPBVthU9uiTSr01ZxRQW4nu/P9uVTRDcvn3MIPbFx70GcuD
DlwvOtl1DrXbTDMT1ZOHPZMZwtffUz0bvuMkdEyHm712t2PITdgsDS4pOLzMVAMK
V8YOP9k3LTPftojjMTU7+64p9p3btxbQ8FuVUTJO/DMbnnux9dJEb2uPfUoxaUa/
G/9ScQdKFMMfHkA4jKJ02JgzZ4lCoLQQR+dbTqQC7aZklQQSTTDN/CtYVRyPq8Y6
K63wfci64WIfdMUerwn1/Krf0REPguld3w+fHHXYgdlCRVeG3v8Cyi1OSdmp/k5L
QTdxZTgP6YYAnb4Cwp/pikNYPZ2raHcJRi740DdmZ9F6mlSGcupHEceF2fKLGY9p
xfRpxrg7Y8+cO9tuEbvMAeClc3m2uPLlNb/7RjAaD/s4k7Ch3AT/rgx8i4MCPfHI
Ebtua5Ie+D3AqzfO4PavIlUkJv1PF21rqUho+z6/De7hifhwB+jV65rkjtT7hpK3
EdsgyFcno4SupwUt95mJHNyyX55kPek8T6TW8/g/WcedQls1MENWUYRUdvxNwNwU
7pzlkHeDAA9mCDMSqEUCQo+2SAWFF5W32Qs1WFQ4U7OoDZgsZtljLNzfGOBZI4HM
9KbBhvUhqc2b2TeAvAz1JULW7lyGWib4GdiiQwYEgv3q6kL/FEBOwUXX1LdbuiHl
Vpj73NczkIk+pXuoQZdkLAGkfuZhWs3mv3cKOS9Vv8KdvRrV9NJjqZMV4xRaSZA0
gDLpelQkexWOv1MYFiGPge6wKzbIDgaD9YTS/fcrM31N2Kl0KzMEkRtBR4KLhqdc
mF9Etz8J75e+0LU+KM4tvnqNLme6txv5LUPK5MOYRpL7/owmG2dy27vTOCYQ33hQ
5c2bL/rTrSLW7zHsparPMY6F2DVJ88jzugN8q97J/v1xXgeMzbw3bHCdK0tADI3a
/o/KgqI4Z80cTr4cmr79t8Omz0wQJsRcuvlqI83afPaQ0G8VKIcajNreWhDRmRHd
AK3b1unn/JbKxMU8s3RI7yUJdavs03XpbjSYIzumqv3Ncmn8yw/mSOGU7J8ia+bI
PxuPuKaDrXSUETs6xmCDaos2egX52o9Ocu4oOymIzzzPGfHazJJFw9RgvDrYuecD
XFZIGTpDVUc9xDr1PUA7zMR4JuvMzFXCHDQsh2Bw0ZdWruMoNTe7kOFFefL9EOal
IJMAGk4PezUT5vj2Y9qmdrf2LDiJ5tVZvoUipi9QdpcbF3aXZazSV0hsH4z4SoO6
RBjCfdhaKKGXIOs1gh78yW3ydPB/6ReudafvO/1kz5OVaqtJ6q4xtrxRW/7yrJXQ
M8MmDwSM4g5VfHUgApQ+ZCiKazQgLIjP7xg50GORedoTCIDsIQcxLW4mQXC+pQtU
uv6YB1TgIMY+V4srGxizaK4bP+X81X7j29qQlcVerdbfhrmHt7OrA2mL7ynnLEE3
MdAXFd31Z7Pcp28MmcYrANQTrRbYOxtniV8DT4R1YkPHK4KlaDPf8cRiqbUDOkB0
KVSprs+2Pwy6/lISNdlu83kbuA8doPJJKELqTsCoJnzixIPyrPWA4Oy5fIf7seOw
MFpokY+AJPezaUCjcbPR9YH3ffplxvgpDYbpV7OuDjq5kUiGrt3VHn1wWSGqvMUe
RSUJ3NIZuFqoVATsMAIo/MZZi3blvSXvY1GnidWrYL/pYHZ7N5Q9CfuDfF7zb5oS
0S8lJwDl3JOsxtUoLZ+tAnhqbYJ5CLYGM+yvaCkQLHfzTvLu9wsRVFttmixPa1nq
dNQkx1hXukywxmUMHSh4CgkMg4d2Ppec/5ZDRTNwNG+Z/Wy5IobbFbaZMc/PXc9l
go8uFmUHgb6MK0Of+dkcb86AIlWu+SQZbZIGT6Kos6u75NLujTtTWRQYuBYTOG6X
hZ9Nvan0ccQlleOadfmZXAzV5ijRL/6FrTmXRUxxYCRmTQfkPH9uN473N4x2bkgP
u8cJlnqQbgoIRBNCdnv/KbT/vCSAhFmZorZwyEOUI4EcMyWdOBwFQscA/PULJQeX
fgJTFyQe9d/dleFULeNoFHfjtQas11d7CC70rg/be1prpujc5W4niixHsJNYSN+l
1f5YZplU0+PIzxO4sQzZMzxGcBQt428I6pZch9sohuGNoz25yCAEUSWqdVT6VnTt
sf/o1FsTTBdhtI95UU0Vs/RBAMinmGx09gWwiQr11AVs8AwhB7fpWIncU4cKLAkQ
Plc0jt1OGZN3jVdkXsNOgPD/z/cmkfUVZDtLe2kD316VEDbOGeitc+25tzgAaoHz
W2AbuGizfkEa++gpF4cuCRvXgHm2N+0frPWT0/0U+qZwcK590GNCFkkHnXrHyJ6B
Fxon4/BikzyoOCtBpnIVSDzLZ+rNMaILECweLKAcew0uBvHLEdvQM8ztItvshlF7
+7PSUyvpRsptoNVqPGu8qY0xDqLQmadK9VqxYCqVAHYRIMAbdk4jtQUZLaxbcZNx
RrRHh+JDY7HHSyc6EOeNTD+P8IxA/EPGW58SpLvMA2mK7C3/LtHebiPVKDFkt8sJ
ayWWGm/XvFL9Oc72i4vI2Za43HNslKe8QjrbVqkoJHZRMiO3aQNeN9UiImWvgIkA
YvClro64jfbG1Cdy/8GfociALsK5jJeatnZOwdK1ohtksZTvjnDAxGjXcya798St
1DsOYKsVxSMxYxjm42qiybTV1YfDqtApJdTwrQeyyCnAREfbNCqNVtShiTegdqD3
X+zuvODWzvSXevNz/MrGc6W5yc3MJR6ppnZ4MH52ZbbXQEl7Cwzmq+PL0u/R3fzn
90RqmWAKDriQw4NRBp8Ncjh42F51BcpAxPDvXuNPAwMVDtgaZ9zM0BHrpzpBmTHG
2ZF32BIFEndnYUK/rbbeR4zg0XTL+qwu++S10o1s0EqArvkULajSspBdtrVEOcqj
0Hu05ygKgNUnmbZIbBpu8XwUUrw1t5ypGFBWNB6DrLY3Z9hDylfvc4+Sy9eZFNUN
lTcvnReTLz1p9VmOu/7pbc6x9IWRCA0sqhgSqObE1EeypQ0gzJaH0eN7WkQ5S85A
0HBWVMoOcZ5wFYTC1HjbMUwRmPVk0kBdOUPY0yJDAcpK+0W3MbK4sIEwRLUtZ6Lu
9z0zJKZdqHkTx6461uIEqfTZs/+UQyp9q16C4ejNIpyZi3/lxlKcHNzD5nec0Z1v
Bwk92WTuDl/GNYuxTGPuuy1bjwqmKPkwYqSJbers1aQnt72IRV70hXWHwSpVxOnS
H6UjhJE7EyqHXgOd1lk949rTpODvEhtC3bYCoVuQqVuNcbBFd7mlAsFKr82Q4UwL
qnizUxYAdhEfZezCAv/fmM+W/J93jnflnm4Ct/lFhGLPy/7YYEIfhZ25om4Z0cWQ
pkJdKR6XAhBfpEB9jHHjPom7h9vNNpNdXybvvGYXXn4FuYHdZTjp+EUSDCDbF5v6
sI8iB5mc7ri0ZL8FIWZHHisOPyTwWSKk8jRKSbMT0h07Wd0DmoR9exAL3YQHMwiB
5Fx3UypO0RW98rlwyIUCYmPLStcM3caNBkWLLF9c7xkpcD6421cJa2cRennYfqou
4VQ7OeYbFuoCGnRTxJcmP5zJUvoJivmLE/mRzF1IZ13GgAdkFr4ivWwLaPZyjFPB
ywYQ0+bIOb1asRugHPoF0fAqaL4v8fS/zYU3BlswnlNjCUbxrcMzVTqFN1abr7Wz
1Lp9cCbGTZV9MryAGmU/6EQu+FGNQe4VsDuQq2uv+DGydeK9yfltCztgK6Dja79m
DOWvqkoW+u4TK1fQJUe8hwrt/G2B7PQO6eKzLmatuCTAZVxMO1KwJPLsFwKg9ezo
VDXiiXvs/sL/ieeJJAmub3p4N+3mU2lXmYqoCwMsYDHE1KNiPvjReIGJigMLv6eO
unCxREhsqGOh5HTE1z8BxA==
`pragma protect end_protected
