// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W4kt3UTycSy97jBNZLBXx1Cf4HtjN0lPh8zVhfPpPch4e8JTBQ5nhZXCNx7F+sf7
Pf43wElzEydocSaPvrj/0Scm8/1QMTQQO4Oe/S5KIT2yU6orXL3LvLTWc5r0bQwW
ArI0UX3Q0LIaixGxE2WIXKXA/WOjI0vZZ6sIObMYRTs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15872)
j+9/qLFORT5WZwx/GDFT8duw80djfxOjK+kYxDM94x/4MiuEK9LKdXvHxRKtYfHX
PArbbNnFk3pbIBPvib3HDSTCnY68jPcFShxx0qAO9xFVPdPOVObSBPRm3qebFtfx
wzHYl+INgXUjXc6HBTeo+oqga74oPQO8WLazxgT+9We5sqyR32Z2az4pPmx2nbmT
BrJ9/XTVmBauoJWR0Q2OCOW8/1HOqv+OBdzw+Zs3jszoqu3ZamzQwHZEOldDBw5r
J/gmXOsT1HWbXDLv7Qr8wRKirmiYn4BbCQLA21PzHfNWk/FONJPyaidUEY6U/I8j
BX1iq1+4lVjwQewwX8AVqGK1SkJrMw849Mf9HtqOsr0N6TI6qRHVY8eWzyzwIdbh
OWCNn3d97aS0MAX1D66ZiDr1X737oOLeeK/VfCm6XurqkJyethL0vUo65tIMsNFc
NybEKa50emr+0F+87KYUByYAKCxAAccWjkT1qssTsPBD2q0H6HGhH81Kh5GKPGh2
Ze/heyI0j0hDcpe8mksT7jn2TtGF5QQnJcsZ8SRogpI6Nz86y5jFem/hl6K+qYfx
4FAttKqcwgKt6aP4xbeifQzS99A7PJvlEJYZlnFmOZlA0BaITHkbM6+pG+fTU+CJ
ksA6d8Pd7KCOoEzhoxg3P/4vai1A+Njy0AbCXqI9Nu1Cg74j53aeahS7SyBJTI+g
tYcfkStS7EYdFrP2qTYeU5w2E6wy8vRM92A4EFRAh3phhnqU6ioa/kbbPBA4gAT0
YjxdIgmoaj0P3BuFkJnNvGEByuIAp4PHyxclfUnMInrFht/8zxWx4UATItkTlZ5M
X3WBPqhgYz9Omp5k4o2qSSNErqjJc1jRNs3k3YkO3Zq/qA9zrQVluJ71Fwnnw2gP
8EgrHWccs9CC6fX7D0Auh11PzMxoHkVqi35P0Gc6/I9MAojFhAvViwWjNOz2vyP5
3QcwL+MNaPBDGBuB/vftfrIvLE8AHrR1UJ1FknjHFdfJ9OlXuxuREdQ4XlGMrZMG
8fgK31jXmyzGZdxB3Xrr6K6R1Gd8JOAEWrRYcqfzmIrUQxX2qNx6baPjWUrXyNlO
W87gMR/cqUIJ9w7Ep6p0vNHdHpFacosQcf1ycnatULIm3rFHSUZlRD7IeJdtsFd5
mVF7MokIXxEvgSnxkciWZhjAaDL87E/wg1hach9bNfKdS5KkVetprhTLfqPxlvQy
Tkjej+NIuiosS58d4HpSBfz6Gd3rUaoIPAcnOgZCKI8reC+9n8CSRjamdR4qTo0y
vcxIRUQLutrJV9abpqyHgM18QEtU0h2RgqmQjlDRGj21OzYcanhhpzjqoCBSceQ9
QEu63GGnp8hE+fh4tMuWCAY+tOrRw8tPrhs1R00wLcCYhAh+mvBmPMh0J9ppUOtC
xH6xHFfslQ9XDpAc9b3bCA1mcEYZ/BwdL8oLwWwuUrjuXWGFbz2v3y88ZYEDYtfy
penkXkdWUDZd1F7I7tlI+dxmP9S+jqOWxaFWEA1RLWtOLRAOXRSlVig3tuGIOB6h
1ljCQkI862TQDNvEpO1wXzLTAq9EVIEyHINY8e6ny1T4hruSfaSWXx3Zr8+Us5TU
pl3jlN/1HsUZMyEZNA6t907Na68XkbnwH2gyiaIxD+eT9+GMb1a+x6XKgoLZm3H6
piWYVUCeClXBjc0iLuHlqFWn9B3zk1AhirC9p5lCOli9oqC3oDZDjuCxupZQ2+gt
Zxfc2xRnOZ/g3awcL7CIoAmxOILlgfv7s8OYgC4cUrW60MPD8uG+44JVzgRYveJo
pq244O7Wrm39ijmXZCoaUSQ1CBK+2qgNCB3BvmKLTxFrIutHYg/wxElLHXDMFf/P
zp+J3jMCvk6q/Tle79NgEkoz9Q2Av/yEhRfPfNpPDRImTkF06NJtmqE2D0/OXK8k
pLRSCywKVO4mUjz8owsKC+zrzMGJ0c4EDJ58oxMObm8jCWq4yLxKZ711M/GOuQKT
BTSf2d24UjRJu7OlMxTjrRZhem3mBC+o2ntHaDDBqqNCQiA0MBSzqP9ACex1Ksfk
UVrkY1SWcjWR5CoXk3YJfxp1+6MVRItESKnvGw77aIuaLM3WsDKzypmsikSjsjI+
DfzWRX3fXuJsbKQq7FHImieTso7Zg2DB+ZCbYT195SXXVnmd+TJXBpkdbBmfz2BF
xZ9Apim8SN/fkENNxIxfkVqN10G1HDVQcPHu2P+OvkyvieN3L+He4jPKpNACOfIj
A+h24/NLnIXcVhrzc9YYRDX0PxCBtife/cnQR1487PJSQR7C/9RDYifI9n4Weyxl
4hNuI9FOBGbZsGvHOkj05Nz2hQIILkpwcMeWgEJCLBws1w8EuKuKjmaP/H6z6q9d
HzlV/1c2oUA9HsIsrr/3vV23DEZAT6r5A+UHiPCTuGU8mQ/Jf+A+m500ib8iSga7
PjqTHV78YFAalxZq4cQdUKqQrOlXKafzakDy1jyKe0FbCM4E/gtkB/mcm6E9srko
Mr3X1mviN8Ius+iVM9uEQwLMsvStyi8EhryuJN1097i/vwfbu1vcQ91F/iQz7Crj
vzDa2nTOc6GXBPTFKc9UOydHog/+8j0ZlnfkiIa92cWJlXfH6pURF1RCtsDTDdk7
0uqcpV44i3xW/ihPkw7umVhzq5p+krr9MFl477nm9AjrE3y9y5uuWsvx2+XGFHZl
tZNLMK15BPHnIkHNjYwExz5YSnlG+SK2T/b02JnJHPQ3Cz4TuVgsv52upVqJIIdk
mcZeN6TU1iMguj4Ey+WXId5NYTK92U4AIvhsKzR5MT0gZOSBsbaWbPtG8sDUGyZ7
L5hMB8rh/s0bcQpPLohCTmnUgERd++rDZrAVL2jnQehxzpgVzYeNDYwoWpVOtluT
P4RvhkHLVUev/pm1zR0p+ovf0jgoYBGdceQEyNXCGD2OvCELp+ddHmdPiW1luT8A
lx/MIA9BG0wSKIw7iZH1wNT8Xmu5n3+lUfQYwWCmTS2yrQH/HtFzSu58mlevRFfv
++3YIIH0Bfq0XFC4JiYAPw3ai6IXA3PxqISwn3w0aLom89hOVxBbSyJ8qstsUscW
t4ZPlhwIkSiNB8FdkKq7CYsWWeQgK691izh6xXbCZgn2qbyeNo5X8fiIQOHfeo3k
PV5aZUhxiP5J60hbSgAA1oMlEt7fpveptwj/4mqLJi98TnD6j8eAAed1HnZElx2N
TarVzCvVmlwBk/bC7ZNXLnxgeU3qFe5sSL9mIjwO9Bi4fHli69cWklgB0cYRZXfz
ZaUTC9pAjlgRlVE0FgoISnFU73sWyfQZJ8GhBnYlQZkeTLKzfxnCxBuPiMxKoXet
/PlvPNN+Dca+1Q1Ldh1Pq31DKu5y8gBw4VhPp3SIAgF2rmVG2vOidRVizkVMstdt
j6pyCvmCVMZhCel9qvNXh2ZIuCkc2kZ/3x98nZw9S6S9uG2vNee6JS8YF+Ypv7Z0
nfbzE7NJOxWbI24BtXv380pqMsgmYYdo8dA5tBLkghOG/wgvfSOavhdnUMoJWUOh
1NmQ28yZnhpcfwK5nOEoJ8oFUVyB44aT/OczqQGIGyrxKiY51fi/CuCOshqPubJj
4L7gjP+fsWIoxEHb3Lmp4kE82M7ZmSNR4QjCGNM+kx2n8FBh8j7uPbhKmy6peEMJ
6wryq2WBSJY1FYBgFEsoJ323lU+L3Pe6JBAQzD3YCxALxxfA3neeHkRixJBOxIOK
Cto95GO0HwpKSLmNH8FyNM/jIgnwmyD/wM4hvlyt+pkK69qexqkTIe5fn6Ks3VG0
UP4lNaUI3bprG/q9tY29jZB/yTjU+bv8La8j7EmU5LDrpAppLN8s19NKU1n+kPCX
85cBQAD8GPbMkbRWvDSqi+OotOxkQ8M/xuD9VquXmzx0FOLeI4e/VaSYQXzUIlJY
W33x4FSvadSAuTL3x1egLXWTNWm3/q04BQuCkPDQphBcxyOMScUG9A2V7j3GoTxq
iTHi7ZCD0blc7Y7wVS9CshakC9M3yrChrpNCbsPJ+353MMAAjxXPLJ9n6WmlTpEB
GdvoxNMU06YqDGPCcQs3pBO7OTl36/ZxMEMmOeNk/Z6iF25yH21t61AHD5pL0O50
bPHZnJr0NKKyedVkyaJ/g19G2iYAe/++jM2U8ibCZ9ry+ZXfoOlWsLAw5SebxXiy
wQkNyb6+JFSvDhuorVT6YohZOcym18lBNZDQo+jIaD4rKy+QbiBsD+Ks82b9/YTH
GiovBvgKlkMMBrfVqEMaaxti1vrrvDPWa0QrsY7LCUv04mwUi5CsR5A/7CYnfVjo
b2gZosFn7xBRR2VQavyiXSjnnktcTaap+7DujTdDJPP5zJtTmWm0HzVu/9giUPqM
tZHkpc1wTWv1TqVQ7B86B0XlKunqZUxyy1r3A8rxqRrxB1b6qvmYLGWEo8rS0dr/
UUxYNl7f4r5wtBSjCraXObHk+lOChMWoWjqNIARxVVwZvfA2xcmxbk3o3EfX0tap
HChW2DlxOZDkSchmfOJjUhrvTYB5m3M/tFce21Bt8GEvZvvPZ4ZjFgdze8E8+W1F
2OFNE/YpmIpAsUvaso2diW2YsPlwkJorltDpfc4wmWHYVOVi4rVl0w2mJzfh+t8b
LQK0+0pJ+mCoxEHlgzEdoW51TWyrhpBag/FabkV75kvvpVbTPh+rU+fC0iSI1ydI
P9sN4dykMuFUIPrZMpUY3aYwjByQ71+HNjMbSiN4c1EXIEfjAlklR+sqhBd6NAO5
ptafyBq6X0Wheg9bL024W2EV8VQvJHB/9l1e9J5tErUcswJVVvusJbs5RkJana9Y
Gd/EUeFDODOKsZP5iIt+nJV6skEtb3k7yAE6bu9yUonWPlnkVZ27Zy5+g7zuCrCD
ZasM7gk7z8uc6EkHc159tT2KnRec/PMWWvrKGO08qszU0FaiUjOH7sOO64byFMWl
/KF7WklyP4oDmoE1xqLH2lokteZFsT8amtMCPELoeTrCnchVj0gJe0WeWM4cZpCS
VIBgW28H4Q5hSqAyVzLucZHHXS5HSrc9LkoZamXgBt5gmFz7C3QaghlZRU7+5evk
vRpDIBal73BeSuC31yYEacAdAjzCXF4s2Wcc1i9Nsxn5V0S7gq4+qUT0aTlbJac8
uuIvYfd5nEvaJ52uey6yzQgyWeH9NG2gtbsPN80MM5grk9NjJEZBYLN9c15zBMvG
yqhtQFK6pPi8376Y/UyZZO3izGjvykjJceujxZ48ozC76SLfbBjv2+DTB7H4l551
8FtsMXnsw2Eh50U4fl5wqyDAEG94qiAryTnLi3EZcRj9pUP98LDbI2+FUj69lIvx
tA4mAHwpEmkVDGTn+8oRN/7QgAaBWgU1+CMm005ZlCOJQNsR0Pr1v2NC830d00Gp
8aDYZkSkKpUU7lETK7BEgKMAI0aui4y2x/+dmlP5fUrToD6wjgJICGUiKxgMXtWd
hF+UfZWcHw0mU3JWkpq93rDcQ5uKQ9FIaY+LcRvpkk+id2GnpigcAMmBTGvS4YOS
/3YpOmXvadoBr3ILqJ6FxNnlKTBxAHoxBGrBck01tvytEyvMHyHBJwdKydrZvV71
Duuawm74ZwlxDH2JRGEXFVOaUxouRPxVqLSe7hC9MYACqfLd/hynJwZYGmUL4Zja
+hB4xOWWZiA2JciPLs9d9X6RgTwcPmfZT9Ihm0rbZ2OmlBhPC4Z4M4mqG8BWABpa
eYeS9zq9oJMaijyML77BmVI8BoF09ulGeQ0SwPFxIf1sqZ0JjA445pKslshus62P
pKO2rnd7cz/cGkAF+N2mTC4Ot1EhWSdfN66fIfv27CZxDgxT8WnWwRMTMBXuJvEL
YJQcjEd8G4npaPilZB1PN/7EqnzC0//4pCGAqLlKJUBRYWsug4P2t8tcBW9JxhnN
/kbnKTyRUsy93TijvDHmbTUEd/+7XJwChrQ2k12NjAeMj1v3St2bdInGejWPssDg
GlrS9wa+Lop+ch0WJM3fzhTZw2o7UVxmfXdKLLXboaUwDTMUPCdWwYl7mEJHUMck
0mUM8sETL3Tbwt+pq1qAbtPW5ZmWw4tL+jpr51pslqSWeG9xthDzEgaUDqbeB2Sr
hbcZvqn+iOYKzZdfxfJ3tiIrLlMVZqpVgWUvpwuHA6DL7vHU/FgqJ1svSxuOBii6
sMD2LzBIcBL+htdVI6eApO79wvGT43SaYZ5E90j2OHYRoTI4SA/olLqUsDmruEnC
mrTDuyE/GPdcaiNPzrB96YGMIZtT7kezzw3gQdvLRwN4w4Y6nAmbN1ecTVCB+/VQ
hwBt0xPoe5AGXMhWUfTgyJdiKYQfdxOSFr3B8o/54rAYvUmu8GQ9tM+J5iIdCgya
6HUUulj6eWVOOrgXzvDnDKpdGBEVPfzLhWqh0slWCxDBzyw7RdUfaAXSkuhYzp/N
mqaY7GxMtI4e7mN8nS41NwKdFFqDeRaN8+m8PBimXE0bkxyCTll/+9SHF8s4a7sD
YxG98n/9Ht4H5S05r7L+tCrDCXKCl6ujqMtvp4eg+2zyYpJTddJGTdq6CtPVgK0E
SzG6nOVU7iBDle5FW9k3LGe292LDzEXETSgRArfv5PohBSUYpeGpooJUBhzyMR1p
FR7MWZ0SknSbhuFFSsvDwaQgfs63g2FdSWNoegHYmfkY01SMFPtMukXTjKny0c4K
lA6grzdJprLsXHXyZ/FkxBy5L0LyVNYae5yq6az6l3GobNDvV3SkPw4uxWzzkL/g
u3vox69xfSaaJSFtA3hK7KboZsgTnDm0AaIBj1vV48U8mS3GI0/9KfNLRX+k0flo
1ZzImKaAThTALEF4wf1Vxw6xIdCUlvlJQRh33xRRms7Wa+kQo6bgVU2Pc8RdojKY
X2hk2mYtaKTUdAOG/d+x5OdWL0bE7aeVpuYbbsFCfZxNuP3mrQ0cgrfuBpm20uAj
UIhsdteABCm3GdqTTvawNGUpMahrmEYMVYHzkwJgaybOOCqmSa+Bhq8MwSPNTts1
Y4fHwh7T8lS1hcGGJzDrP6V3zNn1L412wJg9MjHbGSV2SeAGbF6xy5wz6iX7c4Zi
rsjCrBXn4N5yOwpyJ/G9zspO5PF3QUHmPJ2y8VGIJshOXol9BBepZZvrkm4FpMRo
uJswSYDEss5O7BQqYi3pkNLIyqoFcqPv3Tn0hJ4/V3a3MDAwWjQQS180QZfvVBsR
zFE4gzo/3C57bC+/ckQPGFixo+Of+fDKZdsh242y6K3FYBS+WWAw3+Bxu7c27JFN
kAnAzkol0jwvcyIrPThLTH2fwsslC3t6C6A0OXXlhs+W/Q1qOPwfy8X5lXeUIRZL
QFQPhvyzV6h5+N3a8upnzsCmRXdzqwbILF2a0JcuBIhtQ90XrWAx5hRSqhM9D0Q1
YRVMxN1Ptw30HtNjnFUcF7BnV2li0JRhmmiTZYxTYrTUO83yf16P/H9nmPlvTlMb
s5EWy9VPgrivZ3z3qb/P2WCvoB2doZDMS+YRPVQKBpH5e5en99OJhOfaIR6agVcg
5RlMn6TV8JpeVu8/SzrEy4OfNRVVpjsPrGjVsT6TXqHEWQMxXPoJ5CNlwYfZJZ6k
l8chtqgunaBOMuQzp93B5oWerVA2b3GWLpCqxybY2ipoxwAaftUOToVoCp7ZTC6P
JJgIfhsEt5JeKK1fPJRbA/O9dyRJglA29zc8gSgB3MLzJzkY7IyDNxB85rr4aFRQ
/C0/qW4Ihvbm1sGNFeF4yWiMIWVEWmr+H/aTI7k3jJDb0L5YvND/T5Y3Al666z9I
8XX3QNBidhzVWLspesDy1fz9T/d8HFk1GEPSRd9x9HGDorhDyB7s9xwDiSmkZ05D
Owzagoq2PMAgQs7kFCbNwQ09BNtpKqj/JatsD7u1d7r2VFzDDi8KTJByir/jZa6o
M4frujn/ahCDpPoubYaR6qcCFUk/x0EowamM00/NTbFF+r4kOmFrK5qd5i3W3zyx
Zka1A0u8BvMgQI7EYYZ+wz4t5Rx9A2AkWrovHeeouQ41WFYu9OIdilPmynX/JUz0
Ji02ocSYIcB6NiYRrDWiHvXI7v43SXEuOFdtfFNuMYTRmZzyXvJn7VtM3vXBpwKZ
xaz80FLqqdYc+s4ywaWqgZOaYrnp1DUWB37YrKoH3gwNBh8yktgOBkKHQtg54Lje
Ocrjurj5vl/DmIX3tQd7o/m9lx7w11wCbcw2TQmHDunqOPmM0FjXTprQg61PIL1A
TUpWOKGKuAPpK9EulrKAP7eTzA2TXmnNqokk42f/Eyi5qkj9DLoXbBl8zUlm5Pil
X6hFfJDKS3UNPFx8YFH2Oj97GDrpE1r0KJVGfVpZQxWMObKJurMZpCGpWXWi8FKA
2/Jo/rDirh3q9mRADlSxzdUTJt8pxcoTQaloOA5rNO0zxdoyAzWjpNYU8n2Pf7so
4q/Jj9K/SCoKK1iCFpnLqfNyTs/bBQOtoxqNcFyzc661rSAIJD01bdobVn/aDjne
Cx1qoIv2HriRO0xjuPa4ZKBESj7dNmOFzs7feNvHh4yNQuJICtv/V2MtGWrNVzoP
OuDvSYDrGLTkaEQbuilclxk6YOZ+8OUH30dVayAP8yk7Bk8y8P+54Q1trP7swIYI
YGi/LvTtaR+228Omn5U4qeHECgj+cl44C1K6t7C7hsHUjwagF2eVl/EZ2CUzLP2e
xHtCQ+AF//uMBAeukOF+HAIhfJcCUO52Nv+64KK+Zx3fkZ2LlI8FVXEnQVPYwk2I
3L8KAnnicPykTkmnNsor/mg0tnVpVhwB8A9DEyWcCy4k9WaJPb7MUGRRXzMOJdBd
y5xZK3pL6L8OhWHKnOPB7GyeCCR3cZV4PzaNKsO/C7oHyODovv5K+DccwDNsHI47
YWZ2TjcUOIhzm/CxQG9Wlw5KJRs5gHrZdLPwpaj395jgS7J+jMXKepexP/6HNlHT
p0HjRQfNteAg/kS2TN7rTDnJYZM5th+2wfU6s2GC/nzk/oeSA363aCiTuLBF2Z/G
jpGE6oXgAZH56ftJk8c/tZenK5nqyPGfUJ3PAlyb2LaboNNhI9KnlCcIzT5SVzU+
SYumP6qF4jJqPos7OwrhxHRjGsmdvYMIHDWkcHV6RRVJOScDziqA+jOyF0DeoA6n
6Xs5vIiMOacgbe2bqNdPYmUE44QoP2le5mKUr5r/GwaMCGGoUfiut8Ltbi8PCyA6
yls+5WMmIqw+KJ8hYRhSJ2P+y+MGIXz+WkUjMSld1bqE1Y16t/vfbil9GmLZBY2A
ICHwW4wFVu1pLlQs93nNJ/irKgx30OHuwerxcLarNNqNtXe3j/evllUQutN0/tU1
FLCTudjQJsrHjNoAjTmSI/l9bJEMOjVYA1Bp5v3ypXggMhGJzRChldhCI7clSNBF
cGfPbmeZ6XlkJmORCo0ILZkelttM2KrIFbDJJwUW7tYYjPfUup7XIi0ViEylA7u9
N2V7CbaVPZfmg3Qtcoj7gRgNb9ke/DQvX9BK/VCbrYajllRhJYfbInfjDNtXEy4N
WIB5p5YqlPS5SJ6yOf/1E9Td9CjZENog1HxTF3AwdMcC9FP22I7ZHB+UsCoX4Dnx
WUxC16ARxQSDEK1olkcY2XkqOx7GroGjNRf3CTtWZe9AWbODBMgfHTmNYcXndLZz
3jykL9nG/1UfnJ3P2vh6ctFBjCNEc37FHkTPTkSts/pXJBtHnfrKUE2w4GtXyavn
cbjvqJ+x+d3Xa/CipegdL2FOVgNLT+Pz7vEqmUjtP3bBL7L0rTciRb18J5aQkOp5
8rXi7CoS1o5fYx5O8CC9qzM3k2RO+zITkvnUcugbrMKS+fDtE382IpJxPT/ZpBKb
044dlkIXg/jpx3Op0OYKbwUdOKANiGXjJsHMtGQyrs+b5nJ8nk7FKJiu0Z509VOW
nJ2H698O+0FWyLM3j9i35Yrty4qUYYo/TeYeDqkvRJZ9YcMw2LzMqfIlMmP+wdbU
PX6jQyyoshpm58gkMoQ/NK+dCOUhu8on9O0+0a5VoxoqYYTFF5Kl7Uyd9t5VcVot
NnLDbjdvkW47uccEECM6NyV0t8SPTJ4tuUck3JflUBQ7amvzC8V7fsD9/881yrfV
ya9dEOn7rYB+3kVbE48U4yWIWMcT/ZHsU6rJr9qllA3yzOKBKLFCvfeSI6PfVZiV
HlOlxp52Gxl+VRcM2LiqHfwmveg3/82oH3kPexLYJRhKtrRFyOMx1ikMNJWDKOQK
nGICSeQrhWgvSn7ZXn7kXirxn1/VGuEj5DiSNsO7WTbL9pDsaa6vjt9IEmCIZr2w
9s3qMhHab53KJoBeKbvG05+ET7wHMtcXC45OStCxol0aTBKXPmr79SPd45ZYgim+
8ORv0oO0bRLpgwbSgOO8qO4H0OvVAIiJgLmFsoVJIiYCbW/GRbMHsNrqkz0H2p1d
vclG0S/e4cwLfatXTKGZwosjREpqzhcPcop+B1R2di9zIT7naL+rPlFprsekbue5
gk2xwx1SJsyGubgZKZnVuGqwHidLgFarQJqjueS3iHZ1xL4d/5RE+zuaiCtVRBmX
NoAW4hh8HQ1Mbh5h6EKQiGGYtyAwZ+cexX20ULTMjevBrxd/h5tarFztIOm6AN03
Rsyw8flrQpVaZt32Sxbz71bEeOPNODsWih/Ov77efoD4GOo7oUQUdXHpW52rlkzG
CIu8lkjPUcMOh0LpUSgPk/4/5X7kkmqvwySCflNpBePox69czLSgOGiVmpbin4aT
tq0N8a0uOvqrK6qy9FGGgrGpXirHU6wF877ynOde+mD6i/w35VaceUryx62LdPp+
n/yTGmA0/dA4xJGqjdcRYv9gyj8Z4X1vf8V92+1r/QiPrgsfEgqJsyt/virABJY2
s7Mm+qNUFIlv+A8Grt+FE0pS8FRjJ6gj12g8AXoXEK8FRtDAzN1b615lFUBzaNeP
d3IeoNCkF+JDBYUNrHiYzza7mwXsY34b1bsuslL6EJPwa+sjoXZSjBIpSn89uvfk
/cRldhGuc/kcUjkBrLpH5AL4gr9IGmn7v9cKOCW733D0NHswGh3HCkFnwJP9+DyM
Rt+Uss+zV2CJqITFQfwGlRxS7++VyGycnDsADx01uuOceu95baBE8tr8N7+KqGSY
dWZoAVwmwS8yNH8HYbEeg4i8/Qv/FASWxR9YVQpiIYhJaKEe4Y1bSLjICCP9cC0I
kvuSNESxQYSzQj7zsNz/nIoy1/8aet8k6JnRTgIV0fItOZtdQDTctSQsZTq/qcVY
eV6iPzXdEc7PdkviUGmTohDdBpVqdhjuv/WuAX4Hvqo3G7vQiomMZfZi/bTlVHC1
VldvymqD86r0Fvvj1dtC5BsMnRnw0HwR5bcHZCpubqIO1J+Qhs/FVEdDCf10jpwl
CRqm+XwDgSG4FvKp2JiQW02fxJANcOb0+V2tK4JEqDj/CXW89AY3+XK10vyi1fSQ
VsUWoiLC6CMm+jBrGULEjdBvJLDodIPy5qMZUGQmSuxest8YqRyssnkabNfPUJMJ
vtfLutX41koqCxjMLKoraR76BivsIlq+h3nkRfjJ17DZKNdDHLtJazNSIZCuY2ej
nAUY1zUXk76gwuUIbsSqFh+mfS4PBxTU7kXrsuFS7PTtmC5pxnL+krDZqEyYjHKK
bL8egRdA8YWI8/Ow5wT7BWSZakxwDUwjotTRxZnLRxO/Z9G5wEbf+zh3L6PKTfa/
fxsn6asiuZ7ihpgUhbk/K3+C4JMZpU0+Ziqwy2AZN0KtJ723cquOYHd0ppoRLKuh
5jqgoo+er0pgjkVdY11fsElE4WT31F77L8AHyTvCIwExKihVCmUuklXm66R32x/q
Dp2M01YiucRjtbGJa8MGiXJ8TC/R5otRxAoym523wcQAooBxkiOiqt1PJYijee+R
23ieGkUcFBCQKhOoLaOK4K2LI/HE2p/ueGrpPR0WGm32jJa7E2KeAMAl5Zhs2W1u
FAm4adD+3hBHuZ7FIqXcptVxbnPIo7wJ1bihaiBQmLFtbyt6s1ogKHKQcWwlOF+h
rJuGSsphPQvWSmvOS1Kf2u+rUqv42/4H+a1L6xd4h7lWxO3/J8KS0orn57wOvhrM
B9VumJ+1sojLp/j57w+N4x7VmSJwrYYvd8IFcXW+NNeLjAFj58/Z4Ts2gTKh1bLM
goz31noPMoHjPS4WcPQG7Ku6mRFgiWxjxAAP6a7qhWd7hKRNpRB1oPu+HP1+O/fi
arJ7xUbhdr4YZ/8qoatB+nOnyEAArZrmF7GITMAU36ET0R+HytNEpPntSRQAPxm6
VkmiXPg7wb0L/MPPqF8tqdWRjWpxzuRg6XXtBpLRJu1z35wYAabBty/NuCFAnW/9
NdA/Ih2O3BtochkxsXlT0QPPCpYoLXBQoNloxOYFtEEE8OFOd43C+yW3QHuHtOZf
LZdZMazGUAqflGXd3Mi19vECBGsnRgansYKpStqgWiMZbVfGCVKK6f1Y4pbZi70m
yARRsIy/2V36MpM9t0KV9dbYT1sx3FE14n2nb0xtRPhzZYsx9AVOw3fSrXYpwZSh
jM0mXO7+MSmzZEFwyDAHrRbIYUKUt9e+iMzn4kB5LxFPfZcRXUe329QPpY5GfMMX
mImdmUlFKBoifSGayOhVW97pE2mjlki5oTm7955BY//tAgAL4QkizCuHIsBdHwcp
4PkiyIPqtc/J0Qq/wtzjkgcR5m8WKzE1pJU+0EKqRe3sY/4gc1Dy37YbMVnlR2b8
ZvcQGwsWHhSzy4bgrTHYARFrvCHE68vAB9iIeD/We5+oQWuSx55ycC6Ssxa0Gjsb
1qXuaaKmuNug5CXlpOMC65a2sml8fl29dZj9870m1oVfldUtu+hjqKJnRlnPrL7Z
RqslE1/8pg9abv3KMijG1KVg1vi0lS44qbmPvmGTu6rWLEGt28elLgOAlwvLbuBV
bU/1J1pZhU5ksjUME4WoaLXDGkRCvouSDmiKjTjWEEhkLHVXLfWzlQJNZ3hie2Bu
JipEYqDlzWlptJK1OfrxNHKja0LusL+5lqh2d+kUNdoBcGGBHIPUSEVeToucZeZm
apOJypU5vEBaOdH2tfrsnFpVlT+2S2+rLA24dPFnZ/i6ThNhMQKPstgzz0t6zBrZ
PibVE5oko9/aW4szn6K7rBHxyLlo7lZhGSoryHZvp1CJrxuLcBSOq6ZAGHGriYU+
1EmmQrS40SQFzk6NqQqNgZ9VJGStICcDOt1HLf29V/ew2BOJI2dOOF1rt+K28pI0
7qm3uaGL2j90+6KnWJA0tGConoMyWz18dHCvNUCbmEMTbh+3FJ2TWNOnJfn6bczr
vBbVntcco+fhq2MYlEuPUtyiNdpXPK21aFbGAMvp9t/z9HZ1XtYQsbzG44przZ+5
W/OpRl9+nb3dKKJ+Wlt2a3v2vU/R4cjfq7nKtPYkFMhUpAMU7cQCOgOu8UklUGvO
LR2ytyE27AQu77BoxxWwjslYeqXWmgusja1jlfIld7WRqF5zdAz0RmxgcNKvIIaZ
AFEHXcaCFKwDDqPpuNPj0QosnKf98nVkUF02X9HSsTtsdJX2KRPEC1FnSYgSXhQc
7mO6s0bBGy4I4MbccfuNeW29/RZpuHr7+8+V7kmeZcNDpDafw1lzGtVBbVuRzdMJ
ZwWsDUwkicLm08CJoCb9svE6mrjXWZBzMg3+AUVHmB6Mh8aoLYhVQ13JFZVEBLNe
6LyROQPuiAVNfV11gqMB/IQ2eBCSYZNUGa5BKhmq8JpfGvYhLa57WkO7gdd33H9U
/PDrbYBA77W7mQ6OvC6icJQEHpfGm7Mg1CgCjuWtdQfDW3p8k9uyHusUJTQlqxhh
xwQfX2uptxQqneL4/9v85wKEUUIyQfygIQ0nPOMhl4abDE2wlzaFXxB8pdj1b8RI
88QtUEnCt7PS4dcmukDZo7U2S4U4gaEzhf9PtHoqeyYMneuJ9pbW6U8J9LK2D89U
uXhc4J6YWq7vVZPlvjLg5bLfiU6DYgDXcHRVC9t/Xk8mdSR7N0INTKLQuHaRDE4Z
hmeMVaIP7xfAlqzKSfYQ+Kajpa31VZ/U+lN9zN4q9KCUTe5GD3t8M0bNQo7WgYkw
vW7TWEiZbh3mqrUtkMf8DXv7Ck53jKOvlcJjsOE3cCnKFpHNdvOS1ieyi2SFq3gZ
7kJ9qwYjdItylEdm0/zgS6sBEegyeZ1OzVqkqtqe60YulZOQdWtx9tAUDpQzBxU6
KtAPZcPWSq/2B8iBvkiiWazSe/ce7OAFWQnJ9qmnPrLPN6n2cr/TLBd1jnK/mW0t
iCi//4bZjyPUDF2ab2oHePSeGeYI/PnCgYkO8xdn/MNqTTGdAD+mBNTNduT71NlM
IM3dExNI1axL1uV7CAP6DY+Cm0ST+F1G0CAEMSa93ji3OCCyQU1/e6VCTlOIKQiy
l0HSvlmoKII+1ijV611blbbNtBktoFwh0uQRNrgo8ajgCQW1EUWADtmwAFGwB0wW
9MSTO/5RMdbPPN0v6y8wWV5784ygiMS/Y0wZJBXE1nQEeZaLG2jRT5GbS5f9ZJvQ
VZXsSDii4o2JRMPOtH5KFBLMMex3shj/138pPstUMcGxJBhgTrvwNOhtSiXBl4m0
mw9leFNDTVPZII7ZidEr3Y4LDcE5AHi9QUxDKCYXdwYKj3TU5aYkYsb0OYRsYGkY
I84G+YVpB6t+kyH66iiQLwIJ89zLsV5VaJOG5QKwne3e/7fjdPtdrqpl+yA7nbaR
ky+gN9JlnJlmS2CkQpGYKYSGeYf3ASWo5+JGUfAv7KNJzwSMY3bVsp0ThO/AJM3y
8aKjF3DCrKOPkShM6Qwv73zo2mQIr4u98lE8LsVJv4ECdjEHl64p3p/jp2Z8IwjU
TIA9BMLp5pzKdKMwdY/nhdlQ1T3lpbXqfMkZ3qNNJ6SnfOtDOgmOT9z8++q93afA
fi7mxINYTC8Z3cRCTm8if2lhu4Ysap1hYE6LGlUUd8Cvd6rOTeFFi/bLeMnv7coQ
gv9vJ9E5p4cCC86HZ0U9edRkcQBtUCwqhlUja39vrpWq38h7wPOjA0EVz8R2VfTc
jKlRo3iXIMzQWvFWgzj1I5z6YGAod/6uR6bH5kM3zsr/+mvVjDDTS7WZxo/q9V0L
VQ05B6t3xEB9EssIiunK81kU1TaBTUITVN8n/DsDlSkS1RAwL25ByNgcnBB/zOKs
rhiUZvEZtvZSXeL+WHN4e4YuI0tcxs54zoV5lbeB4BR5YpDuoAC+ab0FjePDV/IX
Xq6KoqiYynfEE0wy/ybpVhoM3j6psjrsUmgNCkZvgSnx1Fd1F9kS84UAW6eH396D
ByYM617naoS6BsNb1XFx47mJj4E4lcWjzRpKcOf64b9GjIC3l/QpNgY72lbvuaRu
ZPD3dFCm/8iJEe3dtQgWojMb57MZ8iUfS3VOS0fgiSwWQI1JM9d6cEcBu5/QxB0a
9tN79JdbbhC76X0Ijw+y3iHLv9fUAVD/UZPChuUd1zNMCegbgNPWX+/X6oFcVr2f
k8x7Z1U3ZGKJliLNjiHOG96tfrik65qjzpGnaznUaanIQsHeFLvUiCRH2LQab2Cq
/8TBDP+tm2NpJxGxBxHoDCa2CpJecXCZvCOoyLDHtv5bA68k2fYKmHUdS2nUPd0Q
yNrUgt1tCq9Iy1C4/kig3rKEfrhWM0cL53nQMQKLKf7qe+LdFD7hrW7ychRXyxGm
KBrS7ndaKL/87KqqzekzDqVnvc4k8DYL6lh/AFnae2C19VYsUr0K3hGw3vdm04b3
d8URUkge/ShiDvBcvxU7zz/WD4LX15UQSZIj0R8ruTKlpxdVVDYSW6kilhwPPmrt
sn+ZygGjlo9Dadt9PzYxZdu3C9hfK/+aSVacFJJHqjIB7sz2ieYeNKIVHKrF0/ek
XEn/Llp6Rd9hj+IuAKaXkhDPykm2Gb6Fac6UV9Z1drPw7NfMGkA9VzV7c4HAPAN2
ikhgzY7KhQ18Ay0q45hOdcLakdupeyOBNjDSzsUClB/MGF9A/ROrZgI1s0pOPzv/
mM4q686Bwy5lGWshhxH5ZJdlRl2IGxK8NuH6xT5+3c+OSlbEu/voJ77/pa4KMQxq
Jujgkc8mJJHn8UF58g6Eq4wty0yf4XrRIYDFXyD8cuosqLVM3CI6kn4mi1VQJBJE
hR5pJ142lHu2TIIcp63V050dVaDPAvFtDlt3aaJ1+axJeqODfGLeEtuLn30JnX0n
mNyDVYjg17R2aseYsxO97LO181GXq1xgMPO63ITs+RhGXA1qhd9cvd1g/aYGqDYm
nNMeo3yz2Ck+BqyGu6t3/bzJidg/fivC1R4iq8XAw+MuUvAKaQzYSwOrrnri/VAV
Bk/kvBYXBgAphJY4XIbnqKlTgyPBwCHNm0nEAMeoRzlwHfbjI4+xGfXvrpDavXBN
U8jhNj/IeutILbxIOGnG/hixf4S7gUymuXxJCo2BKSzFXeuT0eWofZQgF4Ymc5++
GDqPxQwpUYNz5w3sUGV71cVLOc6Qr34iOXFMlSkTXPkIrrHijf8HSeVC4k7Sb6lO
KFegbf5fRHmppgczr9PDMMFmGXdWQIKhOeK++u4fa5b/GfkMD8RUVNdi/iBmr892
vrnwXHGCoj74ip2ZI3YWbBuGfAaFIvLvCYU1liA5tHLy6JaRIcYqFmJVSWSeQ3qL
HMM9/JNaNQECP6XmBMlfGj1LI2Sfddg1YQz3ka5H48cOHtBZf41Ltl1Du0Wd8E9v
QnMcHjuz8hdnLIF3HdQI/UyYYd/CmqsPhBK7M6W0PNq/wgkTo33M/NwAhTJv1WJT
ynKMcZC8sHjfenLuJ1EwosSKo5K045d0mnktQHvn2xw7d2e0mggf7tb0bUVmo6Sd
qFCEGsoSN25h+IauhAm9ImS3DC0oXpMf6/6g4cZ7xT1U3DqYCZCC9HVMjpBiillZ
7OP9mp4ldT5bIECHEqv4x5PpRX7IKfZoP5txSO83J86qD/9luyc2bMVYBTOp3XUN
Pcp4LQaZUpVx4rRvgdvAPT0kUg5R/ReXmw+LCzfunAt5IAWxzDYz2uw3zbjJSnIr
aWbubpAWtbU7UVnaFdsF8VrD5kKHKrTUx2XN2nYkvebwmEPNcewtoOx7pDXg5nNU
F+5muXWJFKpdeGsAEnStCNqI+5UETieY0fb4cDdmdjJWp2Y4q/VoL9w2VAs85SXf
VT2eGZw1FchRg9OPvugjt7n3l4/lVFPqbFAIA5rl7MQ+BuEcBYYl0rKHsJFjXcf2
2uFJPmcXG+/PvqxDPUKx1u7ROicViuJgt8vJiA6+FfjYYQ3tk7JKTt1XiRV4KhO3
L63M7nSuF672QJ88ceLERz53Q3+ODHkv8+taFJKS6tapcErxz4QdTy25MEMSZxKA
JBnmfpxSCFEN5aKicDRB/dGMMNUWpSKZ52wdrglpHmWXDcgEgquUWGKvk5Mjor8v
qftT/u04VvDO5g++mDaPJqRMsWfNCoJKX8tWhO9rVsE2qCAZCdl4nLWNPJzD4k2/
KGpvD4DtWsxQ/e3ym4q9oFoagwBZ5oGX9Pd8QmRt2f5Fi5fDaJkC6ZQWxHNyt5Lu
rfx2dv4wFAsq6VxnsR3FnWRnaGfDQdhjIlpHZNGzWUsHfHIn6nsdfxgliu7gIAjU
Pl4OUxPGU6ZQa0no2aA1nKGee8fg+89mbzAHWMG+Ynf6DjGMZ2PrO8VHCAZZ4Scn
cRK926kiIVwk1Kank35kShAYMZxOdeC44apD0qn3mAzqj7aFWpTiHww/g/w4hpf6
DSUxvCtTbGc/Btpk90NuXuqKBkx0adpznysKmhsoPOK4C/c7bNkEy9e9W70R/k2o
K6mhwcBU5iT4FKQNfnlL6Ht5gpiKnk5224Xxy02usrKAA2L7bzN4D7OUXSRkanC7
6/EtVFS4cLQvWmS+cDU3XGW5Dlgy3cqiZUF4AYOs1Q1t59EZV0Kx7wrUt0IGDFZV
cachOq0Sft8lmoroGSRO1TTl8f7C+dBLXwiqPRW06ETXjjK3Qg8dlEBWF28Kfpkq
3cbi/SASK+s/DMdlo8MGrxZowLnXhnmAyWRR5axH8NMTvuyqJBVIX8mWYmmB9I1m
QkfzSJOeMVagCe9I+ziDesawiVSQHI6AGKxGMQvkBOpAlU0txAiv9PkYjvvTWx2b
BZ6QlCNke1vF1Uga6hRPPESYJFVb/HeYPFOfBRlozAaH80yEc7eqpqn78YscCAZs
zdTslBgsJzCi0sSVU4lT22/wykg4wmE4mUZNwWSI2RwVr0w6fY3Zt4M+60rCnS8w
y5V4UrHzH0t5tHJ9Wr8/2E3VzMieIniC4AZ2yBuyxxoDcCeac3nqrzYvFiMlKZHH
GHJjVAWnvTP/vous+ULxh4Dhlqj8RvV3CFqUpvc/qXpD9Vd1KJKtzAiqNltTkcZe
x1nvM/SIGwaPm5UexcL8AimySsnhGAOLfJ+SeSViyGgREhW+ONqooA0jzqyO1UIv
cmpjkY8gcETfPQaCRD2aa/6IbERPqDsvST3TA43/a5sreqhjMZ07fkgjco3rOoqo
SS1KqFevAPAFNjcWAPZLOHoEImpsvBpH8YmP1OlPgPUt6G46iWkvcXdPuip3zEvH
BDYTQT7MLRHLpPc91rr7/IBkzeAbzS1rwKMLfLsusqRsb4KYMbXqiwl6MoqlKqS8
it8NYK/+C/Hm7ZupnbxfZgRzPtgpWZaxiPNcIUjHYfjxfc0ev5ZboG/jChqO9P5S
GiNSVFFwQvb9cHGmBUsqYFoKKnFALZBY+6R1arsAIbuts5rekWTtyjSuyVFuSund
YaOZ3airOyDHpSncf/DNr9DEUcicMP7ciUyZWyLAT6d9OuNYStSRkTk077yq5mw9
CLEvbAgpxXKANP7JFnAMqKnuHU8b96U+WR4dZA6mYlFivFlpv0XOvkF+6RDgfwVp
dTu6G7WNoFX2UScD8PTsrQomoWpvl5wJIvajnMZrP1WuVW4b0E8shQdCy6jVQdoO
iZvicq1RutCANmnsohCvA7fxU/EOCLjNNzOPO2NjfkWaFzV/9dfeQ/vmkOcIcePN
RER7PszQRTeUpe3qLFck9JJS8KqrSQTQIuF63t+W80j6U5NF1J2nxNhwJ8RHy3zP
gOEhkv2RvZNXQXXn2HM2RZsRjWry4Fczkuc611eF+YCkhROMguliHOY4CAmK6dC9
wSSqWTOEm7hHsnkX2kWF24cP44Mx9Aujkng9XPyhsbyZOtzRHgmZKl3trQAp7Tao
0+WTfNmQxOi7dzMGoELLLcacx17CCC7T32UFbTs8ul+3MzDn4Nu3vEVmFy2nsgMA
xksDjzlkrCrtdVvl2BDuedcXhRqWVXvlyedQWqAruofcUA7jQHM6sqqzVjVGNy4P
9+CP5QpuerCJk6iaZPigofmXZqivAK4dWAd+tQeZM7UEpMEd1gRih4LgBWJSbbV1
nR+OhocJvdheKoMvwKETv0uVbYpyJV6uO1jUgodW+YFjPogMFxpE8/c9N2GuUOwO
vWTkGFx+s3ahwgximDp2CHOEqGQwSWZxm8OwSAqjYWHyN6kwuVzPuk9I2wqidV0P
B6XfUYUl5hKnNac2m/5pjyUHXVLNitH8jTCsGPPQp3qRtiSvAbzXRMhF6o0IMAW0
BInrMT6cVUazKKeEyg4gQLk4OHXbqHQG1k3+ZAvbf3o95X2yNXlPDzjD77vBaaG5
5rTZ4Z4y4WSlMfKIPihNPzy1RXBSZBynOrZVNngzBI5SH5H2CLpQmIKE3KBD6qVH
ivsF4bEjAciSKBXojurEwf/pZ0jizj4lIziuKI/OZVXeFZ+50l9FSFKKRI5tEpKC
ugKJilfuamME99+GMSiYxX/OLDFf+IUH2X00TwHssOOTNXVZ13FIIh122gNGcYCn
sSkqBpG4IgeJCneiSBhWurad6k3rrbeY+14jeeElUfh5jOG+9FHgYmgPtukmXelz
PesUke2+HJi2GYnBpfHr0ovSUsj2PHelNrzhnmePFjKW63jKzqrG6NG10MfLlF1C
8TrlH5D1P/0uYeJwqHHk2Khcv7SK4gaBwLYSzK/MAhX4wqr8yp3EjnMOGcWwIuwq
5KoBKbW/d5afDEmfjQZeYvQLoewE3Ptw2pYiFPxi/d7eYhCDoLJp2fM1P9KMT/ey
CieYVmANDKN4R6zAmvbcRnGVpDTmam1nCCIkN701mPgH/hpudz01LQ5DyRrk+WFA
K/RcVpRmZkffLGkybgBmUNL81i+V/WUersHzlUQo9MrUtiEYDjrb10MdXnv6X7aQ
O8YqS2otM3pXi39C9pQsHTBaXpYW5yTnVKOpK8vlbeS79KgHYf/lpsrDOzmX6ws0
FHIhEmkMD/2ASZxtIqrdJ5Km7oANk6n6joXjlV6geug7VccOw0w5Ncs3EIFM71SB
U6RM/9eUwO+5x1GtvXh4oqZrbldDgBHPc3i90/IeTh8HUm6ZDFIZsbKsOEu7yOle
1BXNzBmycZznyXCaNPsX/lQIfM9igbZiWrofIHS55/MQPOYxQFh1fRoRdCZX5Jcy
mxVr6ZvhUf03u6yTfB86MKAmar/YTpiKQYRgWWx+K1CmPQP0CgQ8pyUigziv1kRZ
DKl2xhnWdJaJXBvDM1onDQV/aTAm/4S1NQ9E3lHa3ZX26XTCktEYVfVJcA9mPlCo
mMR9U4CjcgM9IviM3S42VGf3kc2b2RrnFF3B+i2gKh6aujxZn17xGA1LDZU8cn8p
fczIIYZLL2Mi79ca2XmVW7dp8xOEUWTpJusZKBvWKSSa/zR9cPjNnaljkB+wXiJ3
gDQ/q6ogZf3AWQL3gzbmoQQQz377aCYDtXB3VON99HNaaW3AnDu+9ZoCF0lL9TEG
Dc4Zjc0/td7mjrpIe9LJ6UFzPB0SrTh6dFwg6ZMehmBA2fx8Cxtp84ZqpT1uMB7f
yimkxzazEBBpX1ZMsMjYgdI1eIpM3pTkJclIk0C2a4qsAeNWWGx+jcK1GgiGp7va
lFrlNHPtV916ZMPd495zZ94kNejf1Q25O+QqF0AvUFBuYni+o3fhn+zK9wcJJqd3
4Dor5Dw0HPDnOCrJwNl77hz1atn6UlGJllK7JdA3yvmYt7aE14DeePqK3pHbslZk
sF5SeBSe6yhG36EDKOIABV1LQuSmWF3EGGeRUlW20B79uKgiDfb5XjSGt9C1kqWQ
5MNuHW48VC3oTipe8Nbf9FWuDirWtCERPj0CR2BvmrR+xFCr96F7kTVpAOTGpxAa
8Cju6OD9LYGyBAi7YEie9dLaGUF/CzJ2333XMzH/tQU=
`pragma protect end_protected
