// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OdAGaRBTzzk+innLSWrlBJavjF1QEF1ZhDC1ptKxjD5jDPDVI3Q8fbsR8oDuZ06A
5ywbX4KPcAJsroMGeCo4sTPZc7jIWbnsK+mtcDii/kVKe9DDL7woauUIH74L5/jQ
tafVwvJSykx/112hFMH9lniKO/epERETMYouu9D3ShM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
8bIdeOOZ23/aEeUMgE3G+DFMuTekHzIJeDvsme2WW0rHSOW5Krcy3SBsqynztroP
eXwsiBUUw2KZgeFCDnnGrRh/wzcAq4CGNIr1yvtb7BHYLJrmiooGwocug9r1FORi
z45lHjkmL+1FTBrYk44hNNNxjYY5JMrEWYVz9b9d6oQkkNz/HS3f/HsPC738DryX
DdVGbGNdNgT55Mp4LAlPyEx75j0hWEAcYUD/VaYhKdYWG+E6GYaLbWX0Vu7iPpJl
0Nhqq78Ss7FA2xJ/tY2xeGg2bCsHuHDjqVDUiAj685pQs4FUag0j01+jSSfYFzBi
bfgEKRpjd8EcY6dy585lyfKQTvcvcJyjqVooomZfhz+c06QAQQkH0e5DSULWZBL6
hRF68XXEXwi/8TdblG7Lp1BIy8z4wDirOc7D6V1Ceav9/ZL8lU0r/5OB2hE44dqn
mgOTsvbxqAwAhDObOIUEmUzJQDWzmosbbO1SdFfDDVqw5uRl70Qoe874MiKSkYE5
AKmwW208EyQi2Oin2L+D4wu7sCDoRENPuCLEPF3pDxBRtbYo9MvaFq3sG4GcxvYq
5KMLU3MW9nJucJm/mwexosLJTylNMZ0eKL8hDtORASfxQ/wa/+nuSIR1bH56fHWC
bajnF1efL8cCIVO5EXxMplJRWa4GvoLwNrZKoMHdgZHgOrWqV/jq72Tq+DcSyz7y
tH5hZhNR73CNaq2lgva65PD1qI9FhCXsfLrqqbZeK02S46FsgqWyN2ieErP7QCbq
NLX/u9lMYjuddAJ/LlVvp3Jeyv2ViE7j3vsK7f1qEsfQBaAz5AfQXgatXGFWSCl/
Uj/z9OstwF2ZLrIZ3HjLHMIKdYWKKZUHsduWOifP1GFGOWADGgXndeRSevORUXHq
EvTyC1xJzRnliUpZcKqTctpTueDf8vw+djUUbpnfd7N9tuZaJdikwSC4J47saWGz
WWts2EgtDqe3YrqPcrPCp9Pkf3m6DT241WQhVhSHVlcXCjKbCmMmAhFvHxmr07OJ
IY0tsqZ3Yud6jLH6vXr+8MJiHvdwRl2u+RlPuvKnq/mkqN7+J4b9VeNHu9S+6uFo
6jYbCoDBtD3O7C1rVWT1rvSs4GWtMDQ16aGc+CsAG6wJY5kQqggxAh/l6s2WrqfP
fHzd61CPbOu3wDL0W8TWKFITVg2CPfSzRmy1D7RDcIkuNYdn2lIYZOOr6JDA4xno
svgroATYQIKuAdk1ZD+zmFTnkKQQ5OqcvnNtFleLZNgGNLBhXtfE6CdjJkv3oqgB
kV7CfRIEVT7G7+Wmev8ITBOgFEL7M9RSAx6XwS087c9JZJbgij1NKAUPIPhLmPbd
E5/PYlSf4tCPLzhoIhlb+XMzgMwu7pUxtsSeN2jIFAkQ8VYYC78MEMBUPnonRC2i
TJ9V00ZC49lUB9HshZ2PXmK/5slpKuc4J3kWeiOCNW4Aa+KPsAvKK38/dpjhjr8w
MxMuAzL258zhBQaK6Xp9mEIbFHH/Sm4x/+NFCR1wtR8s+V94ZB88OS7yucrfpIMD
5ilTYynksyAtabmXEA3U3hxEArrlw0qfD+ZJav0S7n2CHET3lWU835zY38s71kPK
HHhAQdLoOza14gRGXSt8a3O6oFCL9o4pCOgalzz+i6NRr51Zpda5gtUs+IVpWKCi
5Y4s/wk2rSQy74qLJtoCkVoW8kGULl/fAf/lw/7TKXRJ44j54aBIKNsxnNR9JAsf
qsaObtX2lQZrpnQ8k+Gd2kZQZ++S7nYWnfBuqxt+pxLuwdJzKsosu+FNaSvTDNRX
t7yIiQydozRoSXQ8+dTJ/ZBlbLLphvfnKPAs2mw8cOciU0BwVeN7Q5z2UBnbj0wk
mYw7P2Ru7NkFS5WGQ8KsnhnVfDB6B3BhEUD6btyIhHxi83w70GaZYw/HqAcfOwHo
52sbeKmJAmbNrDy++vA3JgCPnJSETkpIrAyNjC/1ZP2Zu1Z8pcI/2rBUnaZEHVcv
b+/VT2gl9nIcqV/sIaaR9Loi2T9nEP50EAmUU0U9UIF3s23UslvMmx/50l8+ImK9
4J02ixAKP3gFuOKiXIwYrdoyjjva9ZS27JBVLwocDpfB/CSBOGkRLZOC6nkR0qUe
AZdj9c8SmV6lQqypDop6Z9bJ1FxuH0VJeeIXhFohHyUN/T7qLUPe/HJeaqzo8RA6
lp2AaFFDP8v7PMZ+vd/jijee3OvRtcQz0qjcaGqbN1AlCgd5djCg4uAeOwg+y/Sz
cKICTKiwhq8X15s5mZJsx3DkCKkm8HBbRVpfqzwc3XzeADmvl+svBaAY+qLwLqZN
cKqtk4CmwkaekcMxIhIw+y4XmBEqqVovpBVNgG6HBPP0RgNtwYjsG4iYfHdEkLkD
Ro30Nw3KrxfnYOMIpcnl38RaV5EDWPCRBYxkyf3URSPAfDtVzYQMqvSXjQk7C934
12SQllhneBL4Jfr0ZOWifxkMGQmpe11VgYN52mGj6dKXhko1t8XlKjcn/Q8J4aDj
85F+v+1inLIf+LFRrVyvOI+nRnj6q1gV/kXBrDritcvhlp0R14Pp9YCfSWWFWWpV
+q6YZc/ijaYY69ApM3cz9ZriL6ZCRx9sngOMredBWakV5jM8s28T3WGZsH3Bs6Xy
pEgpuw1q2zrIxca/YCM5dn/g0AmeNcsCeui0OIj/NEmsjwZiisYfhUXqweNd1wQ8
vNziT8XI/wFJyw+JcVZFUdnLVCjcPwrapuprtG2Z7SBZrfODrbBX5ZtOu1JE0RMe
qWA/l9cQ+qR/ixNDLi2XsflLM+ituSyr460cPQubiubnd4dz97WhYGOrLyZd4P67
kCtwToZWhtC3LaSK8b6zMsDrlQXeuk0fopS127btlbKI+/zPONbuvyaDrMqAAoa3
xizPPQHJ5FxJ0Kr4xz97nFRmVcgDXhvnQM7FKC8YJlPBIyOMjXau1vVT2hjzah4T
mh/pP/GkTg631ZtXZEZeRNnlUhd2iUjxrOjak9oRMUH/rOraM5suGkZqHl7katWi
eiOGy28wNLKmLSogo45NiA3bdscDnhAYZYvsWso11HxVLWQlX3J4mFFCQzYACj58
LeCcVhkf9BJXm3c3H9fmPU/uYqS8/E9zcoQpzHXh+BPMTaDPQCs5M0a0EjJ8CcOI
O+u+J2lhzXTNP0z6DCNjoohp+V5o0ivV14UNp8WZRuPasHiD15WZaGO+AYXftwiz
onrmomgbcKIC1I1e9wmN/MySx1yXPov78uIE0wKn3/c429g1R8Xm4/SDlXsRBl63
tEXtsKHB95XBu9+kxkzNsUl1kKgTAPNRK6oCyO1y/EeFPe2QXY+2dHthWZQbySqa
uGnaDgrzaOQcdjKKzgtwe0Cwq+JCOeJb0kx6orzDukuhYumbew4uYBeCgBgUQrMC
A0b91Wlu0Hn+KBg8y0MtHb1Muz1JbLZpf+8lJ81elL2uFz4eWZ07TIm6DYYo7TrF
FNnc9O6ZdvWeZk4oHbaVEezvG/JOxgMxXS2adnwWVq0jkQsxA4tZSGrL15CjA8r8
7OtiwQ+m7j14kVnCv7mZWeY2hXHykMSWvpTkF4oLwmQpFqTzT0Qvlaar+ydT8R/i
omFRpnnlR23oHQqWwexjZ9/rVu2P8VsMeAHakLkwBjAzYrpLWp8r2Du9I4dWvuyp
KebEjlAMOfn1LU0HG/5rJApVHk7MJ1dWzR7IkG5vAVxsmRAzXl4BAjwM5XhOJPB8
qmWNxfKlZTV+IBlpxJ6/rdfBt4C5it0cOXVRvs8VWrB2oRLVNQUiFvC0xHlQ45AJ
qkjvt5LllDQHekFu7yz+evsUhQRSnz1DV9I1w9KlI8CqODL4uNZt4tJac+9jN+2z
Iptxu0F0Nm61oGBkTrJfA5PUmwrXGt9azsfqp2BehJpS+If0qAyOOzkkK5FbQ7cI
48dZ/G8S+niRwbk8Kp+tIIoBlbup0IHePExR2OQtYx7r9Pt27eMM8akuTs2oci76
B+JtyFxJCG0UGq70DTJvGExTtPJ5PQgdRTHat9p2ORXhAwlVB97cygMnqzxD1sPX
rRmitqKJCp2ab5bUJ6d1g+F0z+VVIOEs5TlGUQX5NlLM0TJyddTAu7+EWmirb22L
YXDe374NtR5+ZUDUuabIZobiyxhEdln8GaOoQXCGun6111dbIlZ7MHSc/uUI2+oD
KcyfJyWbTeGyc6HVOFs+RiZv8huTMDtozmlsoiZaUzkhBLGAp3uewTjXfSetlQKM
TQWAbnK8Biuzt3qhxwwNXZ9/ZLVHeBAhL8GWdZQKvHH81tZrkNq55Y/ES4chsEOV
9hrtuRvZDMRaevdH2X3ekRa0L0uEV+gn5Wlx1Pbet1xPB5aJ+PFKFyNNi1rKTw1h
ZhOrQHVHptr6ZXf1WRgdmkya94WNRhlb182Y4IKLnJuWv/dtKC092YJpVJV4SifC
z/ktSc2CoktBnSlLtm5PuVoMqqoZbUkQQ8OVy/Dd3W7kdYAcjOS9XY7tWfFCtwAG
ZFR46uKcwwA9EJhDvghoZuAZ5SkMh5mV6WJp3DHZMcncJPvw+hQ8USRTSitdW06d
R01qoMMlPvHgWhzze62k42a5OzpacYX4sWaIqvq4wRLdRnb7SH4Fggyg4oAHiZh1
y3qDaQe+YFRIrgXtaysdWmk5bLgR39Y7cdhWnRj+7CV2zbNIjiQaUICKqH1q7azv
EL2cRwB5vkjCMzUYRBzLoVPQlmgs1+KogoOMffrN7nedBj3xmqLoUWt64aWfilzd
bxoTepFzSy8aLLs3Mvr3MbLPYVyutBVKQ4fkoUCk1iWWIwinsuSynVMcSHMGKAEz
22ho1Olzn+3sFdVqZZuQgp10XMnY4aWgauq45WQbL0s9F3cfxM4eSlvNQD5VSyXg
NGcGPF/BFhPDCoCY6uAFFjUebak5wEwZSZCaTKCs7+B2pqNHSgSaDi0vvBsr9h7S
E6TImY3ER7rirqW3QjiLrpf35Va2TH39Nt2h0DZ4HGmcTGZxfjhyT3bFZ8HyRjcy
S9UnN5dzbaXK0g4pIeb+27gqhH3QUKvD/VZUq1kjwJan8aDyvGyQRFdPrfNLCPCR
39U9a41UX9nRYy+Gi7oiG9vtkhUa84YS5MV20PK7QfnO/ymf0mJqokVIrlEhoFt7
b7QbDsPIg3RgJ4WPDHykW4PFkt6Lqfs+xNM0aUPrwnLKzdKuDRA1nOB4JVAwEiE9
FtbDPrq2lpZDtBj2f21sKupLYNM5suEAWDRjz5d9Gtb1MKbbyRdeyN0MZCjagVB/
x6ospxgMR75l51/UAGkminU/oZ6SDbnaAfKXSFQS4dwVteJ0ImsTqsfxbcch+2Rq
3981F8CCTlncxx0UML+vaGLGSzi+8yYLVpLrFLvQTt05F/sA2GMnDFHKQYgy1eDI
t8m7d2oQf6dbILqPEjF6vUBHjnpAiPpui97vESjw1dHh5YAMkfa604Xezj5tRzbT
LBbCfJlj75pPcTGTuRUxcpnZrXLiuc/cV7vQ4tuDmL+tqER+DyIQq4ZUw5rlkzKe
WnUx7eG65BaoODUalPnp2h6BHkYELtszLiOLzndAS6vxlsEElpohDASBPlrdwcZL
bL/4y56cujPdxDzg0JuIv9eWDzhSdTpzrHvbmEhTBmMZLdnkxkFqh5komQG+qK5p
vxY0AHDUnLCg2yGBNmKIXFuJV7isF9fIMa09EmgtjpjowBdEDBrINI6xIw3WrMpm
APOzy263gebpsCY7l8olbm42M4mBvNrVVjbGm8LuE9SkZUIh2wZdXmonma2VJtin
LrK6lMsMnwQofvrRxw3cpnwW8vbVfhD1wpFoo8hBsi3+tTUtMTfuF3nXD190wfL0
XY/oBUmnjbMdRg5tGGU4Rw+rcjph/kHKuL2/baMQ+y84NJykJZn8yhPHZP48//HI
K0R5xkNrkkGE3Di0FVZ2EyFrDXvhw08aFIc7RDWFR0yOlAy45XwruO48HpLdvYD+
i1HpdYWLC+UAsNK5vod7d5POWMZ4lmFht7W6AYCk6uopRrKjLGDsgZl8BiHPeQrO
oqiDqAeWCs9GjP+XpRFaoPqmBxDEZl1TbvSOmWfqOnt51ZaUpngX/ckoR9AJkOE+
Uc72Y3vfHEICQ/olC+UEmVoGVVquiTVk8ir9+TUriNM4I5uOz0GicMZDTZf13Acq
dry4o9e4j8TqxCnk32N4xCv5fx6P1ph36ECksUFnP71NIpbuPmACPurbFkGdC4H/
IQY98dzZ8kRMBKYod3UGoO2g0QETLVHNFWnELTY1FwLZLso+LGvBVQMwj44IEkru
6dhlWd/IUAQDaq5SONwHDU5ri/L8/tFgYHAQrfGscqn8vVR5dcO/VMIDtcY+SatV
nB55OiAaoRcbOXU6tIGnSk/aJsZwM98urGLODC9DesmxPR+VrzY7e7KG6qjeuq9g
uj4Q/JUR6hRRPPppIiPdyjGknFBjUOyGJSKnf7SLDQ+gsaBFEiJJQOkSh6+5OsQy
AY1p4jPh0ZvnEUyA15HBs9YRm0Id0dWvtGo4Tj7P1kKvZ7tRcWQYH78eUELULF+Y
ntoOi0IjZ1cMzo7Z0zIYHkWyKJV+j4vm2+LvcDth70ov5g5roE9tz0Tve2/oD4ot
Kj6nu345ZHZ0g0gq7dGI5I3DAvd3Cu8h8SMwbriXWM3FhzqUZ0wQLNHDdGjJhxqC
wHK5AMjUMTyVCEilHboMQgSAGE3Dzq58bsEGSLyN0OSj2pLHGWyPKeQkPNW3HNqq
zlhJzWjJvwWQSvYslSdUtLQ1QCzQinCfxtkKIm0bKFEMXuZqZQijYaVN4tN8dwEu
YcCz4u+Pdg8NvdXrC0sS7U/t/AkV9GxXoUUSR4oSGNj8BgKa/XCpBUKDTAW1kzOc
0T6TP/g4m2r03zUXiqnF3TxKbnN2e2yQSp1hgJ1IRr5gsp07ECtoV9Pn7+5Bjbj4
jCnSSiqmzncspjHCDzuIg3LEL7Gk2BceVJgSBhs/NZdLsIaYvGOea7f+UOguTCy+
0sP1meJuTNUUYy9++D5zWT13NrF0D+9rSLIFArnh9NVYyzjyr2PoME+qzSj13aQW
Gg5mlCy4cIehTHk0/AVYIXGcG0l8pvTnYoagNlJpel4nwcV6GUPT/8g3mhtPrvVQ
+G0MjerQXVbbqVuMx4aeJuUxgD0Um+N1nTwkiUfqz8u+E5W9vZ1nWQNRGv2LwOIc
fsjIOFxbFYq6Ih/FqLif4C+LBWM2yCI/DdlpeKUos5C2BlDtFSySlEbD9NojnXq0
MbfvJUhiyvL6OJ3Li3IoJF9r4PjRqHDtwKDONAjOjnpfu5wRmDpKsap+PnFA7XVz
Llihpw6Cw1FG2JiIucePHcm30mdaDk1D5dVTs6GlhjgYfrEh3h4j6mSFQc/Eueiv
4QYYyYinMPU8J/0EezpqOKSBgr2+2AzzqfSFiQQuGpcEzfxcNjYe00yBkYTirA2V
06OXwv4KEv7+s+PLE/s8U2ZvXz8YkksN60qA2q7ydePak4sYGTeib1nYht/HPpoV
zseUrGzNhgSRlbO8AETAhw0EsNcRFojzAWxw2q/7FOf7nqrREibiWdwA9timQZ3X
yNizB4IoSJDaRQ8rb70zMeW/AgHskJ63sL3V7Zb+uWLvmTIsIlrrO7ZP7x5m1VL5
Kd6pGbURZn8boKTBmxa+LQcQRp99J5kRWz4ZW5Kq3dSn68uIBiLxzkN/4P5A1W/s
OpE2gKr1ip806ZM6pFep5MKqK2JQr7cUqYCIc9VJ4cPUxogqF9OTgNQjOil//TZ7
fVX28a+1D5TqWBD6yWZGW2kRdHLwThmdGwqwz+32Vis=
`pragma protect end_protected
