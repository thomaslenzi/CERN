// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YarES3aG+fMsqli08sa5gU+YULmWCw0fTu/gGGp2Tok0KgBtVcfbmN3T15z+FQOX
Zczf+ZErQNOD63IOO/7cGEbBScbQglFOTsGBy12+HpxZf20cDKc+Xuz+tXJHSE2l
i0z5jELSX5OBKucEDn7i/dyC3XVYwDegOUAFJZHvYHg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21904)
rEInXFIDNPXMLpOo8kIzeV8APqasFKbXHOIuAV+s6VlOv79lWB4Qb83reE1plgnl
ICtmWwMSGKXASdzV7bNsqnYMJZVUWffJkMtiMXIbabiejBgaM2zwbNIf59Yr/2wF
TBeOFD5IWuNkMOvbexoNbEXS+n5sdugyPx8uSVnXryj9V/O2fwNJGtEvzVjxuBs8
V2vXDBZ7jNq/oKRuAS4n7OUgCmQH3EzIn6/NnKK/uCtKGy+sA6Sb64N+5wmbCAoE
Yei/gyzGpNUJsip6KLo/g4AlxLaxqhNQFDNXVfp14r1iNUHYHwH5Y7uvy+oKNnVA
V87ca9LYKjE8fmo0Bq+u7+MTx5AD5w67wuQ785k+hswQwTJ00as+1Kv7oXHu451U
wYeg+RULZwJN9AYQH97tmfRMf11ay23miQf4IBLUDTewaCF4DIrJ42YkFwyj4iBy
4osXXAaDZu30cQpXWwXWRZx25Oy+wlZ5puKjdksAJQE7/+vKES2DDA/BBbqUmaSa
e4pyEnK71CFskQsZje13yIycUXoig0bh7Vph6raN4fmAv5nXj80g5LmtdE/SgKeG
9AmiMLkvfJbxqQ0aDD2C+eAeR5aBP1lvRBAMTjYiHjQLBGFeUW74bl1z8tjSC4IN
9rbAtW0LDJukeyDrwzEGPAPCEnubv4Ob6DekTXYqTjG1SzelF109Uwj3Dy0R1BoC
aw9lYvp0WA9Rn3N944fI31mdAeGMl71Xm58zOuu9SOiyB9rx21R+CBYcXq0zr1zB
IOKOL4dRCiqS/fCemJd1npnzWjl9HlFwdhN7d930XZLBLBpvtHaD2EBjaQlXq6Fx
RVjcIYJP9GWGfhNTdV9bTEQz0QSrDei1VFHlVU1fuPzI2LWk3APYK9PmC/F4Itlg
boUAln6lcp6fpSbX2RTIpG1tiTCD5W/GGgmopbLRavR5JLl+DdWLlxRikO/6f8kC
PnTBcaV9EawrsUxlUlVEHvXp1xZoug0sIPKDJhGdFj0wxvJ8UZrJjHGiNWTZCewx
wsh5K07DU8rN728OPeG+Q8Nfn/a/1dWJpes+UDjr+ErFkeuUrArTb6bVEYdCyStP
aVQs0RXN7z7cD3iB3qVEw+vC6u+O/tR1bcaEZ1JSarP0Mwu0IKdrxzpz1Mgu7RM4
5s2Z19mIu6wKoE3KKkvVw+Ln1dt4kYdAXQL9HdV5yJGqxBUOXXmG/Da9BhAUQ4hk
lZKCq6jw70Jks17Khm0liHP26Cnr2mtWIt0FRAjOkpBtRjmm9ZQE+HYR18fzlpEy
GYyVT0Xnyr1Xtndr1d7Jti8Rys6ZlE1a8zR/ieNEwpO0aOp7fDwNwoDvOzZneYzn
Cjxt/iWRTqU/qPT/ugWLhg+EPfVhTQvjl3xfFnkS2wuCgQ+qzrSY2SjFGCehiohP
uocjgzYCIosD7yd1tpxHY1kMVVETw4UhSnKLDK9SOEdVhPDKyKzIWw8R5lLmKCSV
qdxup2v/CzGWJbe+uLoYPNV77+kOMoHIgNZBg1T7vhsTrI5oBtk4zGHRuoSHk5ss
63c2W788TvbB5Q1w8VLSzQpFIC9CSgM9hsCFkLUPNTfqdhg+sjbQuXb6YTuVDeoV
KNxDph3Fngbc762gyqIenp30DpmKNIFHU2RLLQliLKpYVKDXsBO/yf1Ew/LIMTUz
PXPoYuH07gxoArmjaqQz2npCkDmenGZr6mTbzMtii9S55Eoj7nKWqfVXoR0BbSrR
odTnyqFLyO48MTQn8nRS5Ub8qXdA4qxtXBnacCsNr+8hIc8ruBy0IuKyiwE7IFwp
tavSskqHhRc9syIt/T8b6VKOx8CicaacE4c48aQaoxcCQeSC3tp+9ECWr8nq+n3W
7tXwHiCEDfkleOzqPE3BZif4Og7P7FvmGmhfDulMbXwYqV/V0ZFXt1cxrqFxf0B9
hleoee8NPhAMIP6Qy85j6At0Q3LScJH3eVnUvlzUjhzaVi0HCdrDboqE7HBqabrs
XYs5EhaQIZZ35w6GbiAyVzLb2/CLVfIbN4B61tWd5sgT7XRPGlCsC/8D6YTS+wyP
bR7o8EO3ble74s/4j5UzugC/cA4/uJTIpeSBD48xWb/ilRmGTrYJkrtH1e62n7pw
r2/cYQ+7SRCczAsWrMAdRWsJnaEu6hSMYsfPuFkdi+6wBwWILK16Ne6mE80fnNFG
vhoWqgtA0XPIa4iKRFIqXrhNFY4CXKfZa9Xnzf8qZFMn1m3I3ZxgBqqV4/PR4BWq
QbV75TMZJ0pLjxsNJxq9kuTcn8Xg3OxDItvqVRxDhFepPnkRfZVxSWSV4+aBg+gp
mDBFtmzFc+nODUBUj2PVgwE+VFK+71c0lhuHOfxFg9HNBDe2I3A0S3+WiIUNgVSf
x4awV3FtBnAl5CBeK6Y8BNMruiIbIiYaQuPVOGrqd61KB3hH7N6My3it5xn89u+s
OVUB0lxQemIZ/nmWmq8NxBEsjRG7e5zBOPg6OVB/FKOyb2qc7DL3ghkTwh54WMKd
jnOVuujNkz/56S2nfdU7sKWDunzPRuwLgRoH5+vFYKTMUHiK7Wr5TY2N7XJLW34P
h4BYRY2I6/MvOIuODcZkXjB5zRp0qYodfkH8WRXfhJKHfD1V0IRvSGP03O5ElzjC
gIT6vlGCeL7sF1t2RTG8ftBFwlb3ui8uM1ZxgCcynRQNYcuy01vwke9WAeaOjcew
cvK2ZZaxvZMc+2zQYSTY0bNUKO7Kw0YICrIjnDg6T9S4vurstCV4T+pfXPkL6YaP
05h9T8fu2PUSrxMZH/mFtSc/2PGghIKRTs7aMryrNeVpbi95cBSJMfh5s/b/kX71
tJ0VsUVAni1p4JSrGsqhizfokC3KBoHJulKxvSkcnPVEjHbXt2Hp10A80vRzJHj4
QVzKEdroeKbGAEp8wmIeTlDU788UaT9cKCn3fnig5r7wSuX0LAoqj5nVS5VZMkZ3
WJlILQth7z6Gp8EjJUyIHSfIXzZls38BGXiPzv4VNH4en6cJ1J5GzjyW9v3zkQ0g
drrWrSNhGlUaa5C9qOWdGAMv7z6ShEmdMbDdZ34fqtVXC8tyJIQ8AgYwrUJI018N
IGCZrrW0/jKYz8ZYUR+aDll+WolOiLoppwW6565oYAQC+S+5V+9lQAUgKz/YEsaA
BMh6vJxLO8wVsU6TQGtB2lIudRKCYgJmBf93wzGBu8rkrqpzyBlM8JfgBwGk/XqB
ZWQvA2jVBWq+KUC95NbUKAvB8Jt0MGKhSazcSlgk+ApRfSk5/TDohYdt8QVVHN32
rbkqxQUF2cM0lwcT+kZwtrio38CfWR35VKPLvUhSO9+ChrF8E7jZfHAZdufHMrAo
VyKEazcGWG6vDnfc3oR3qeU/hwqOZtrAfu/IDzA5J3f9cXwXFpttKOGJcvjXlnW6
QX5D8jjwfGFzkf4f1djMZwjCMZjmcoOSUQk3LVGvy0SNpuc+2ZbQgy4wu3/aQU/w
FL8ubJ5NC3NEdxKL+LYH35+e6ITULdzH7DJP1w6fx7svGljyrUAq3uoI5HpJexFe
UjVBO4A29Bc6wQqm85pCDzhqHiH0/iwuZ4XsSesB110hD+mk1JDvAdqMISkn/F2p
nTF4pBF16UpSl+Ltp72smvwkgzscgmaGOjQ5Ph3u1NsHZK9+q5S46b5Y1qWzJl0F
mCK6zWCxRZ7Jc/XeF7udp/GDYEavYpeJFawUwwagABQWpiFS0Z7Fj/4Fj3iE9zaV
H/j8NNIPxKsWgsCsl4OMWBTyu4rSwLuR8FygwVXO+c/NqYRiKs3IjA2WxyFBitt2
PPc4YRLajCsLHI8wmouWKNVXP6lMKw0+FDZNqLDy99EmV5js2aBa1qXuv8Im+j6E
CR13OAVQF1JhjuVikD6VwOqjeSXP6PXRII9owNV4WOMRq5ZkTfNe2WTu6q1lB2wR
pIeLrC2l+yvFO1BE6DIRsnS04U8KNS/moWn2m59Bgtco09YJ4GbbJj3R+9sexE2j
b+cX1XEQm+zPl+7WwOXV84mS9M0aH6Xbz7aRnqyAoU2xWOkbcUo4hNdgZOpwg4hH
pcd6/Qyxgt9fFyoe28i6uGs5EPNcdm+NmOYObZorBADgsNPwenqtAMuhib7axc09
K+ehjMg/UKSNsnv2G2cWZWlVQhPCOaaEXEZ1wuZZ672I2kXXXQ+UUfD0iyNMJIa/
KC9WAWc4nO07RBknKX/sh1l8mpF/ZTJalxYdgfICsUQx88iZjV2N4CLluhzmWAqb
QyG5w7ytPy4vTNr9qkJpl7tJ9jOoAo+LkYUpxT+Wh8qgjgqZZLcd1j4xrscdDg5y
+IWBmqUKcdOfOOMBaf5s/+aGNBOTD4bEQBjaQ9hQNnE1FtZ50crfe98i0kj4mIZR
RFSCggn1HInSng3O9fcPjBgf20eyqPF6LynCVek8efmJQDfXVlysTI+T5qzfd0br
V2lgA1nvBvvfPhlIen0N3Rn0cXGtZe34QQQ4ad3S1QhX3MPaRwGN/s+Y77jBqRub
axO7UgfOUDrT4AlWhwEn2h7qCQzYvgLLmBTdKdsQLyJCDnGV9YcLbYQy9YbkiuaO
iQUiVXBzgacc6gQEQNMbkysCBbH6JL6zkd58lYaOcTPDcngvWKDjEsxqzDPmD9Ie
DZLXoT4GePUvljbisV2A5+74G1URdddnmfHHx16U37ek76mybAVB2dfEnxRmJwSP
mQ0epdpPaJ3vwzGlHzSnGTmMVLG+zjmS/vr4Ty13aa7pBk1Or7rWUXLdVHUaY/4Y
l3mGbq80Ya143R/9EhJRzpkDuwBHRc5KipSvchFzWAu4L0Yw9+LZ35+WbcxB4zo3
WNnblXNsHxOQFDYQdEI4rJxLQUJw/gXHwein7JXfxVZ2W7Sa/in6eWbceZMOGgwA
3t8HlWfribaT47IZ9MJVACRRYMcyUY8HkH15XQky5PDlHJjEOycn+XIaPHo75IgA
yJROgWVtp04N1fbwWs56gyAWwNPS2/kNnDbB/+5ZPeJhgKqik3e0AzZHS7Tne3Ux
5/nxHMBVq4phveHyChoCmC/KfWzSbHBal3Su7A4LK+WJ4OZ1AZ9zgapCbWEkWbES
iE5UJjBTDPAtkFJn2UGBwLXOhvkyByx6YRvGLOeS0iX+MulUrhcjmGERgADoefdf
+ksHYuKyLCJdhYfixUQQaRpCTi6m/fplQaBCIi/RXWaBSidkKlm8saYyE6oPE/9d
XFNGAeXSUAIagxnL+3CEOXeV6Z52thWks7KJXkuA9th08RDvmpNd29VvbzucoCVx
6WN2BzusRvQQOs6NSDMyXjtE3hp7GPWsDm9XncL7Nv+Foui0Sk2Go3x87+6DDnYd
JkL+dLWPmhmS3bvwCLuUK3b/kmkwPTDqDI3kV2L6slxRFsAEii6r2SMJIR6Zm7Yk
XTN2E+HTevzus3R+5dCE6UMqE9OLNiBjFX6qqRJRRCFoY7AOLI0Bll0ABg0z/WDK
1Ic7JzJgfqB+wh6+ICB8qFUu7fZ/+be0N0lbWm5yOuT7WK0wYBYTWZJgA55AYAHf
6tybQPkcymRdm0X116+2Bv8C/BIMMgC1a4l/RpsVpIa0FOvoOWtOQNCRQR0vGmCs
+E1jJ0cUrsrQTYT2TIalz8PsYSAvbnt0tg1wyJ774MkJflaGjRRV5MH27BFnO7x5
UksSmhkKzJ7sBruWbSCpkmHs2HC0f3KuPRrczOxgimTg9NdasX0aW2jAoXJJ61mR
5tkVPOVyYbf1sQ/7kUBxB6VePzUdPIz+rabNwcnhTBn4Rh2kNR6as37lrDoqT7A7
IMkQmZKrIG2WFXmFJnkBfhdnOplSXYCZA5jkyvAuG28szRiq+Ur1mKT+On7dv4zs
YlibfPfNbxAkJvja/ojXgzYNnP04SmHnGObMHYXc8VEvhJeg6dq97maUxkFSTooi
/a8XYGd52gp/1J1ZseCFAn5jEcoyKrzWC14OsJ9Yjokz+QnON8vzKZNWRzxHzn/m
VidkYYxHMssjQ5l2wg5CHfG3Y5IxEWwdUTzcAVVOnINYhSCaMomKj5lioo/7rbGI
IRQlcsarc7DIM4StK6KXd34GCOQWFti59tT9xyAPkjS352gfulJAWSFaWcZKhdkS
OkmhqbBz/i4JEGTMoDxbjbO2zvQl2fvxX7FoJBfvIrokDWYrCLUUhYhKXH0zFgCH
VqGRKZ5H1QkiwnJhdN8+lg8VWrgjbYzitwu+zK3AmIa+lR2d3rjK4fcyf82k3yyj
Xer7jjcT8buTeBA1AvDQQYsXTcv2oZAp0UUNQsmbo5Wgon47a+bzVQijVCRkzLow
p+QXkdzRfWMU1WmVQQSGBV39htFYpGpcjL/GN0phque/Bn0Aua4jgi/jkPLgjSX6
mT/VEbQ8dpT57r3CcBeOy7XJqgkwVyGaBKh/ZCQcBhVdiRCZtSwfHVV+RTFkiEZP
SfF/Eexz2RDX+zWP4Zfa8nXGC9izEtYUgXA5qkUbKfylnK77d3zreJhKQg4YJUZn
WoajafPwEsowbbCKVqf1G+dUFmvS88xr75cGWziwo2RBTMvfB6LFx1Q0/9pOI7MY
/sO72wiKaXG9wsPo07AfQscSGDG4GyxVr5RJAVmehlS//JVuVWt9YULcuHOlAJn1
Daf3VhrMqjU+haUZkxdWddtzI727sJGMcd/mUs/e4x3xN/gwBSIeHUFgnFxeHJbc
NJBbrqo/eLsY6bijUgCKnUANryL8EDt4XuPMv8fTYicYBbVzqMsV2WtO3OJLCAUK
+CK3+7UxknGl/Ji6/lkpMkA9bXoAa5cCebnkfxCGE7GTGqLdWuUwUJdBSz8BsCyi
NEs7zJ1pQEPaaOwswrPxg1ApyWxviKkE6PyPMPLyai2x5uGLfUkw1XrNWLA9vsDN
Xawp5m3c/M7MiyajkfnN2J4BIwYUytOztawwdhgerMSivdMSE//aOFEUcFhowmqy
thKCoTJ7Wc+ZR9OsQhsq1n/uDAihRc/ILNQM61DSfPWGax1APsrexlXRzLbXbp1Q
f+iS6KhyhiP7umFGxR7V6XEft6RKvJAj1KGfo8b4AjE5KsRYEnqn1nOd7QkRlset
xGDk5A06EgcOVBV5Fn4TY2wYRRfrihAZE5Ija0u42/l4phoKDKV9/F3XkugnTSW9
cUasKxfyeUl80NZ/HvltLOE+4ebcT2Zbl7YV4eDwWJakC9grTIgSjj3l+sGRrBai
cQ1Fp+nvyEvS8RD9nBuEprNfehCUrhhcw1+9od7Z83Tu1GcyezarAiHD0tQaJHaK
BaBwjULPCQPo3rkrxPTjU/MjaHKuRLM/ZSuRIe0FYYG1mGL0S9ZRfUqZ7f/W39Z2
6XN6jAwezklttxH3NynJXoFxEHLDnW63pWz4BdwPpZY5AJliZ54gzx/ZiYmeoWcu
pdqdKiPKCUNj6KkqQt90MmYmQqZ68b6UoilFl84Z1p671hkZSd3ulhrqeh+teQsa
QWxyWIn7/GpWifPO6h5Vqg1wvxnqnOMon+Y7wrUgadVr9WGhFutdlcFUB5GIjA/O
ADxOEHJ2iNo+QPR6079U0qECkGX1u+Fn2LR/sD7Aq0+mEUYHLU+RehNqW2pMPQ/X
orZ3EkOahSe+eVW5ZwjzmuopWwlT5G3CF1Kqh58SWPlaKvoMAq4VsLJzXGZk+mMT
IKpIPMp7dYuDEw18I2Ve30eNTQbrqiODWuzHRf4AhXdsyAdMYo3Rb05G+POb6g5W
S5zgWsYHd7mYDTNgz7RFPCA/P0cfJON1Lb5+cOkb2KHEFHZW+An34h1vXxNEUrm+
s4pX3wnW4xPCI7Bz71/OCGnigvv9XcFZo0LtVBtThFeDOhMQWjaD5E0FOirI+RIo
vAmZa+UPQrrh3kLWV/ZHHeAxqQdxRqJBCBwynxwR6FieoFFOPLmDXwgRS6VUbPSc
QXl0ROgJzXuw/LV3uIZGNFJLhXvosDUj84u8Cwtj6bCA4v0oQwp9ZMbmILRP1l8x
K0Qlm2XHamqzz6M6y+2vsp9pUv98wqUJsfMyTDI/2qF4y3PSuk6Dc8H2qVE+OlgK
y336n/Rs8LkwBNr13m6qOHESHM28AkppdFObKsAeFMrnKQ7lNXkc9DHsl677mQSL
f3BD+/TuO1RdsIdtJnimRNNjMfNKKYdG3Ccw6SKSlq3HLIemLkP1wdcsJLikBdPt
5gnVzbu9gATR+NVIGBEwluYGTktO3zWbrGkMd5Ax5NPqlc6UGqQWj10A8740rCTz
8BPvTJaPvstLvdsuEBuRUAN4awFlQDSVuw4iEtihQqEUWZgPzw7Pq2wiwBLizTBF
wv3c6/HEsnlYx5BZdp2+PSIk/mS4Ndb5JEUMFs87J4H/brvEYMbb+QaH9KyOWlvO
9UmyY8s/kF1xkJuween04iUVG/dWgZoej53rIaPNIDIykgIRvF4/RazocJxqQOyc
y5LGNPyPaYFvV7tQKws/ITEI3/HZRtS2Cs9gH2eBGXsa3rnWgA3Ab6KYOzgxPAlZ
dcmPWsAsgYrclck0OoyiEhmnOyaQS9AquYUmKGI0e7P46VQ6ZpKN2C8K+cbmRC5j
tyNSu06jWx2/SnXQMrP/J30zBaLYeZVsmT0pASzHkoN8T923i8jKXGRNNnbI3qH9
RPu8W6l8dKpYspwZ0B1QkFq6xCWcj6YscRJCTOJb1VRGBwPwUZ3S6zICSU1uypPU
Ct1QEJPS6M3fnwWNuWadlXeJJfgd45mdJXqy4fS0+62guam6Idcv8NCsYsV0sKec
+Z1n1/dKtf0JtgmS14A3ESPetMv/fGkYEO9QWXiVA0IJiWd6JFHKfAUAEKiYf02s
XKMEJUvhiEuqWgtjH5wna95sWz15mL1TwC5YCAryeWAQVeOf5rgyIQRnxNNXSht8
gT5LYPGIT2spJO9KmAOxhnHqBfS3wwQMG5lhaGtJBQG6n1QSvRhNIsex7usUSp05
bZg8SBpQrCM3SuO0WHAln56TUx/krgI0mrYf3GUN6GeG2cWLsGZkHicRsB+nEr3/
0iLGwLXcMnBZ8dDrXH7x53Z5UC4FhtoYQdq1SHz9rnuO15PUbw1oz7+tUVstJ5og
TC6kPR6C7fm2WyD+1BBP0L488SmdZWM9MQr43uaI5H7x7Vo8QUMNKtWeWuf+enZ5
214SJFz2qRoYWOIi8+9F8S3hfxNFNiWoTxCCgfUW+gX4dbxU0PI4raxNjHD1smKP
ifC7mmdg0p1ftNnXFB4ZYwm7qetkJSIOHn2JqWAoBbSgMkt92mOCZ1p3cmhpRu+y
38o6IX25XKpPPMRezhYIYFrry9w1dKKE5wb8WQCmb+nGJo79ifHO6cPwx9gYiHbp
t55Hy3bnCSLZBtxNnvtlPhTI1gXJgeN0iLuD4+VmTf9aoAaG/tEtlRk7MaVxwhlR
akg7JEvKs0HQoyP9peICkjh3ox2R1Aaw+JTtSQLMsjtmjYxjQ0KEn8xTbUo/wjrY
+LHtMDveiJnXP77ItI37TZZ1ra9K85MjXGNmpTJsasi8T9vqjqBEcKbuz4SXxjsm
hDLah98zFb1WApoMmI+fm1KCfVhZ+0PskL9rLF9/d40p4HI5ewCYvyq29iMzj7Lr
+ehSFCkVwi3crsxIha12OZo/3f39+7h0bFahvzcAsJ9W+V6HL1OpY+T4Eku7fitg
+hUr2wqWGklSiQTkOWZdEqXoe/uD7sYJVASmX7V58afoA0efsytVkAhKOtJwxD6C
MyLVJ0UMv0x9ZkYwzIxjbO+27Lon63/saqvZL7TjVXZC8RvWqGUWacmMNOXZnO3z
Hm4kr9Eo/CQHeFv7zW96OJM3UtzuEynG2xNvAbzElYfWCzYvUDc8v8AP/70K/J1r
mVVZ8fCZmOpmGh6j9FZR/83RtUIpDeqJz+gucJEZ6iGLVQNpB/T8VfBPwOnleZ7E
WPkuBgnJYBluM6jT5HHyAbOeWnSmii616+zPBL7Oo/uoEWNZ6H7bZQCZRUtYBx0r
AenZNCKiPychV+4SKI3eMxVHj0jIGO6pxSns0oKtY5B+RyM4jNz/gZbrc2E1ranf
hzPvaQFulp6B+x7cpkvq0IOA0rQQJJofTFM8BYht3aQPYi9Q5DfkixsLoAPfoThB
E6Nlve/3I7w2XO0hXA/CeQcq71swPRrcLadC4/Z4pzUnJxceIqQGW+QLoRfgFMgV
SiRKTO/o4Y+KUj9Ekn/MPvPIrOQNlvVETXM+je+nmNQniDxZOU4CIKPMcwwmMgsf
tljHre7meVZwg6O5FypFHAExEN22mznJ0IVETwmWj/hrMAtJzZ0PHyrkX8QMSR/w
rGIL3nuqMsrK2PYEIup6b64MYK1JMBkg7OxkryjrXR1Fe3D/zHh7wDzyDrFGN3ZY
Z5BCkzqZytHYkTlCAiRkeI5cPxIGkDlsRTUSACMEbP4Qz7Bf4+IQnKV/DSzW75eq
qK5V1SPa/DjZywBbfzoA71VG79J0rDGvZMdcCFOAQ6mKQElQcXiMLODJLGltJsey
FV0KPuSltxEDYB9mkc5r3UzLXYAJC3VRwtWF4nVgIo8BONPSvWCbgsAA1ko8uxqq
7K+zLZmTLUlHc9G4UBGd+Es5i/lh+eCtam4T3xLg2fL7Omv0LmyJIMR2cDoGrHpu
zqw9KtSaRmFe+gz3XykW0MCs4+Hq62JFJDXKXOdhrI2+m/t3oO2xfZek2XomLRgH
crZOElsVbXd53i41W6CcnV+CZLPrJSpVEuOQ0wiGtLPVn7xaPFAzEB1IUUClKMhh
qUg6l5HxdSmmMLJwsSE12IIOtQYdqlAscNq7oAXc3a4zsyHEQzgA5XJwQzIv/8Zn
vS4UYBwO0m6uCYkEocSK9m7Ezo+zZdMzEZTNxyexTTcAkk+row+URQt1ZPtYkOO6
Izd6YxBCRA3fxxuT2IgeSI84+4xfiLmJsObXu5NVgYbhx04vomAq7VJIOiRN0HWX
OIr2nVmnNRLP1beqmAw32hGNZVfv/zJZBhiXho3oiUCMdHsYmWLxGa1SKhJ9ouL1
diejU4jSNWryVPx+lINd4n0kRS24FnqCA5hfHj8axG+ysrfwzyawiL+gqVB1/44Y
sccve4YrpGm9g6lN36xVlZ6YzXV9lVypXzAToCrJzrrHMMjQl+7IuAPzHaklBHb5
k/IOwe/6639Zcw4Ni2Q9/ge19F2wsjiR13kwIvteOKuWIr8acVSVVIPXdiaK8lJ5
bI8TS2BDVs+xpnGn284nVcsr8ICRWoGm7GSc6TAmOm6f/RGQLPPauHGTT4wpMrN+
xZ+yq/IXKXakyxi27iTp59gbimsUIsDrxrMemhARlcjrGH2b3HF4+DIze7CgPR7e
VQpe2JZh1tjsOACR92SkNHC6SkNeedoOmq3zDUeZGlT6n11rlBh9gm7r0hyG0SF8
cAZaiN+D4F7AmyYWPGo7Mg+FV1WJhwTyF7xU9MVVTtUIWqZf9cUPP7SzabqJX+fZ
E98SBiNMcw4BrmnoUDUW1YkGC1sOe5q614V+/+hDYYWzlk6PsHdBPCEVWo9OY2JT
UY6qg5e4nDKPvPpR90X5US5AF/B0mlamQC5vmyRmOraQXrPnhX1tHICGt3e3ofga
6O+Dd/9eIktKjm1ddMElxWtgdLRaFXFUsco2uGU3bQAq6x/q/FNw9zL8x52E1kCD
gKsrjjqrjWj7EyLVsqIuym8wTkFDBUhPJiSI2JgBz9Km9E4mjtiaW2MOoRgnzW6y
rA3vzPzZLDGXDDxciBkUGlB4tjgAu+HZy0PSUswAI5h/UZHT38oMstCV/LxIYaP+
r64ijyTZgZxINg6O7XA7ouLp768wn04SYQby5x8UuzkwiClcpaoSVxCB9RSyM9eO
UnKUE/qroQHciVWflMf/h/EKXg5RmdGRYyyq+eSeLowRQBaFfLKM4Vp0o/SPfMH4
5ke6u5DffbhJFbQRkGajCadV7GqLXHxlC4J/enQsEzkr4ZnWnnuI8F1E/vMKOob6
mVwjcVBY56ATnwle7GAZMd1LKD+nRb6Ft8T0a7AxTXP1ePQBeanrScwwq5EE1+X7
ZO2yNL6YEVyWB+uaGYRIsn4gp8dYv398YSvyFjsat6pMBcdxoaSz2cm0XwHpLBIx
E5Op05zlPkEemvRKcrCxmAEbFDgtAmPrjoIpyRsiZQJ2GBgRfcWbw/4Y25Rk3NQ1
WdhXq9Liw6JWMrOIENPdH40bKOuY89dd3IzmxixGCeHgpsvz6UyXW/0oo2E7Fpsc
yP2rjhurkIcV6h7ToBgLoT1dzC8HcgBnTuaNCBeeDiSfark16FMGH+IZUMV7ThV8
3G08qWgmtkuKb1gpg/zJgpfL4wpcEkhSfVOHGWJ7v5A8LTDowqv9/dBCT5qcYSkt
MSIUTKuHfA5OK0lH20YCPudNa3ZcgYlYB2ZDsWmcS6vIvn57WXApD8zsIxpSVHuF
YXq7LBEm9hdZ4Ts0b3zAiJF9wkenx3G+jc/ZYoyPMokvq4D0DJOxAs345JCJCar5
8IVUuaocaexFt9FOVVCVlwimPF429fz4fXMx/9dk2yvw4OgiP5aUIJ0WTZ5DpUgV
9mrO5gUeFBFsGeIjjI5MVPBkxsnu0AoeOvlyuTVQrJPccgKdJ3UIv7rJSMlVI6Ug
ZzDnt7rWflBAXxPgaT7aWOQ/X50taY2frLVxd2zp0/FwNoXF/sdubpQ5rkzK4Xm5
3TTlaiQd5e2F3kMvjDQr6VrdgZwPlIz8kspOazzkXsqItBEOj7Rk2EpyTDQnGYJq
7QWjvoE2Cg9RwsOm3Dw3giyslpawgP3QN4KmGoLmM0m0ahWikMUjBfFabTLSbu6C
5o4SMF+a7cIVowj4IlvG1OKpjfkKPG1UufXDWp0h0TuNpPXHK+HX79I9INyVGSpF
X7gdP9v+pybbdzoYSFTU0cYxbeRPS5MJyImSQTskYn+NpI0dzfm2T9X1pRirqNPm
MdIUFTLIpgj8cH9ebe6UW7JkupOk33Q930RAm3hZDFAm6s9SG6OltHCEXHQcfAfx
f5U8SOzQiKCfipaUhpmq/YM0br9eCVVK/SKdRiY5I2abTZ13cWrxov7PArasQiDc
HA7xLjljaiDUPwy8ee9p4UU1aJEXB/HERo27wsgakxMatjOsbzF/R0yU40JzfbiB
CrWT7E9xSU0w5D0MnkqQmVFl1J09fMWWiwN48TNp20Ouq27StaJEuJcKvQx4f4O/
njCShYWl+DLxxCywV+Wnb31SPxjqfNCZiuyCYrXHe+oeFnKWvVrgdcvCdH1T0uVv
Rcxs+SfX+YSD+awci+ZAyGEsTpmTt77EHQeybOF2lY1f9J4JP5R+fE8Kp8O51+u3
qGPEyZ0TN/qoKCcgUJuf4ryAlA/Co+cP2hui6dYBkv+cdmvOvsWGyO/o7dEx/LE+
s30mS1DYM/ibPNQsdpbZOFj8CbqtCWPCOU//bfYYb9i0hPpTms8Ae7/TpQT3BsUt
BcO1w7qnVHgnQdk/QQyw6AUwcMikscV204av1SdfXAEso8uvfuaTjfO9B5u2p2C+
br4H8qZR8fXX9IM3z3eDgGS+kjkfXMLPMlGZ5Y3sUv8S6jWKK1w4SfwPnd8TbHAc
DhqC/WRVVCSuY7g90/GPGrabxq5q9n6YlWYcHKIULWYUqVNzWQIxedqRzXmCxksl
e0lxrQnXqyV99AcToTeRmCrG5os80PsykmDEoEZI7DtjYsLsHJ9n1ZNfrH1TeLs1
EP218v4lJ/SqCe45qGO3NXwzYNZ/pdXAj+i1Ic5So+aI5xZYBViXIVdO0T0PaVbF
nzUZmmH5gb4H/CtNizyBPTt7+mHqsb7mzOkobGuZ9e0Ejv4PDhUwnRZTxKOOLX47
wHgiiQ9K3hHCEeJCTIbAjPdGylUH939bFMDEC2inLAzWq5f3IUrMshfOjox0wzYN
9e1PhwFuGy2uQWwLNY+PU49K3ZX2EPyUCImHDQPXKvkGG0DTkYmb1YyfeekU50hQ
C5xCzJZL9WN0pqAcBOlg0Vu0Ed7QTUu0vNB/hfi24/QOuyBgBLMOm6ytAu/PR0id
bCU7fEUr4x07bh8zEco4z5wofB0p6WURca1l7h6zrCsVwx65MampZuRKRBU+R59n
zTM+k6TvQo1rLVQUXLDOPqUPzaDl/aQ2No8wVcIxUXrw9nc21j3VQlBiGesq0YJG
fNLmR8JSFPnNHwS8RAYmNnN9H1AlKqA34CwLg9H6qPiKFdtDoWuFyPcYGA0bDp7s
/c2/sjvMpzk/3T/fHwQ2cdIPY19mRjBdfH4hVqeBO1kxhvPKHh0qVeIn7M8hs7UJ
mzHTNO651Gl24LV46sUfkZfh+EIooYlR6QX/osh7UrQlNL8VmL1Mca2QFw10RwfP
i5AykNxykJ639XnL2y0osIa859iz6OyEgAXYHv8ceuI/RefRNBvCdi1G8UkwJ6Fj
RUFKxys2Be8LqmF+wCf6qtohiXZd8HD3izlhZCyxyTpdi+uqWJ0qhVjKik6pGOr3
Bng2e+kqfJRxFf3tRlqjiaN6djRVydR3MeRImitPm0y3exw33i7dPbstHy3Zd97o
9TDJMVAKGToraC/y6vKX/+DAHyl8d1OC+UnmCrFxJ43fC9Xn/cM07D+Jq6Mx8aTF
1DVuQJmlvAT/0ksU2+83M5CUFGJoaDobn6ulutJaWRkIJZ6CSf06izeP93QIIIEi
7NVIFcykK744lvmKoyPujBl7k2A/uLbxexl9lXPFooSYfOG0QheM3QitgdRz7FjL
LaO8gnqL8gIDUIpudtJ9iPsB7e0TmZVHCRxKghhqg9WV5R6UZykhbihhxbPZY0jG
x5dQN3ZsiJxl+fvcX1P3ISnuQdLlGURvUgH3/YLmiF3grEydSM9L7iwL/wU8JT6K
WJN+5wYg5T08AS+d2ZZLmk66RP1FFrOBMYS2EXGcuI1gkuV2cMZ+WWHpes6h/57b
eIQhmqj8AOJU2hokRZDYACN2lAahsPseOaXcjKz0angFMUsudDoJp/1dvEND/Xm/
T5fdCeyij0wSb4qFh1uIxai3hkSHiZX/jMtjAGDlN/a5EBDZ1hyqqdx+IyKxCdA2
LgYqa18KM79YLHJRXpij1MGpdOSgM3HuU5GhRl6agynn8wgL9kZ3HMXVyGErgVVG
gtyo9mPLYpwtg2SwfHH428XLpdLjGkBY7weVFBcZ0E9otPEwkB+Z0rWUdX4mCsLY
nBKIHW3jUF+0CoYslHBskJxrufdbepMRCfDB9yCWmljIICvtMesMNMhlZVP6E42s
V/Mkv0VWyM9uyb1EH8UbE/5pK8OJpKHeCb38W8ElhCm8gXOjXt45yGx3o3CLvLXo
wC+QoDJbb+YEoJ9a/HeiOAOt/mOFjvdcjmB5FuZzicczenmkK2BvUiD1nc5+5Yc0
p3LYsCfGmzwvwBEh7SmMhZp5eqJUmpitmAXO3glkLPhna7K4Q+hDYu30UYEXxIGa
dSehUJ0Vxvuhcv3TbKnKJ7ibwo2ptEJu+u1mwL25GvtiEovnKmLSuGduRxCRXG5y
Sf0qAGKAuEaxSg79dWz52VBPy/yv5WVuVqBT/O/M2VC9+GdYNhSxfwX4cRZNP3zD
f6/xLieE4YTM/7ORo/+gKUdThgOTzi5LdYdefSjRhSNjI1OliOXvbBeiRdIkMwme
KCRPj3iF/+JcBFPxuN0yGrsiHEd+wD2FC8y865JQZkS04ivqocBOe+kmtzHSNBFH
K00PR3OQprpcSQ7OG68XldmqLfqj+XN7jLwonLxavKj0VGBCA62QmoJbLygHyaLF
UwZrymduI7DJnW5Cmc17Cfr/oLX9J5aGIKXnIBg7RUaaheAN9f0h48+YiS9pA2gH
2GtP9UQClt6PuMArZjwWbG9UtO/mTV3UCro7yb1c16AITKgbKVMDMRGTFeFFBk/K
T71TDLqKO1XJfARTysuEMRDYoyEFRDkIbpmuHmSw4Guw3vITPupOG1KSV8faJdI/
cIQq7dfS+Cl4aX1rTigXtBdkleY01saL6WDLkfW3CGmYKCUwYy7EDLYnCTe8uhrY
/KcMC8GjpHE67lngVus+/Aq4opnAWHnTDqY2k+QO8XkOjtxLgci9O90ll1nArL7i
j7hvQI5vTq2VqwzHziXnlF0SvPR0eBkIBm0cZ0TodInS7aMyPguPcIg56/32bPRE
DuwaIiObeEpy7+nK+LS86M1bTQm8f6AF0LgP4w1oKOrGckNYgi396r8k4+Vv767o
RHWieFp5TR2HYU/dXxLfrvZZpYxrjsQ60uB675kkaLSoUvqDmkvZHsPppiKzI0DG
KDxsUfogaY2QZ6bl+2bgoYHycJUnhhuJ7qJJyGPWvA/W5UcKjxHwQPld3DoVmuQ7
sGGdmEyz0xarDcoTR9KgchoY0WdcBRCaFt9ATR9uVziqyFkow/B76oykB7jcU85j
5lg8iOtG6r0KyvNQf0QQveM2iUF5Plj3kdbqFxQL064DqDkBzD0hufmty88+cbqO
By+0XyW23iBA3IU2+c2O5jmZLDoyQnEAuNMLY8nR74H+oiS/OYNX1dGStxiPHfUc
99+S/oAsBrmF73sJBczEvX9jcPburN9qzGZJSrUiotz6Puj9wGkF8hd4ifZ1MbpI
zJdJI69jQjDgFDtHtTv9NVa77YoAKoeYu3gP3L+L40dYi9rXBDZtEC2P1a0hQwmB
vrBf7jCDWVPDpznHtK7bAGCy/syYfPJ+TS0+kd+r/+4d8+hkpliDDbZYfQyVKloM
b6wCeBDc+OGNQSj+lhsICLun5sSAdXe7tRKFyQOvLNyQ+hUnzDMsZ8wQu2Yvjh0S
MULjpQ0Ycr5/aShfoKcwEJk17SLNEck5xe1lfCgXvRaKff3imcbFjnjNF5sPH0Ng
U07PD4ATbbv9smRjUvDtQsEg+xDKnasv2ACB3uD0p/XUZ6Q7Qfy5zsqpRxEdgxMx
YY9ev00U4j9tjzy8kqosAK+j6DFftNxOcMTu7KKraK8xm+FjuVt/xMGFtFBmj+UN
UhkrANd4YosvvHRnXIhbTzoQmGbHRiUIU64xGaRn9i1Sg7xCY7RXVFQGRi9Gm3Xx
QpUz7WciGWtZAFmYRxHB6FlsQBtM0AdvKgAZuYAU1+Tnbs/kb3uqALLn1Bq1pwT6
q7ln8K2SDVKW/mmmUty0y61XU0TihbqqWsXQUluADQHSxj9FM93ZWWGVFJ0mWGm2
kd4Xh1uQRkq0qPocxjUUFjgp8F+xkmk9x82sUKZ62VhpsFvzdpm3WFtaJIND6oIM
bpqo8KsUpZBdQ26G0yLNbghNxHCib2FnTsWs9FUlp3rPpohJRCM6OVXxIjR6NptX
1y31r0+rvPiPyf/eL2W2wceyoXOhXNmr+67bXS0kEUGc1Wy03nMXds9VNVeSM/PM
cQMuRxs5woOvlj5e/CaR3FObxTTsNAozbFco4oRbLRUrWZMm3P0PvhZ0LuCpSnD+
+PIVZuE6E7TrPozX2KUKWuYLio7uygW8ygj7Ro/NA/YftWole4PyEjEdNzaofqfr
UMbdfyfLkO9KEkuu+fGN75jj52KJcSH7oPm8vvfBGD6G9wwH/UwHpNKsV7v8fYUj
aD2P0wvqEtfyceUFXA0xCkvAxMl6pBuV3nb6lICMmbmeouftztOm4PBrhJuasIVx
pXNRXjezb+TqcunWV+Oce6WHxDWmA+jQcMSmy4Pigg3linySOtuGsjisFgDbS/IW
7yY7TIIIgAZjaLQiReD8XH8XrzxMVuwJ5WwU4jlj5XlmASCTXvhSYCo5u+shA4fQ
x7YFJvLO2HmrAltLfhf1xD2hrRnsGnVIyzyI1TZN7Y13bhqbjGEtPCR5nhFMnHsz
InHWOGe4D8mitG84dc45xmpPn4CxTD3B3+BC2mJdJ3LIyx7hWRNptw+1cntI/epG
kktTrkZv0HxVtZRLkT9DcRaAkvAkbDJQqdH47Y2ief0kOuOl5cc7YyeZWxAFKK9l
Nu43uSnydPQIwzImAQxzZPY8iP76chOybfMM8kVQ+m+tppYS37xBewXA+J8he679
G1M2PYjx2c7NkYz4hqxE5UN3+mgUeQwSisxQezIpmiOWipWzFUSmKwPg3AXZM590
31G8ilwnKW93Jn/dkT3geuEjmBmQemcs/E2OJ78phh8N+CdSu9bdQXDXuwpvlswk
JTTRwMmPTAF6g8dmqs6QfEdkvFSabBjhJrCQrcVFbQLNQ0D1ZP4KTVnYWRtoDUZh
viKOsuxBS7GkRU8k8kS0I6ajZIMwlg69KMTVK3OtUUrtzty+c2BqG/IaR3K4fspi
fSYJnKqcaapnnQiNrAxLHWBD1BLwffxPutAJI+7kVFDyhkGs2S6jjP00O4komcSK
BV8Zi8kRQjmRjqmlkU8TmW02qPd53X1XcAfUc1pDidG6+YlHu0eh+F85tLZ9ZzJF
0rIPOL1AwtWcJC9dU33jczqB0ardYSJj2+PqImJ0HB+bn/yIAXrSJg4vEvurqnun
W/jPKPvbkt1LR7aPIL+v7yBcDZlGNA0cYX1m6wfdkCZcer8qWybYVu/uzxCkrrPc
qUPya73MtN0aUp016uidjdbQ7/1CN6F64t6MwgxCPX3VqlmzEW7gYnNOzt5roFzW
vcdY8PXoYf1sRgiCJfLu4qamprzSTXpOopvEHNeJzfcF4+YAVn2E3aClPQ9Moqo3
eyW1rMWeIgD4HnDYOLssiUeJzwbbnx2gMOAm2ieAyCZrE/O/Wm4hLVHFAFMhn7dM
mjaT31AVdSBIRh7q5tKpCnn3GKCi26ZkvsxxSKC4z0IfDZg3tS26g6J0Dag2KhY0
DN12m0iSbSbEv3LzriNalj9SiHSt4NI7iurTA4woOIVRIk6mFmKfiVbBgw//AIJR
EivlvNzhLDaXyy6z63+OuL9bAj9xLJF91BO7Svms9df0wRAy66MFyrJeAzlr6LO+
sO8gPTSfbS65bDlbwmj0igbUi/RKW6zaP35Odc2xWPLVy0NrorOviQ4ds9g9SaA3
1O0lZWYxQI26x0J5DUiwgIFlyKc0Chvvj5rWyLmSYohxKQgtqqqPv8Wsq2ZCy0Y1
2wlavsiDz8dEDX8uRMPpJHYwrVR4ijKxtK09S/QRJlvc/qc7T3QTfUhtQ95j5Z1s
3kw/aKpy2t0Ucm4/P6sSZoLwtrJ2xwbh4eIfLHpXKlQxUaMI3fE1UY8L0vS7Je4X
INsAeY/EU3QeRSh57Qu8rFL3Y9LQ6+n0wBuhVzmhrUyBKPerH0jTR2+B9UWEEU+n
1fZxrm4v5arF+6adPlSjyjDEqmdvl33Q+jbKu8xCRVCZnyRFlFSmw0FNlhbrLJ58
pyo9xm1cv6KXmmbhnaxB2jrbANDWRKoywj+6f4QoLd4geGiyL7sdH4HJzsMp6TcX
aD/XHwvm7Z8WZPERkCHO4n8WiKWy+tsXBgCHlOPptIDYWridew33KLx7dPj7+X6N
lTkfHnmAZbl0xm7X9UE6UaLQtguxh9PKre9isMCFBacVBwW86VHssJ9OsMY+6EZq
/ScyUNiMW35Tqeuy1//UXn58tRXel6qApJ/a6ySkBJP4OfE0fiH3DvgoZbWl8VJU
spn9eTk0CRwWjDSJ2xD0NYn81jqt9hqiFThCYi/QeMg8A4p5Hj5VBNpPiFSSp2h/
pRWnSWp0edEe+ilxSyFiWqL/equ9KI7Htce+oPt8QqURVD2pQV5pGD17w226EGYD
nQhTzr3Pi+vtV4dn5Om7xwRWPQNPM4rhjekgAk7JLsPbhH3lBBs+Z6JdmRBo681W
Ib8uB4S31YkpLjfkfI2wF0gk7cgtRSbNXc30Nk8iD5Hb2Pz+ZWoGvrnjXsEG4fPt
QokqgKtgVQXX6P3WlPvPNCfJleSfN8eY44zrWsS21JtdOty9vT1zA3l8BXrN2NoE
2xE2otr8DEclCXZnQ0tmEvgbw3JIwILQq25lQhMDjbyWbZV9HSSYaJJa2NfGwfCm
U0S8PB0x/rHKjmWmLkNzKGz5mwZA/ebtwkSjYSxht6Aaz2eFsYZZegfCCn7d6bUp
j9yf1bTYxHPKnEft3VwcTidJteOGzIxgwPAXdlfwNh4fEVTjZQsdCYNfhs7B0IY+
nYDI8QOqZPeEGXDB0jCh5tR9uVI/lEUWQjrfZBpj6bK055EjuYgNFvcEknkdsa0W
l0VYqIXZc9zfuENlpb2z+5f1KQ5nIKVVrsp/w67SOK6+Kl3gPUMfLVSYtlS97j96
VLd/7azRvojZmNa9ONRUnyP+j52rJ6YeMh0Mjub6NE1MAubj52tJKE4QZm7XC0cV
z2W0gs8VDG4vY82W3MBbqwLUV2u1XtWmZTiHNKSAAIG2C+baLdJWgKSAfv+jzIUt
9JFLDaSp57/273tFvpAY2Mwa7VwZcgcAAMDg7JDysS2GyVmCkRXdvdRrqaq3OIJ1
NjlD4wqyskm6RTVkL02eVISdYlPx/Uuts7kpVwvKTjEKjtKvZPShoUsPqDMcu2hm
oCQ1/uSBDQcsAIo6/K3dN5vSl+lNJmo1YwslDd7SVyCNdydXRNUsre7y6nr1JswF
99dWQK5x+RQrAWd5P6Rwyir27x2hPcYUSQf3MyrElsKVDlsks6OnWRhF7BEP+9iV
HKnmyrXMWhxcTeAq0WJw0Cs4H6SUhX+j31oLHIjdWx7e9FtKbM8Gx0NRoxsePeuy
Ue8kvuT/0vdVYf1WwwX2pZVG0e7MSq98xsykDzk8dj/RQmQfo4oj1Wac5g2lHa9T
yavLfWIznFuIpt8VnMh5fzkI3IuXkp+bN+Nql1oKy7vyjeXskwBK2LH0I+3/mqmf
bER01Dmd+PvFg0xgKUuswUQfALDyYojlltHIvMGWrdFwx+AD35rwsgcJyiye/cEx
5+NnW6U4UfTApVgSzN9MXmN7IaWtUd/XUn8IrtMYKi6oEPibfcb2NUx7NZS+oKqL
x/23mOmdjt3GCfS54no9XOntP74HMrJ8uTZgnGbANP4ixfZIcLFoh5jxnhFrt98E
ziAsdqVSRetssMfSXS+aTzfRl6+13Sti9hmjMvWD/ZExKrd5q4M2kDyIwqCSgsi4
iJvOOR3ffmpqaxppHMpLtXfPgxe9DpqRnj9KU19c0osgIShMxip/MDEAu35JVeEe
ZMhuO4RZA8J6SbuTALOAF9eA26XZCurNt34m21GGGZJAZaJD7sEAcDCOb64i0y2T
iyIOBUArk6p1Zr7sT69Ff0AIjBK4+qyLfQ8yvyqNfPgORA5ktmTzcvBqXA6cp+8b
3P8h+/DGsEwc58w66dIOBnBmkeYPa1DuZlwLHQqB4MSQYFk29rjub9IOTGRwn8J+
sh4E43OGQ9mlJqPSM3u1j//er3PFv8LzW6OX787JVtWY1Ci2kw/sc//Bbk46Ob7Y
nkntM6fkdfMymMuqxiKEhrYSI9UxYi2HeSa0AmC6rJY0vV2iZ9cF+Loz2zRswGxS
iucoRIbWrBmmzrfzWGeJjaO8nlNzWsFl4gSSXOgMb7lrxoYyC+k01iAXDtzZd3MH
rORs2N1OqDTzqWyYqjU/sP7K2adaUj405C5oaRxyudIyq+LrNrg8rLtAlWpEA/cw
TJU1gyq+affPrkkZESRIH+PEvMndE5O1OvrYrMbiphodfHrWmVEswxEtWuhTX/vf
ZjKsdpBqxvR6IQeyjkc1lgjtdznqrZ5tiV/dcrs3AY50opKz3500AfE7pug9wZ3Q
q4fZfQkvi/Sr6UDJ/v64d+/ZEJMZaKDw6qGBu3RJDwZRu2RVey8fRJHp4+AshMxr
qBMQJPBHt1eJmwNOgN0cHg4H4Tnbi3Njs2avxP93vyjgVOyZ+amT4HBGIol5r739
/S7Kzr5onL/zs2zkVF5oZccN7/N7HG/xP3g1FSWRCdzBDvrkOR+LVmI8Fls9bx7z
VSrgeZh90taI99AoHJmoJkR4QF31hDQSgLymiokBPYsGwNxY845qodWDj0KhvPad
9CVACna3wWVfalKeCdu5haJ6xezfpUhUao5q5xvSP8aplEOzkN2WGW8qHBg9chz8
6gY45CQrr0jxOpLhlJrrZwUFTyunwxNmICtUGM+O6tqj+U7MSNxNd0iEmpeWd4+1
50d/0uv+6GQrsDNrx4rvVlfXnkjzZ7Gnip3EkyDoA64AsbwYGUBjKHxS8h69dbQA
QnnWcwGRCDP0ukBszZSDOiIyaA1VC9FzvrRwRd0/S2eXirTFmmxPRvL3bTSwRQ02
dWFetyjnJu8sNpeFiDs1lk2RQOa7Jt3zkMVcKf18u0ioHxJZ36epZM9vZXlwun/3
0D1wHe0nPdjDb/fXUlsJdIDZC8GF3fc6zAGgHUN2Z9yme8Tl9K5ImHwJjqs0pric
i63d4o1bz8h8IBIDS4p2shEUsMqDUEhkG7hH/d8R3hUwLTo8NlQOcAdVTHMGjixp
MVNRgd+gGheM1DpYJmU7zQaxb2fdSR15s04WQ0Ak2+y5E09XvbzGYwTT1rcL6t2J
1qIH1jIPFmCvi4iJ8KZSshJZN3Up/j3PZpRXTgIM5NBISgxwwqANLCpsnwC+5Grx
DpsYMVrR4l2UH672s4ZaQq8XtP5TIWvTDuj12cVr34+bd8n3aYbro8C3+UoRRbEQ
qp3foewZhnFhOfLTWuq+J35criScqkdVjmmQzMM8HTmV7Kjdpn0qWixtortzKB9B
0LaMxMLWJxjAHKT4RJpyL8WY3tmUB+K7zyGjewlQ/CnslzKRDEqS2YU024b8vcl0
hP3BjPcAJQSJaUOJTuWCZ4waA4NZ88qoro+Q4JdwNTLcwcghPAbq0fMmxL8hLz9p
+OvtnUPSCynN5uIZpdtkCxCBO6xXm8ai2MgFB6um5QGpPJxUpCYx0iW0nLikwX15
wlakt1mOYyet9kWgoTM8Qg1rZLOn9Vjp7IFGqGTL9i83uG588K3hk1RY3gTkiYdh
+UwmQsmthxtPvWM0p4gkhO5Tk2oHMuTqLN85osePOIduynh9w0vzbUty+dMTc6Wo
vyGNnF3CT/IqnUaEogfJSnK4Ocj86Uh/FwL2/f4GIBBn0oapBSQbHySoG2rVL0Cr
nQgrB2B/18tE/QvKtEcDGhiyOc1ZFCjJ6N6NQaSSQhcSIaBKSz1nw63s+Ej7hj5k
L8fbL1lv5s36IJJRfmaozVSXthK6VOSLBEf8rJHlmADedGjpf9vhTQLc0VQ+4FYH
IxXZNZanUQazg/g7rBfDFEHKqtRpOlERDf8dKSUisojIEWXOTrUpUWyYIMG/nG8h
MijEhEbk8TXDbIHqVypPzPEk+eRr3BsMO8lngMubGQV3dbVMcdgGgGK8VEvv2YDj
YfCZpc7SrgVUbCPLW1cDykWUHHvZivU07co3d3araUzS1hmQTi2uX4FKQh7OLvrU
a7XWRf19+UkgR+SB0N+ey3TPOw+H9vEephJxY5HobDmt3QnF2IOFBmkZXrfyPirC
RCiYMypvBTVZzusZpND6EzVNTVAQgwoExEhGcy0pu+PjTNenuIujG/uyxcvJwfeU
blVmW5N27s0Lqdq+oWhxIX5Jx5E/js7OI+zpS5lK3AyETKvy5OK5/oiHRE+bCODB
CSprkfkiyQaliWDOw3BsJm4DLPb3pTUOe11a/i9yb5iaBjtLn7IgUZwb4cPP0uay
FJJExsbcaa1X7pRTVx6qVEPptgivhOuA0dgiXNy74Px95sU4oi6Nq+mjU01BT1cg
HoQ5C45v6EToCVFpBqaZlbqY1EXw9LtX+QT8PkFl+XWrW9CZhKszUtS9zwwNUUlT
DD3A9X6l6tkOPqeOQjN1GF16f1rM8E3/f/f0JnMoMvH/2uTGfvW+q8cxxjq4BiXy
XaOjduzLs0V/imqjYtudvGmS8fyKhKXea2ChMUOzxqhyGrwLb7r+HGGOCNrqbTju
4xX2/VkJBNXckxG7Kqg5M/oJ4A9dkXgNwMDtiVi28LFmOWwPtq2kFqaVZOEvrZyw
/edGBwLYBMl2CgsTlLXhyaaWr+IbsYbXxCzL8YRu8TtMPAGFi2Ia4JaPCLTWEDZz
w6Yc5WZMkMQ+GzzLew6cg29CzCwWFZhS7W1afjPox1xU596BuH4ZLDsALPxowIjJ
nWFZzhWyOwrzHMpH2Aj51kKXfTTMAR/F18tgXNpvjHqzgmE8H+eNS6mcV9+0juX9
9AzST7KubbJCGRQstBsDOHfGU/XYpbrg1A4BpDZTB7H+/tVwQf2xNUdVEIRKf5BL
IS4MNTJlX6U95mCccWDWh8IdecfU2VocjhL6OqtUWqDKsReENbPLtTur1FwWU0A4
3hMPBKbERNgWI8PPtswTLeZk3iIp14CRtLi0UgFqRrJ4D/SiJNiTIzLgdGAimLIY
XCaGFldXe10ti0IYlgYTcuKDVJbbP4EZApUhPg6nPLBY6OfUN5xFx+cFYnik2Q7v
RAZ9hO+L7NJtbq5ZnGBl0r+N69h7D9BXXtZ5FM2vBLOE733LxEuqJl8TGSLsYLZr
ZNICtiK/yJ0ynSs5yh2j9PN3xdLG7YOTnBGHYOnzUdGW8CLh8VfzPew9A+aZ2aou
jM5irGJa8F5JIUKUNuGxy4SHSfKfvPXDIjykApMkUc6QvKm7w2BKEO9RAN7TzTOO
cj3gFzjC4uNidSF+688GM46UCEPFUp3P7fStXtwS56HlZhIf0G2czHT82xiXtEn+
XLgX12FrY1aiv+qUK9CcF/6H/1kfkMWNARlPcQbij7y9+/BGJvTa19SChHWawSbH
vBpnYkE4D3/Y5+ONE24k6mwhxkVT3NNmY9OFJsZ3ZOUHrS+GxZcA5IS61KjHcwbv
o+f+iujS6GzAxeO7OZGLgyZ82aij5b5dl5C4cKuUgml3yCN1VvJgEXNXHHgBw1nv
Pdz1RDPaFu5yR9/S8p9+7fuBF4rSPOv1Silg+M+W51IEXXIXEI0hCxVYouyM7z+t
7P797LdixsKc9WeztIvkUOBVJWLOWRZGX0t/6eibbKJ3fMLptdEU+m4+oxrCBBQz
YrK+ejIBRY36AFJOTkj4tkLQQMqhheDXAe6OkR16LDaLMJ0sVLdxTfsIzc3w9+8u
K7GNz7zgUARahYyJWbmLq0QGPbkwNeTcyFyzOYBHQYIxG1C9ohad7ip2OayXbQy2
irGZF85hUqZvqYxQHKC0bK/X3GR4aKvycDTUPSogK8GlsJpKX3lYzxcbfOs5ZG2C
qE7ewVbe3al9hVBSchPn2JKeet1gL3Pi5rkrXs2o3b6LIMXCD2NB8b9IKyrZmXG4
RhjOkoIvfwvXE4TuqcCx23gZrTesehEfKSuCjoHZ4EaW+ql9fZvBJy2ETs7Ak2xX
Hc5DsvfaDJTGkqJSpFnuaa6891LtPB+KMOArSCcKm7g7yBUUICRla72bi3OkgcA9
rUyo39RvHF0uBuuJU+LwxvcJ81KzLtgqnAf2eYRAjVzt035ZaKln+64ym+jQUDQ+
mLT8opTresSxTkeGfaohKaFyCnStcFsLJrYozepjbAnGw5iFyVjMBqr081+ua1Jm
RhGNvVBJTA11M8wHQTsTrqPo1rDWbHZYfM9d4g4mwujAdD47TzkRdRQpcwx/H0+b
kj1wHbojQ0V8PhRer18h1KbF//hNdg9KilyEa801F+3cPbSaU+NwphYWYqw3TWiK
k6ZZmqpakCgZHcMGrVpKaXg0DaVmS245P3aqw9aSfLUve5jsZaKhI6iZ/nJN+s1N
IQ3auaDwv68qO+Rm8YGZsTHj9t0vSv25C8DNo7e+rLzkyAAw53RkFww5No1PSi/6
kClDSbKjokmMx7LASkLOZrFtxYDZ04i5IklvcRgSvT6UmyQeGcgwxcHk7oZojzTL
ZrbdPF67g0bE2wZUKwXtnX7dWZbjIkbAy/QPr7XAPaHbTVKk2umkcnNi57EzeSfG
Vpwgik7ujInxUdUXWBqfo1uNaFTxklYcUQcZ0b/XCktKnalGCk32o6jcRMDuxWEB
PYRJhTpE+ZGEx90oh/k7UFBBCukLiww9PeW05xmC2ayr0ia+MJaY5ct7lqBvi7V9
3YfoOsGWd2HfS+8kX6dSOyf2XmHG2hcZ0CGQWb0HTenxTKZyEX48vpBtb8vXX+//
J1GPU1l3ZXSX8n8wFYSgUgUewpT+DODmuzJTHlYiL/rPEnvk+yeBp93LQ6Psr7kh
Rxl8b9paOaEPiPi1d9AfRVtV1REURdZlF+dRCci+U1FwefBv3FCkviLf/22tkR4D
zLFiUL23Car+rBhpOlZqsW5aFQaK2g+OK5S+cFGI+xAfOiuIBGZ5WAg9H/VgvlV7
CiDWSBQfjiU+5GBPO1hQHODzu48kExL9KXEUDSWm4jXc0zvRwYJEwg74GWuxGC0y
9tRB4S6debBBc+FM4obQRLPlYeggVUtUe0b2Qj0QaPCXRSgCDkQMXdfbj1Jewm29
297EVnTiCi+/bTZ1bIDlvd39oAB6efP6gLvkiW4NKr4zqloV6oYe7NLoSWgxguYe
m0IYATc/6jy2eNnu/fjgcd2NtgOKPXCWefRuDUAOE+zcKqWHk7wCt3e0LXc299du
TVmSxxj3OMlFzijvAyGT74g8uhrcbU2LDpj/NcDwews1DiKOh6hhQmRPjBcvvRIy
FNHjAkeXILWpydKNwUQQCSi4EY528foUFLcRXtAbxHpM/7VRCxi9PBLN6R5Focxl
1UsGmZ2R1R8textA1Oqsj89ZR+wqaZ7v1g0vqeWweuRHdp8+AhHPjSGXO4Cx39ld
ysjv4EvJBoLbnX/boqSL6kDnltDPKaFuD9FUAxCqqBHa6AF86Dt7C26qE9fgGSiL
ER39vfwp1Lh6Hh3hMCN66wR4SDbVFE3LCEwt0DGrj2p45/A5fP1C+9e88OlEEbqo
D/93PP3055Y3ws6U4VxS3lSnZAULbH2zKKW6mGLlyeRBRlNjevHvfyEHlU2K+w44
hqA/ZosfgfvbdBSjKuIMfCVJ68nNNOc+FFqga9Tt/rzqeVdvG4YBcyQc8bGqbSfr
Ruv+ZaHaq0C6kzyhlYxUMdRSt+Hd6Qmeh625VpGDxx062Q/+sLRyStVvFupVpIZ/
hhu6JEkd3wezDo74t5m3H5Qq4McMj30lQR9pu636t3w/Y9E8LNgfLi08nZ8rDp+8
zn4k35TIh/LeaD+eKkdAZ1VdNwbqRUiFC69ftxO3cA0OuRDvdr1QAT/rh/KITvRe
JvZhKNvJl7wUYdasm1/JO8XPUlopiqpNlLJ5ln8Ty/ANE3Q8oXbUo3ltudbi0H2f
gf7GUYgy6MqEp03A/xLGKgMBEZef7JopJ9LskRVtW11lIrAR9hpVwIqMVLStoxOl
ohFDy0XNbGAPm9BG80fnniWUlLZHGsa0qmF2AuiVwwgyjBBJv3nyI56IT12bUkUC
lCqmiS4wX6ERKS1mlykJB1Xjcc52rbgwMDrU5znUCp1gJj8/ql3TlGMdcQtxBYMA
sha3/Rgv0PMMejOu20w6WqXUJwPSktxtSGthCKQibzHF2CKDiMH2Z7b9TWx5Bk3Q
5+E3HJvtNoBx2JwUg08YHjnEPpdwwjowTVfANKHRXb925/5Rgt8rtoseweVNHeFi
dOT2NvnVRrzZBVI5KhAYI+LGH/UvhkWCUbht94ulZ2x66/VMzdE0Rvjt5CDeKe3l
6mcxN8zB+q8nz+/oAyxmSlkpqCemrrrO2S5S3rSpi+ZvWeVi1c3sje8YZ+et9qdT
4bpKB+t5LBrzd5+kzE+pljqtIDRz70JlNc0xao3t/zW/ubj5/IkuG2RSriKGNwCX
iriLAf+BLVpGlkJv4qDfiT3yJLhOS3vDAs5+UUsIqtJnb9dUjqTfyu/4GzrGw+/e
eV9YjXP/lQNf+sfOscYUk81pqUfwRducWAnzMFNsEvCFKSN2ha/u53icvS50McFN
rPUHclWf9EAwNeYBvr4ufrw1hFxJWLoYY8YHN+6dCpIol2RYRdHpapwtPPMVafAj
od6pUfzsrAqlL0oTERtMDVWqv0XSJnsaEONcDdz7eL9A1641XPHtQL2jgXWqSFlc
Kh6qV0NYuczvzl6nbmePUPrTabFnNisZy5Lo8utkPtn/vrPE5Qp43dRu2RJTGEIb
RRAFhq950CcHgqpTTD8RXDGIrC6IVez2oHsdRzij/Jeh2jvEZ/wWRZc4IWRzqyb7
Il9ds712fK8D/WrQVjHwcPveDV0b94NknTLN1Lu//o9usjlb4U8GCXI1Po89fVbZ
/O3g4lJufK0nWuFJm45w+OQvc64n/fZrUThuAcRh/annlqX7VYhMC1Slz23RlRy1
Z0Xi/CK2cRsmHZsQ9FKfbWvFbHPW7ROrjaT8XcwDWRrBAC+MKOnvO/iWaC2tNfQq
8DmU7y/XtI6ZTnd9aOF1IW37XrM1wkX375XTnADS0IJJ1N4uGuIROKGdTz0FaoM2
UOT08N6rE6Ncvb8adTefHYfZv7Rut36jxz94jsODzS5N+G0uDmCkM/I9OzS//Tme
X1z4COEHRElCeaqABp7bHlE4mRkbcXHH7YZd94gbBq5+lF3bgAXb36B0FZHiCF1z
Flb+OoDA/U8bbiFSMam1mm8+X/u/UI+jnTU/mTkriiGPL5rwQZSKVM2ZnLnLdz2s
uQTHqRPR0jhqb2tjEqgWBltBBQbhCEAH6Xpx4YV6msztp3WswdnHAmPOpTfgX7MU
+zcSwk1PfJy3Uh8z7JlM3Yc7nflYdZRqNxLSbaN1DY5fMsJrw9YIIolJJCch5ke9
ubo2dMJgL1mXJqlFBF9fCRQcCABdc7Ylg8cVuJkzFiZhjXZCJkgQQLJ3iZw2bK6W
UM8N2MWNPUDgGtIhW8z+7ZOocp/Kijg5MO0hVQpLZL+fkbX6wXwAuqEL7PKzs41E
g9x/21JKcssjO+pgRiqGZCKbXIhA4UqYf4mni6/C2Km3F+Nrdo2gDKFsX7MVe1d/
eq6S0ny/9bou4VZRUGUFazuvUqJva76n4ijG+cO2HBYHrzRBK48y9noArouyZdzc
cw42TzbCp5Sli2/eSlCry8r0Ld7tQmFSD5qOp9sifl59G48myxYKArGcTm+nPr+R
L4qdkTHKuneYi18ds/D96cIfymWT+NT3X/NZwfU3bXc2YGFkpzlUO4+E8yPYbW+J
BlLusyJQeJbrEjdlpHpxMuh0OjYfpe/5T2kJu9+jondZt786rwr8f8hYbWOFXmOF
9mHAgDM0N3muJ0r1tY/xf6g4MkBSkF75e9Hq9aEingMpwvjfbGlyzGJ27ux6uFEB
bQzVZZqj3OTzalh9VjrbAOy1n46lQGouFxAdinPKk+8XLhb1LlhQXCPcNqITxvsS
wajYMk5+qQ5yR/QB2yEhpO6A5pWFRh8zldaUS1OD2Ez108KmC9vvjBVOtXuF/Kvr
zM6QCnyDfg3cKu1BxMDSEg==
`pragma protect end_protected
