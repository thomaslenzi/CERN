// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:07 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gMw9sBUwk93bk17Q27q/jUbETluptuW0XVFz3JVZM1WvFxgZl3LDYel9zlisrtOf
HIDne/bExllQR9fWZVo1oJHzHEXBGweEUdK+MryBWmfBl7k/xdemJ526huNY1s4e
g1RAEfiKlqp2MQ3C8luCUxVLZPDbFBfQsC1W5+MEjwk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 196336)
Ya4zXoWmJ29NcubX0Xn7FTFK6OSzZ4XPaRfJ6qfPkocZMBtXGEnLvjkSJqdQDJ0+
NjzWoyXF1dop5xXXVIDmFBkiGDWd8IzbtTHdJFKtj4uihkEwx9FORQB5mIGKSTVd
zWFu/ZMRBVEtSiCbW7CzcRwzxdh1X+zS+XXJ1z2aq60cL1aj+NLYfUFva3DumXrO
9l8LG1AHHyg9F5Zil2iASxja1iwDUudailc7DUupvfHPYRyzdIskQnj1oHfnnXtZ
Y1wjjwNmFyc7J+9CXWizBMn5+vwETeNHNAfzxlS6XUm+iz8z4QQNZXj6UqqqHaz+
s00NbCradge5SA9xT5kAQJrcg3kCTb8KvOLoXThgm4zxK5XNQ7mcBoJaL2y4K6Hk
HqazzaaxnLi8vpv6C+vmIXIlWrXvrsXbmMh6QjsG3iYG5ercN3GgpcRZPkRmSKt0
fxbU7kEFKk4jC/4YH5Qht2JzM6t5OCkIJliTZXn4r84dDwdXaW18T6ngKr0utj3U
5Ha5M+yTUCBkUXnWORc9rpqibfgRRJjZmfzlmtjlEyTkGJD2RuPxm86BiRyvuhOd
ek7u7FwIxS9d25dwfSFUtqZrIy6jgl72mvcokKNPKWI/9Vd8uD1gcDWcWX9dGuOs
UHn+uxEUifTSmCAd6JWgswlfa1w7JDPd/Ud5Am9li1GJU96n03h9WfIGJ81s1rD/
zSsREDAxlNOCOWW0cOhhhyZFXp5roYqKg7QFZNp5up+WNbOSWyuAQx4LYCr8qdz1
acdj3CI05ptxjULxQkpx1xrSTITGJZfhF1xXA+kksUFo3tojvLlXIXG9H17W9JkG
xOtR2ZDCFQxC+BgNHCCizeSnIpQR5uh5cmJAkdo2gig36/cKURV/ReQV+CeJDW3R
HRcYJFrUDwwdYifbZRT10Az4mp5mv1ytNh6wp+2iKKPpOQnZ8lfyyCw5K/Vtpmm5
pkTglMAgt0ThXo1g28je+hJTNViN1bKEPAr7s7Ohm5pBhVNVGEm0WvEJS7hGzKkd
OPrfV5gKbxYfo8OXdrmsTv7J0S5MgTZ8B9vLuHG6tsIuUVrSv+VVgOlTG2WamsQA
M669RPd+DT2BiLwTIDhUTa/v2UFcYmQS4TrhHpAPLrY7+c8Pu5ZOWZYYc37gUo0o
7xVd5ML0wy1tnYkRAu/Xf8Sw0hZj16jyhKivn7rDfozjOcXqOSbcvTHTWqHyY6uz
yd+pFQSU/vT6d3nEAJ9wHGQcVlOkx+PfF1iLqn3e2aEEaijjAAjbiYNMWyRNr8CP
Q5RHirifmRhYW3C8dGSC0t4HiHuWaL2bytC6gQA8rMKgCzQW7Rm92fit6uxLi1sa
D5YPZDnH859bH/aVlEJLcakpGWPYKyG4cfhsCybo3Hnwpt5uNnJM9CHxFdyefpbB
Wr0+86AeA1wRMb08ySSWsAtYwCa5IzWcRiwLlNcg/A324M3mQ1hZz5DnWMw1s85/
JH3hERHCVG707oDZCRxZ1MMtxgeIWjz13TsdeNBFGvroY3oRG5F/2Did8ckzbAAL
C8uJe5X+ydvIfrHnk4nZ+cLiUVO/XL9kdmgQZnMIzkCHW2AiKsjMghM4z5VYfT+7
B7MOUUaw1k03JkvATgoGZ3fIF0QB78OgoBq1pOz0xfdp7AuMktpFNO6NpqEeH63M
Q81zRIhWoYBI2kdKZK1DXgYwwmncQd5yq8ldqCvz518BGmbWqDS2p58ZxW5CyspL
06klY2LDU24GcHJXP7WgXSHDKivAvt98EwU19/NrbLeKfygz4GslO7h69Tjo8hvq
dxZDvcHnUNRO8lUG6Nmt0hI2/zlrkArk3eABogOUEHmr9GYMWiXjhPG5MadynO0B
L3WLrK7LMfdZHfK1HRx3Rx2gDgxry27E/lY9UCjDkRW5H3mmJJkbS3mGqeT6O2jS
CNrKy17Ddeivub/JkPVFShUiqIyYMVuuP+nKeLPd4hai6UQv/PhxuUnQAw04j0Ao
VXF949FtACXqLqLRf/RFk/ok3yk8weT3kCg+SzM6b+hAcALhq4FhMtDAtwc9v9qj
Q8r196CnCmd3G4hVf1L00DWnN0Hcw+yGjHuq3Psw8NY6qTtW73P5vJSYOA2oC0+M
YtrcLYeCs3UMlPPN7dntQBtpLe146GXes/I7duI+mhTtg6uZlgSeB9U1EPdLpmDc
GqLBGr3lfEBtGK1pa+76I2j/OmxQvfA3D6PN2FmHbzxhcuIwDyVzpIZitWurQ5Lm
GY5LMqKXRCyFia94s8r0LHd8Uh1wJCxEmulqAUNAdHVlyWFpTepmMV6KZY9V5SSp
vht6A1P4zXektBRZjADScefpXbdYtgtuW7rGIo/ZidAyTDzPYnpZdZYJbqERwlI+
V1P7mCXX5Jwy6Imb1l6OMEctDfwk5usia5Ij08aWLoej/HqSHRUZEx2+RtE9Ficg
F2A863edhoAXH3MzdyHAOiAJnmGlJrDIZfcN1sz5TYL3UIrMhgIkqXHh/FoCw6xw
1SBLveUJF4+PWDq//itomJQTzd4nVjwl4YSzo2aI2Cz8HfYIrItkONl523X+rQWR
N4e7QHwvM8wnFyYmtXzgLfZExryX+n8bj/LPXvimEVvnlaiFxWRoZ1GTryfLMLLz
wepKLFhDejbD+wngGgMqeQrefubzsRqeI1dIPSqc/zceD+i+TzEt1neoXse48Cgw
4sNHyV5Esl6mDeeON/hWuLNAZNN/mhRYPUpKZGvWj7/sbdbBAgnuKkRysqm0uzM7
Xi0JN8i9Cg7Z29H7c+KjHbnU0SQYPDjmfsVhs/DneNmzPv30ujqesaUS0/VDfvej
+9RmJXkai89xichgKHF+8A3usjfOM5Hw71HuEDmgR77IgGsu2xCRxFpXu9qinUoe
T1LqY96/Yi3bdNl3AssxUZeknnT4gOmK1cZpI+MHiO+uBTbjhK8JpOc4G2HEPbaU
y1ntvH+YVI6hYIhDttjiyRVy6QJwZsSl606KatUDT0P3Ss1ENXjakTresPVic4/P
Q4JabSTP439ae4aZap4BPeCpb7EnyzXn/ehpPDcRDH45G8+EI6/Z44MxybZniHqM
yzbzu7la1HJuasL/NgbrFJaW1+FicRJjRKmrMv0NLD6n//8Ph3ACKGAxY9jVqx37
lbIv+BGaot9onJhIPpRgRF+uqV+/RykYUQslYLVCcaaYmzOosK3blcpXlc/MorFs
eIv0JJLfgybNJ0VMWRMgqhrZHHiAURFtl2+FOzuwMrFJw4X4vs1l08Mm0MsdTo7P
axirkNAbC8n0VkqFMumfQZUrW9Q3rcvpXJN5oSWnEcfoaNrzdsYM5nKK/EcMpXMP
7HTIJtddHIKdoPUwyetiB3sy9D89lWnI6RgXl5Euaqmdp5hOZOEBoI10GTP67szu
jvmj2Ox60VJrLdrua1KSa4pLcMeHdn/wVbBAhJwYTUWxSBWKHrtaQ7LYFDjz/zZ1
MKRtAct/CrNQPpS5uVYh4Qf3UP3ajtBYWeZAwYkMC8ezaqJxqU0QMOqLRE5iGIzH
7Dd/wYT+0ATEE4ow2nZeRzu6gy2VW0OON40jK0yyGaP2r+pBgzvDipbXKBAjZtUq
zFAtO6afVsG/MS/qu7sL0jYlTGeBCoHvE+qM2oWHFEi8PTJQxAcUZh2CLqypEo4F
SSPSk/jJvGyP1w+OShdMDE2d9aYPEiw5frX1/Y2oPnMHvjHgWJXDsbgoJMRl4Gf/
Wpz5agqbTLhVDR05gmtfJpHbQu7LfF1HS1ADV5GD0KoGezslhnN3YlO+8/6GOR3u
kPTfhqyntWg4mU8aRy8Mye4QbTetjEAUX2g4SJ49JYdqVtHkq6mUgTDwu7IE/a4C
RcTStoJti7keugjPjm2/6eTQi3wxh6iP9alPKBfJbdLO04ejhI7g/d6VwsZv4Md/
h6u8b0xBmy/0dVNgV71GYeVC6T0RfbZFDYe+b6WUDK0kB+0guUmMnZ+i4P9zXNqs
p/j17TEjl8JlNGd6MJCm/mg4jtB14W409Tp2p9q9+bZMcm7XINwom1QSPeR8g3CZ
Skt9Y535zdzLEnLSbScDM4jlG7KKuXpTkXxAOgmtLgc3hJRX7ytxxGMMKjiTsLDH
ijPnYbKCM3RmnN68T1HC1jAIh/UH/JywwLbC51gncj/vpk/9QPM4+JZDAEo8WP6A
IO1VT9x0qjBhPtbuYsyHWeicAJkKBLvVr2huY+U1wosp3SzjXPpSiR3fA2JZYW6y
tDrKpkpW5sT4Q4e48tAOpqCwI/zdrlGty/40/Z5LK531EKnKJ1vqbO0y2miE+QFX
D+xELRRnjJLUXNaw+tprg+zk6lNZ2rjVXVxKBJivxVzwK6Lz2ThtEaIJBgwJcSKu
GbVd+PF6S7pznaMCl8TldA12wDMLcDKzOV9wb6TvmzFImBBCkrQEWrffCRNCvJyR
pjG6yRJ73uob8Hl+qdPBmmVQyihIrjMNsw9oqF1TYZjTG6TrOx0w//MJv3vgH1yf
jFrrfNHcHh9auohfeOjQxee+DZLWugUSITyr+Gl3GSOCMDpeZhhX32dClZC5IU7E
QGeZMZcCpgR6PFr01aJQ4AW1vK+4VICr8lQu8bA+cSGbhD059flsAbY4S+vYg+hG
qgcdMhGM5CBJvPIFPDOOavJr0Afncgc24OMNdxP7kO9xo/Yxxs7KoHv5i+GV9ihY
ULSGe2nDwgD1UEWdAi0QAO0KMUGJ7Mu3H2F6sy5rOlo/3TLzbLDNRqpAbxhfgXPE
o5XBPgaFuooLOQOqyWoOdNRy0Mf7r/onUmqfq33TVNpSjV/B69jrdNU1nrxcN65a
nucY6WADuWLSaS183yOYckNdSp7+KKM8N2rleIbCOk6evorIYIJJQZLyXtlITlaD
FIRRKqkqJHDMQ/TY8v/befwAka3Kk1l0dOdiJ52vUQXQHqD5sAfONRJJqwgobFcn
jMZlzWfU/6VHh7jUMsFZaQ6dLe+5+QT2NYnUYMuTy/67XpzCXRQ9raAykx301uRd
CsqLYE/ySwu51x+utViqjqX2OQ2su367HWed/pkYpHKkhX3lknw5Eq/kX8TjLwUN
rPgxtE1L7xCatzx556sybXhKoOXnKoboVfp0dBPQhgJQIM3F5m99JufkB7WP5rAy
3G+MbJws+/gOIKDrjpRDLNBhyV+T/Z6wwiY8ComYnx7oXLl+bgYugRwKHchAO7o/
bujCkTS26sn21rfhShb4Lw/MFeP/Q03JNUCDsVSmMI3FjZVN+9M6kihL1u6G2Wu7
WP4iXa0wTGSqYV1uLbQMuZ0hKIWqTyEcWFzmwz7Fj7ur71GzYua0hXtu/DP5nbdr
MxuIUM3UsU0iKs/Qp79IotqeKHwXMBFwR3e7PRqsCwp/a007W5PYU94c/FjsA+Oh
+9Jda+Xuu4dDNbQJFvQ0WgjPZFKvV8cYpo0BPjhLNVsB+dBZ7IFk2hX85edzoaVt
szf2puEl7y+Qy8W0X9m92YseHMMPBGObL1jm7f6VRRVCQdAo/wf02Zil/lNO+7CA
8uf2Z3RebvJQrFmpX2SP/bx89oVzW6D0fYbaqyn5N+LEqglsmpXabdC4RP81Xy6q
v5TGhAzOqUKipRzL+aYXipPq012zEOM7LKF7tBcYfb6hO08I5unY+1/IOeB7BxPl
SF2LvaJm2plNH3Lx9bNjzW0ceuuWgxb70jtNjfnqp9MVPqOieo5CafNvWD3GwqDa
gaK6RpC77sF7PxE34pKiMkQ2dEjXDc2s0zDr53ozgKoGKOFQ40GLDGs99ehtOoHI
jb+RAxcshH8MgtGl+wpZ+wLzCFKzt/X8bwVZq+VedEh/kf8/aqIGXyJM8Tm44aCm
zG35/rh2kWJygZ4+8jMZ7Dk8xM9bfd64gL5TrpkIXMbFFt3JiQBj9+mRcUNryX8/
M0KILI2tkQ1AwYYzzdK7giBTiYE0elHVG9g0Uk9K2AfRxZw7FDYHTtEE4ppJMo0w
qj5IgSR69jMGnb2PpW+YRGWPTHSrLhxhzE3xaGQ2wLvjBbft25v5xjkBJlNANlHp
99W1KrbRNhLmnQJcu0JGSB1RMpFgwHLkdITMYOIX6jNL2e0CJQhDHeYcYU64UYIR
pOYoiEp4McZ9Qptb+kCvuMwFb3PIjww1aMbw4AYOuoUMq9+hTQMzTcJ01rkJ1eQH
p8llAD/JpIq8JtURe1T+MOn9/LEgQw0BVPRzvLCnVum8Uz1bOGACCCVhctuwL0At
ece19pHLFuVFzfE9ZBNgreCr9+cyw5pgmb5irR4Cg4famQHHMwH3sEkcbYvslz7T
k0GXLXB4hSxStxDGso0tzPGkqN3paLgd7oE0jkD/RZ/NBQDprxcKp5t3lAgosX0f
kCZCDrYAglRaAg7MvHiNP1DBEts9SAYabwYL69WSR3LX4LQOI7ml56mnHahIWYpH
4n1wepCy8iH+GF5WXWLKyIUfAZyH1vGmP4ZU83A54FtDft1mOs1mY6+WKUmiVY/c
GVHI/HXsQ/S2qlGzgBsBn8uORiG9c5buvjpl3KeXWzBifWeCCFALj1+ZtPHcQZni
Q88jnc8cacaxev+ISNrZ0qNXws3k8kORmrXUNtJexylwSkvR0hCR2TwL3sbVFJ++
FSEkgMfy9TLvPCaoPBqr6MPVkWiaAgrxSQ7RromffevFMiH3d8sVHlqTZQdEFT+8
JpOnuHfL1tPaolVBmnEH4TrVQI11ewvZgZWXcvJJdnJ9d+PIy7M1BMAEjpJfdOMN
zIcxvBw6hmyrm3vMiOYkkBB10ja0xcgyv7RI3l9mdrpnpLstbxicX59z/lUmFdjz
uUHmpZCht3I5quzZYfFjTsachZGinWphCE9wFiKhlJNbisQw+0lAWLwEI1io3JQf
ClTXza/vkAFAsod05SPmXLIheKaoBgPYJi7OlzCJivNWGu7Li5kq5xrx2gvhkk5/
q0vHkNHGosZ7IXL14OyN+XIZciVso7ixW1tu8ySODiahbTub4+63bTWzWJANGPuN
LSISJ7c2ySdfKYMRou4DAZEPnxkEXIgbHTeXKPjfrINJs1DJphyHjh6UkLyk+TIi
Bo+Z4LO30YDfN8OPM155h9wcrSpH8S4x7Ls7RBmwbnzlRS/ntttkKoYzF170oVPu
y+p6WDgSxlSsR3UICoVdOkcf9r+QgMbXAOdK/5ze8FKLcosFX88dOIBzg4UBGsWI
Dfhv64htE7efj17HmZR5TkgtAZ/tqmWgZuy/Fa0SNNX7buWU1QfsCAYnkaN6sWLq
WOqIkmPbL8VzhOd//89BljHpiOVj/SEVQgWRZJAFnNPXbFfrczVBcQQUx7aUybuo
DJh5zlD5I7aw5k2a7pp/RkZRdRLKamYlylkx0n0B+I43jlDR3MfQWDwYsZUxf1Je
FR73POqa96yXDjvkeIzpwqzcq4rcNI1NDHbxfBnS7jTd3PbVHgAj0oBSSmqKstiy
IKyibMVocq7j0ewIDiq0Kro0bUC6Xok3JcvshDQkhpiql9838rK3SgwBN3o+DAPi
BGzjkSiNX9gY9azpvuqwAp7H2Yws74YtK6GeZ/oCbilIPc4O6LOnf8lDnsPYZhPG
JBV4SAVwWBKvkOowWS0/g7SsI2Wcfa1yfpYSLU0/GugIms9tcBxeD1OPCBWsDWko
vekd2+OvRupLOsA6HiPGHuxN8XeqZAJ1xrXShotgxL99kIF0T6eWSqlIXBSQgoxl
XPm7irapSnQ7EX2xunXXB6502gZQ+DCik8Sw0OspM1KwDL93BjG3AkPzoJHcaKaM
fufypifKunBjOUEUdKmZ0oNiyB65qMyScHi8u67B7Jqt/yukIXrEW7lw9J+tjvEv
hKowfOK0Zf8PZZeAY6FdMnQYfIDVcHwdtqgsXJhdUUZwfVxDJj5H+L4/ka6t0HFX
PRIWgzNtfcj5OiOCzo/WNZQyiZ+kIqNw/yB5uF2aaSZmnKUz4s0t0AWQ2hMnDo7X
hfexTXMJb4Fsf5HgJ/1JngnkAwx+JU697qE1hFMIde8zreiuPNTI2icPh5wiyZfL
1FcZCbfqMKI3wvV10NoGBUtyhJc1Tx64HhEEYzNXj5e7TXzNjqDVUc8IwqQQUx1Y
Aw6AnGq9tFrcpbx5ZgDHka9LWxRM06dOjaBlnAdPb+9e6VV7m4W9FPHQnubfMUJy
qeWuzkSj8na2OK0OwnNT1MZZje41/UF1r6IgwlXywPYARLXu31v6CY0lhg+6bx6V
BjGcS+wJw7XsbYv7LaeIXwF7YbphOtEKEyP+nrgFRAZ8P2/Y76SPBdWl64ZhTufZ
GniRhiEwzSsjmKjdX221kHMoybRM4mmoM2Juc32KQ0Gq93Rykh8FEgAYlCATbhkI
bIWpuCehz6BXDo273Hk48n9Qp81t2utJKKHfYRFUflE2JAtNaXi7wB3OdLskKMZh
BvNWCRMHcXeeZLOlpVskRhdrUCUVu6CkRT3mOHRdxa9OvcNhZ8qlc6N0eLOgc3vQ
bdcU+Ue5Jx5n0QE/7eCEIr6BtgMh29nQHSQj6XFvRkDzRxHIXKa2mB05DyN42GrC
ZlESnFAr9bFVoBphRlRcYazzw+frGNxoou7RCwkNgQb5DhbwH0amea4wnVja0/33
tTTBKcHTT23XuBoIPMh4bLFUU3jyz/P3OVbytBZK++fFvnv+LgxK3p21kEsEnhSM
p1A0iIPEdPXcoEEKirM4zRf8j/d/x0wfAf+UQSD+LiqLmFiWA6uKyi5h/rGrVjc3
ExbgeM+o4Z014tO6xSXk1f3lpsgYnhGicNfBTaBgNlORg/jQnulK0ZD9IYQyFJNe
jHIskp57BaGbunm9TstTfo0yeUHDJXodWT0kriC1qPS4Th42wPHui96asTA4S3Z0
fjpsn0RmCO8FN1F44sTkZNdFAIPWgbG7TGhyWxFN2E7oy8E+yNHRB/Y9Eub7lFmD
FamBUMexkXxNv6P2VbFVmRHxlhP4ZMI+j9UG98rFLdJ1qEs2gcyybF5POwymGNnH
zwOS4u3zOZq/q+1TIix7D8nEF+mxeC/WZEMrYGtj3XBZJPbIJ3ITdJN3JsCSDuPp
Took0FMOjbyXWRGItq9invKM1NGYbs7hK1oWyIVv+IBtJBYQ1YfEbYnOmUMqxlTS
9iv014/7Ky7aza6fMYn5VyvaIv9DwNByBsYK0W7eU1PmuAfa65oVSq+Di9Qbuhmc
R6D1a2ht+euVTTc4wDeDAMvFU2cBE68MNV7lzahwBzRywTLbozKN9uF80L5CNZhY
OaaMIXvvihH0ERPankmq6iANLJH+TDJDwJoy0Usyx2Zxlgs+TnIdjP632iyB8CbS
DfX0zrViNBpK6TN9cDQXn9PvGhuizjlJrWJLWaSgLYSGvl2Wl40oz8zVCPV/ZbF1
eEiXjxAKfcj1dRIJsFK1od6MZ7+40oeAIGQVT6D9RgCdmE2lsDSmDkuUMM82hs0I
ekMQHNXXTH3sZaLe2dA4u/hjsnxGz/k/QJZLDwJzJ87vFvdd5VNquRbkAZIarolx
wAf7bcg6NpB0KXCQmiK2Nkp6XdiV7Gff6qR0PGr8UzU29qjP3jXt7zhwA2SVUyCg
O+CdDqmDn7tbuI2HWwdVM3iTQ/ky9nP1cHQn93PuazxBYhC8XkcFDuC/HEt90gI5
B/dhl4MXJp9By7a5v7IvkEEI5YCy1l+0U8ZEh5r63l5cpb0xYQ0d1Zt8sryvfZHT
8d6w6ECzkGu6qZUDfFfLcD7X2BpozjF/l9ya2HnSHX7AGz7CjRm1s5lQAEdTbPUz
rKpDegpMXx0HPUPU5pgwjce9hX77alQbjiocCP1Y3c0KSdsLnj+IIUeYOm/UIdyp
Z4WOqFNGgJbiKYXBRAwQBHy/nPjSGpIldoWiSfyHnvzv4x6Bt4kpiekzchu4X5gP
aibMaCG9dX6Uvb9ISqn5CmuhzA9Iwr83eAQwFnvNdamRITcYQ3ZJae3P5hzuqvop
EHJEepRFG8sIexvKcydLFFPIBaxCFlWVotvnF+COrFQKYFysWMyPy16O66j4mdE5
antbIvfL2oMKkzNpduqYAyndHa2+FamgsvAQcqyT7kB9zt3ueRlMxPz6iijhygWi
DW/VGa07lqsfpH3QoEYUIiuSg5ibGqOFklvfnQ+f5PWhFBmoK+1meLfU7AhCknuo
DIj8CUJFTOCdgl3ZWKaS5GnvRNzlzGeN9LgOpPYZiwN8Nlp2Qf/wm/fzOhSIyayQ
iwaF8fhia2wmkePQlIPynELUexmsx/g9yAkJaBk8a/spEV/jIxBfvrdhJ2cf847A
E9Tbw0akf5zEOeuMa06J2qRIYk7jN1TPTEwgjtbZdFmvWtM3nAj3N18yu7ngNSbv
X+vjwZxvxVlv0iiM4nx0fAMjjMmAQfbKipMbgZLJn1YwO4uFnkGNdFdYpLIbK+2l
MFUxCgM80Q4/NmrZWN3fHAwX0hIPgqso4yJk8zvTNy4GWwFDyylbdJeCG0/hQaIo
ypRFAEmCfCyuLgD5S7Eny5MFPQF16JMNwIogbcxP5SyDSO5YpXNUBvom1ReFMdgE
BSMMRH6Q2T2zujmOrcd7N8jp8vgQ62t0wLv53yhv7NxR2I9sUAMlOe/PkbWY+Ma6
drqLWO85mWJfOPYzic4WWhsjC2woUI8KfaaWIMdTEAkE6NLeAY/s9Q5ngroowCwg
eyYqXg5lgc8FocPsyFQdMoCzbkCNcfTETiCZXTnoBdmMrGuuV/LFLnoLbVVcfShM
m4C/+xMrcZU2CBEQ5hIM9GZJZX2FR53xxFe2IO3I2ER2bGBuhhc5GB1ws9dgUYPJ
nTHLQGTYFqxvuuEPpOA+HUDLCmB19Dsp62m5COUA++AJcmkhw4K0IQAxJHTCfniS
eF8ZlMgMTKD/6wPli7yNki/Z7BAgKRBA/KkAsoaUzj0dKNWSgLwpTIJ1Cc48SNZb
4C7YYO1IplpTH8T/b8YWp9xzo5LkJ06se6MmcnQ0xXpH6Y1sAA6UzASS7wuMcz0E
2495KNOI3Ro2hEdEa8M9EYQgm/fqYmBe6FY8gCOrXgVilpvzC4XLhALxm5PNBcdY
NjFly/q4NmyxE7MwdrLCyK+Kwq4yo61VtOCB8qubHCeTwf0i7Kf+v2e+jHStMneg
bJpVjBcEtQF0OpAxvuz9FY4M12WJj0vgfYPqAnTBiT1R0c2p2UFgDzgp6EtbaI1j
bJdx1lIyq3byesuDfRlZLEbaz2TXsSllW7e8BDtW/Fy4uDVgEGeRU4Ih9Nn/lNhn
ZtqWhc9MMu6D5PkXuJqGK8iTZVn+9bgVtAjIKEqOf4/RwSGQgN1LKIyElY6o0ZGy
dhvlfuZLPVaSNVRBDbb40yqRcWagXB7qBtqtrk+sSD+clweKLCKEP8VT4ojPDL0d
8ogwmyV/bOzdQcknUjUbVBW2MMtwDx3LNPN+eF0PooYVaRIHhSe2wVRgRKYGwlqm
41CyK66VAOKyR1ezlKTf1xCEKCRB3BnDxQryZaV/tIaH6LSUtVOcd7xjWjPFKHUc
XR3vtDpcYUPFTeNmdhyybBWXrYgeuYUFuUeBgX/yFUAy2cROnOtZcBJ8EvOn8Iop
jFjdiAM6Xf+4RBan6HI4i3QqJBMW6eVgskwDZ6waRBGhrqD+sHjj2IAXCVaqQZ7r
QCBzGd/0hPbapSQNniDohrH+pLxRXWoQxP18R8G5jni/ECoYsp+uSz9GaTEYIskt
KdD3ypHtEixa7gNAyjVkDDIlw00rpVp8hQe4RjB+3X+aeEu+cEMFffbxZy5vQnNQ
TrRNtPJFzjjtrpkILYUMoZa5h2PPbuIq6QTKET7oWxUv/lnlOQyJ3Lb1DXMs9igk
TurhTAL200Lykcy9PAAC24fn+rb9leoUBqZK5ZTB6IiHUWAC60oYY3lzjVE00NFC
8LrWU1KV6MYv9klk8dgzI9cmP/r/rJLB8JonrKnPg1TEY2zYrN0rKfpUk18KtXJW
FEIu4V/U480Cs3/YPBgKxy4+YHhm0qjakURGnYjyiToKPxiojNWzStw0i2Xbv8O2
5k3JYXFP/hU1SLbPVFfWgx2sHMG7YYjRHTKEiK3iE4b0q3TheST3lcKPM7p3vDv4
iCUEcsngE7/myJVc62L92c6/kKzyfhnzfYCgnqm+yhewE/9jtv5TL6+vphXQT/Hu
MM+V5hGiirYDNVAgATxc/S+OicFrUdUcp0xunAufSk7KgYF02TUHLySihcGoka9j
uH9QwV8QOY6ukryYLM9M6EqDsCsFiFf00/Wg/ofwy6oZyX1nD1Z+AVSF45x0+8VG
6k9XRU4+4mLCoBxfWhs3Gyzoz3wtwF8Q0s9qeiucxo/Pq48gRh8BEXnSxpGyCAbO
8zVKi7clHW4EdAp0sY6YivZBDYAbZziavfw9gKRUqbdXzG3TYA3smwrncS0c6XVJ
5ElkAWt8I1SEbiUjz/JmxfaA0bcQvuNHwaoQVEmgRQNNTkglRN5VDIVrnPcbBv1+
CO+X8jCxDiyrQn/WFa437NPl+HZDSjBcmtQgi9yZGjCNRRhq18M41CWgTCfLeHJk
Ql//dYo/L/5n101fUF89tNiWS3YmyfevduMaDMkFyz7yIClQ6IECqFIvZNZrQQJ7
zrvRH+o2AW+HpDj6yHylPlSGNUP9mDS4ADJDBmTlt6lHFbERV0ioZWV5VhJ0plZN
yEAVZmH6UDNk4QQzwLa7yCMkO6GiHHzr2bNp+8oud2SrFm+GgdQGBYnzeWGG9bAB
FlGd05jacrvJHoJ5J0gxvvnIlmEfNvoJKjDXT79hLVIoXXZZs57/vtScDrReXzzM
j2vwJbQfbZMfw3nz4NXbFN+oq5diPlBt7tjiciysX1DIUC8PuSODVW/cw63KuZK7
7FnPGt4FbvklwS2gil+cVQ9SFjt6O7HU6a+Cm6BwAB4Es2zdKbRRltf8LSFXTgLs
g5NGBaMThgxyYX7J9Xf7tfdvYHh5ubI6MI7+1WDuqQko5tUfqdJtDHYG3esz9ohA
2N+mzefgznhxzjn14eUj/RKyYqFVAYALFBlPHPzStZ9iyjr6X7GeR9bNNxVtXRur
vwvhj3mPnxnyHgflRdYV+3uJnsnkMGcaMWEr+r4OEHyANCl3KdGh35tEV65tk/FZ
h6mzz0f//FbSTPRfAvHebiehMXwTg4M8zd9P1oJXKAkZUgppKGD3zZ3+2xUcA6hA
IBP7WI6uKPiwMvgYFoRbIJ5haSvNBUOGM06Db6nk6p0iRZz8PZGanqumLOF93pPX
U84T8M+9vYpQeNNlzh7J1fKJXnfYHFKe3yEpR3tIia9Em2AdHhOq5SVvXl37C++4
zY8WnZnXkPUNgvZKmg1prCtAwOOTnWd96F7c4ihejLm607Xi43jjNI05+zJa2V3b
ftfT2bwDSDrfF/6LKtrBJUeKkhUELd8rGNW7JKjepXwJgtllhRCIGnqrE0xQOrRf
Xv8GWcV94hIWrxfchdZeUc8WJLBSbRjcqYKMtXFpytqfEN8ZhM/1I4vrfxrZinN6
wHARhQt3v5vUHUVzRajpLcPzFREpfKePiqYIDXckjUfTp9gKRWOGZk4Wdk/xI8US
roNUp+I71NeOrfmZZNUWmCyM5inzmvh9uG9TGVzWs5GIKZrZMc6htIo2YcPQfIul
VWLrprKjx7KShdh13OhO6ld9f9OPu66yPnD6AnHIjO0dC5sGjJDtwWeCEmWaAURQ
k6L/ZO/8g6Y6gccWuM9J5BbURRAD3MaolNMJJjSbSJcm60Yw7UDumWiw5dLMImpc
S9GB0tn5KD54cp2+kNLr/p9Xl2EKp2pWtAbwwwLHyjo8mtmedZx7RT6nuyAfWIFd
8t70DH0Nx55C7N7YUOwuSZlIIU/XTFgRxhU0i5xtbpf5uTvoZeC909Yx9IOdew2i
LYBmiviZz5vzgaeaJsybmC8cgB/MPSO8kGu8TqewH5xTLeju/n88UCUoRzEmBTch
n8R0PBHIX03xhslcv/VhdInRbqq3RDj2K/HYZjXnkTh8yutig4N6FfWZbusegXO8
JKMY5oOf6sr3/R48oSls8d6ys1vncKYH4j2vNJ35VSB9dceeCZB7LD2AfV14uLdX
tGkFV+9tKOKjVi13ZCJN56zylLjQcgnJE0CZXf+rO7/ps4o0IRjUXfZajtkcGLBp
meYbWLVDbdp0D4o2dlxopsssEUjbRSBpJ9y1AicwRTrFTIMA17dkhV4SN6GT8IfK
PfGRFFhHrk8oZrA0csYTYl424qVrX65S1V93cxXXZ1+wOAknXBsMqUsJzdn1OVJc
PIqAWHOuI0bz8u9eqMniZzaRdd88cdlWTcwKdHZ3m6KpjOcD8NMMB+eQpmyAeQ6H
/U/AM3YTz+PT+LneW/3vcWZUTCZcNQFwqRD8fnZZ/1h3pW+kMiNrxiWqxFM3Yy5u
KxIcKXz46ktuQ+8T/nrWewrD24lVMCF0Rl2QcbIaFMQ6VV1Dq4x5sbKSVwpapVMM
pOzXN7cbck15+Wl+Uny2IruiW7T//Jpk0gD9aVXptoGseWhf5GolpDg5bTOgClF+
jk41XELuNuB7M4hAnmYrFwATj2VZrQATuumPvtLbdDHsUe8HQb7jx+zotT06FPeH
TQ8dsCAo3JnlO4abaKldsIJhdVNMbwdQelquL2W6y/VeYfVBMpWVaz4ToQ8OAe89
YAlsgabpJLxy0pZKcsIeaSiya4Ti9twXbmXgl59xjuPoee4pLU1ECY/VwfhblUnO
0IXjA3ksRHIrCyQOZYLZeCk/i2bCbGY+uqAoRPKI1ZW5DhNd0y1RetaIyjgrxsK5
0ATrEoAvBqObSNc66V+gpItg1YUmGEiiYMi2le7yO+X0wfjRsuEa105OnW5CrZcP
Q+P1Xyf1YuIw17NQgFNSanlIzOBX+O2rg5qT2suICAeB/77aQ705QQOIg2aP7EIx
X+xMnKq99q0pZj9CIbcE8sdkrLUoN+pPIDKbZD6CIz1VaprZVqGi0gX/jO8MlS/v
tB6mxCK+us4hCxJiX2LSme2wZBUiUcTXSHK1qDUBQj/c49/OtFRUEavMmPucl86L
BH6cnred3YYB709sPGUV7CPBiyu9pjk1Qn8gSYdqwNEHMTrYZnWzpUzivXd/YGvX
kAlM5Vka7zil4njE7vF1qo77s9Hp/xolOV9J0w+oX6qIMax3wzURyf21uCTR25Mx
VtBfIjgFCr6LpA6aS8l7hFKL7tr9lfP9BC5XG4neEoiSAtwAqUYdN9sgl8fDXkoS
zPeFYyY5cpg4CWcyXkU4zUSYmn6QABl6jVQtSE15F18MfS20gOREII3qer2SRGpM
0cT0kDgmkXT+1KrGwcqKZp7q8Klbx34ZormULyPInqy3DIrhV6mDuZeKlIeM/Phq
mg6Itse/LEdadf76THsUK5JQK0WFtPaBmsRgxZ1v4G6ok5+wyvUaGm6s7u5NZeVc
AX2tj2qXzJOeXvF7cSYDX8qLTpuhP6UQNT4a9srbmO97OiMDH70NV9p0mtVFL6Zw
6KReYXb00h56sjA0SYL1C1uv48hIGPsU8tRJHoH0ReDFazy8MwPZZTJbVf9GhJMk
zMd3j7sQZ68slKlgmCUtO8DvyGdtO0eTqjsowqJxXSsxkpBczrfcXlMkUBS+d33f
UggV0AYdJlH07YlIw48LpIG8b84c/aaS4PiBV5F3Iv2KQjBWr+rZlZTC5HWCQOA2
mdq5Qk8I+xETb00XmViTPPeYH3oZsWFb1z3/gPfXj6TscDSLpCPxU5bBkkihLlUX
txmMtRkqS3yJ90fQOF355XqUjGuo4ykGVlI8CR75Ycvt1eVot3vdTKconShNDjFQ
Qfr4mhZZ0fajqr4m79ouzAUwcrLWVGfub3m+QqbmgwiZCXBVGMpKvCeq71bKav2Z
IcxAFzetLXN50ipXiwfrYhDhtv7P4foNhvS33J24gTsHv3sPVpigWj4Efg0ogBt4
7mTq9yDfVHPFyJenTcvA6OlLF7VCK9wmvxh3mG8ZF0m83G+BVpFeflprwTFn8qEQ
/dZv7CkTT9OlFAbyKuj6JpJC35/QkGrRdp5qbMl3JpvcexhQ12MGNur4tyrLIy00
iPR8aJiZThPFV71I5PSDILq4dPsjDEkm9UWpdgRueVFWwXf7ECBCUg6YJJZX7nZH
AR5qgd5q2TFSZVLIq0Q9R04ljXKYdoMjFvS3To9zwVlt0KZrikx/Wh2npMDsw8Dn
Mi7X5i4Ag7phveIPhTciAxO/VPWRIyOWqfHhKL8A7gwRf2btMPsmTL4T0TBl79V5
KSNEOM5uia0hsgH949c08Zo5D1m4iesjvrlPefaElEAFNbCWXNUDS4UImWJtl7qM
qksayvtqHNYvQu/euUz/iQqw6MuI4p1AKuovIiLEvcGSr9hSpgH+pMIQBHEjRYWX
UU3qbTt+o21/Ve4MqJZtmn4VPznuMMizQLDEIaHWE+SjPrnKtLphuMH30Z+JJ9xo
pqFYDmHulk6BBxD1P8uo4/KrxKph61P0TriZYo3FnkThfNM4C2SOXaSHr4iAOKkC
WeoMVpGnLfLdyCQwaktsIpw2Wyevd9ZevUQoYEDlY/kcc+GeWNSUmkVioa7wPFT4
HMT9dkviF+th9KwkysTpqWRN2KZj9pnihHqBXcbtOvCScn46fzkMLJDIeZU+CAxV
i8/jCuAJ1eEgjXRIOurKsHo8e1+x75gWfsxbIF48t/POLZuu1Z6lvwS6pVe8fHyS
79yMRPZJInl9mNjgVIDNX+C8uuGYORKCLT5ywEkI357DlZbPm6uLGBGBIC2VSAg6
SyeLomlS733DBCFFHEbUVqw162O3f7ZqGIX6nLBskq7Q8/4Z/TwjhZVX+hjfmXBW
EVTymdlRMx0fmMjONZYysiQbLluh1I+4w9wl4w5eMl24cE2NFCggBZBWwPKAdgYg
HenD1JF1ix1UkgQCdksvYsbMAcybDHM9liCrj8bazBYhrsgL1W1U+E0maYGq2kP/
MoaZbU32kOoLJ9EtRBfnkufkWWFGlB9RjsbbxdYhknBMW2ArfrL645oVyTfOr3Z8
b8EGHg81pkEK7LBEhz7dSIvQgGbiIKp3T34w72hMpgHa3/XcFjS5vLC6rrO95weT
NC4TekBp9Q9rdsE0OpQBAxeh5TMOWyEMW8UtUGGetX+l8FAwHPOhQGbBt/48VTeu
ptTo8gAp39QnMZiMrlZfzRDHUfZV+6SVIv8nLc8O8nwUE9CqG53JVxRuRZZs4TK8
lfyGpZaH3RVxKnr1xUas27qUlPznJWVPLJBIVRr3JwW+m5zvbBahr9mjqLpoypKQ
UQctViiPpu9BCyQl5m8kveOxcuB+kGgbJ2DoHVYQTaxHk87LLp6tAyg+p9tf/dAp
TzEM7qYHTEDu29ojqy/01aUAD0+5K2zsmcjvVj5gJ1/U5tNtP4+z1M/WOv7tfO8V
53JOIIpYp4y+sGDXJxIHRQODzxZ08I/bU4ze9ixvVLyyBWkeyb9WQ7JkB6eB08ti
d8rEeFZffA0S6AW+3XJoMx7MLkVDMGGW74rM8lqZ2j9LTiaK5LWY/NMX7N7sH3mj
tqFtCPkAQ1xn58LkbT1SiUN+WOpJgwEczbotKWW6aal9VQscY78ZztgPQ5PkzawZ
8ktfoEUhW9G5j9zyVPiMRv4aDWLPN8QtU1cOJjdv3UpZmREg9vM8qjd3AoH2JNDM
rwlfwN6zYgr7cPi2jeurtPJIkIKYi5SLpzH348IgdcMD1d+oujpujybpmRnWN4Yy
cOv3cAjSrq05K+37pv8vRXT7iotYefJBQ44R+S0DF7zunobYRU3TVBHv/wHRuhUW
CdUB4EjlQJZkKCQJwPbBWyppkIGd1iHJXLJD5BwGZh0G+3LLW7QYcOG6L5Qgcw+G
5f1DknsJICqRktGbvRooGalM3O95j4pfmtja8KtdH3rJyaIGJOt5dvNLj3EkDgzQ
SG86e5mFQzuqF7fZ7zwA+l31XgVrsq5+nqlCCq0oPloKvK6taHamDJwBpcgfvb2z
+6I6FkwBx/GPkNLO85Ry2MXjM7VTPp9e7yfRLvkZhRkgihQ31pUghknqnOMMTz4P
43m8TvUOhW8LapbadaHrWqdnG2gj9YfgaBhHYGY5KIqV1i6SD/5hzbo22LpfWcXG
g9vdhlZDc8yol0MAUYW7wy/Oz8GxZEk4jixD8Wxi3yTL9p8ZaXpldWle9ugi5BvG
O4uVlu07tuuKVV8WnzYHT1EXOhlO1RwBcg6Je/C6MfCA7viW29d9UPv3p2GKNE7h
Wco5GTgkHH8zHZe2hVFOSR00lwtM0X18Tw86XUOkkpyQOMCjT4BPjJzjqquVfHZi
2S5uezHncWjECRxQvrLCrs51uB1FDb+VA0kW/8zlTYvy9Z+N76WKt2c3EJnGzYtg
KPlyEbX2ONRbi6TjY5KCh/BWJp4+0qxVGhhZZx/XR1qVDJzC+uE994Byaayfufq9
JswI0hDmHKYaMheCpSO0GvkfmRWaTlMyoOmgB0RvkOXBE3oDgB6x7ecL4pACJfC5
k9kdKS7s1+SasK5MOg83OtUxlVJx5rFcDgpvbUfANwSvrq60w0L2ByjIYGyhCFqb
MOgMhpCAhlXquvjhtFxJEvmVM5PUpuY4MkOGUJ095At6rRlDqMVTN0XY8W33Ju6U
n13wyq6shdHCOi/n8j9ATTWZurns9HZgdd9kc5EOWj/Go0wgzACvPUbU61Odvtli
zYym20yr6wryZGOZnfoYPO6/HkTh6xaRoRdA+1zB+76BVHbg/RXmWi50nrCSbFlx
mWMf+sWV8jEpG09TVwvNwKEv74piN/K1Wq665DDfpYgfRNxitgrXwOWFT6F/3PNl
/JJgFNofZRrxzS66bkAGPtbI8o8W+W0qV86lnKEIlbZGYyDK/7bF53vqZnzcdY7U
cJs17IphkvyFl7ZQcRcAdeCsueB/Zetd92DAuWikFRWdTWVwBsBrdawbd/gxsbAR
Vdt5KP3ryofKwMyrfd+PUfw6hoOy4Wx8Pp+fsljLBFY4wyEF72w47hmSHRPsv307
uf8E0K2r+ywk8fF6jhoiwxFJMVwuQp3w5k3O8IR7/Zx/W5KxHmN3hiQKLRlzBByF
j2H9nXCg3zodOyext2P/sdOlb8MblXq/2n8R4As7iE0u8Ib/9R3KPd37ZhzrKmze
J0BBBPKeVFBSHpnxHSGkHDn/ksI7nKiqN2X+TD7NKcXdoVh1FkmVmjZI5Wf1NaLu
FPDaEylifMoWOjASB1wGuorhVltIVkXisVcWFC0wbuSBH6wt80iw55c4doC8mlFM
p/PPKpA2EUnOGkcWxlqKOG/nO1nG3DEkuqlZrRz9WxPWa+dxLu4brGidCyijzF35
wSThgCapyrFCUN15vFP+xrIedaQMLy1K7E2W8/vkMro5argr5PL1Mc39ZjIsS7nn
TAjUCdcJu309NJSKF/LEQY77ygL+ufTkGlMmRy4rWaS46QcH8vJ5URA1guaoLEMG
iOYDUM/KDyCQh2SXn05r4cajTLjzAibMU4/Vomy65iW7NWE58DmLJY+xsyGv3j0q
61jjEoivShO7GlMJNB15YbvA4uE7mtpxKZVNY1Z7Va7VsMf5KKP69VyNWYQokBsh
kHvYiIVYtbC6mhEPZRN3XWnC0SU7Y+9DXSjrfQhT37UfJy1iSvA2KMMgjvcivKp4
qgcFXU1PX9yswf8A9zCilnfh7TYjiRj6DyvyE/+tt+uT1i6MX//dyAUmqWoM5pfl
nDl7cgiPG2bfdtRmHwVTpXrSv+8QSWTvYNuXuKQ3mLSxaop/S9FdM+eimzEGKYd1
22F9d/TZpKh9XCe/08H8S8NOo7d4wl0aYB7mPYxG6a0l42cxSHUgEWtV3eluILGt
F6sr9VJ/4pD9SZrXBNB8/5nzsRDBKq5GO55InCI7MR58miphPgBErBYMPej6/HBB
a1w9OIdtuLSO4DX49L/N4n7o0buG0HGu4a/CxGS4v+MCRbSQot6xZdM4K7PPA+pQ
rWRaWZZg7P6uIRwPyDj67G7AEuAVoTop5/m4bag83w99sJEkiq2jmvRF+BqGST0R
yAVm/yboi0cN3eV/sur4Yv2be6sR/ESeWeg42oZVOyJofmrC3kFT7baWSmufIO4e
FM6mLG4CKagmXZLdLgRUpiUfvTKD8nI1InCcxDRkBJTnKv8UY8dTTzGDrKFeZFf+
NXaLkeLY3OQuaHJpzxv6nZNMwH7PT59IIhUsPdcyTxj+GEdneM9IXCpAu0DzApRG
rUC3R4h3YfxBgvNvTx4IeVRDacpS9WBch5vIbwhrty/VvUlwd9utDiGuKEWKM0/E
UZEgNvh/W6Q9GsA7auch6Yq8Lx0Cc9xtHQF0CpwSY8btyfBlyIM8EicT7GExfy0W
yEJf5wo5A9aNbXuSlbM/7rMV6/ZOdh9tsURziJ5C61gb0ixJijdUO00JOkdNkkXR
SyyzEXDc3JRXc0CBSEJdle+dNl9dtIeNOAKRVkFYpQcshue9d5XAC2pvvqflc8R6
62MQUdLZz5EbxJpNBfoDVb9mMcvjXNkP0qbRSv29TMlPC39bG+K3lisRVcK+5i7H
cd7C0ZN63YkxdlNDBFw2HWcmLtJKtFBLPaKQ62h3m7bjgngT4HjY3PB4bToKr0Tx
roaldeq3G6taZXKyU1lrKNi0N1H50a3cC7iA0v4ip9gUEqSNje5vBOKhSwPzLFEF
KwWj6g9sqSE/P64Z6OON/b09i+fiDyESmapb6EM4q1yMGOl5tO3z6JI4TiREtZ3A
ze+noZDII3mQUPSC77HlpGViAWeyDcFWSmkrhM9YnYEcYAK38wkI9zgbBHuGRknd
uh0XPxDn900M/DUdobWRzRMxiA0HtSyWkCkRoq4qLjC0Ibnfxb2UvFrqBMPMj+Zb
Yz094iq0jF2sWL3AZnRZQJmK8DeKeDmp4/dzDHgzlHtDnVKrcWezEMhBdnQIx/FP
ldSbJc/d8Dpd3SpAIg10AQuYa3nD8huAj8oSV1UE60TyPFOPsZli6TD9bwsHQWxV
2RkmRc+C60/OLPC69lbfvlseQGRQp0OcP0P7rA1eOeTQmtwL4qVpt2UmsE7F3W8S
7Bb8d7v/p3jEstj0KZYaw/SZ2/4i65PcmX3RuPWYQeQ2WePEe/gSiXqQu92kXhVT
6AzqCA94zinRjzo7qkH7Na6jRWUep9Ux+kwWZ4k/HH3xZ/IBJiMkSjf62jJy/r7w
/Wam8S9inqumW6Vi50blZOgnuPrS9CeBs+KaB3A0MHrpJoybFV7GlHXpc98ysRns
7C/L8PDFAsaO9+vIO1itQzyrBjr+tYgErH+haD6UZXVlr+HJZu2Hlzk50YYDbQ0z
5zZhWzltTiChZMi2quyuj0Cl1hx3Gir7RcT7YH10VAxPohgn3KboZ5mFwom7ZSYY
51QEw6EiNfaWkKfBhhw9sQT6ODUfLbN0WOcGvMzCxvCB6lxDK2gGNeWIwUramuKE
A23nxi/6aZodlW2nPFyJMNFbPaLZ03/F1bxkJQdSOUZcel+lekiRkZe25DekYbx3
g10XnLfHjyu2KILzaWG4ZHhavnY414ejAHrKk5DzRRMVxvNKgju/OFquGcmH8U9J
sNzasledZcs7vrU0YNf1ecs/8OIYymtFVSq3gr6VhhJdmfeqraIyfF31bDB1mMuY
93NWQo5xtYZt/OLoGKm7R01Dzmo4C4Q5KyY6ezeXP4tifTlxRg6h4LPDe03pkAYe
WXzHOB0c3PCHLPnaWfgJFquz0BkrlEPqy/YZnSjhPwBm9XkTGdy4w5mlyB38tVL1
8DkAwbM5PevHVHQuhnWfN38CtNLW1nUPNWJO6HGUjSAABgOlyMrbRySJgJI+4JBt
QsWUbBu6oF7nvwccC1T0FPHsQybgy95y+T5pfhAuRkUEFVQPYOsdwbg2XGCljpe/
q0JoNjsyxSdinpfLg33E6KXh4nTsPRTyve2pJfv/2bAYBaMtD57NxIKpYm/eiExK
YVZWpvi/J+h3zUO0Oj1+xDq19or3oEHfkQKAWfs9JVcxPmosrcm6R05j40wKljcu
Hgzbd0Zo5Ar6marmtpp6s/nXhrTUGWk4P7jEkkxA7r8SjXhlhaofuf0nbOGLmAgC
djH/L3esm8u67c+tGBBGPzopAstXJ13GBMKGBVNUpmkmfhchZbARx4QIdRg5mAHx
H2pL++eLiOtmDjineQmOag/iQ+H0HyK/fbAHn/ZPoQt4TmDWcUaxvvO2wy9Y3+73
DnSeLroC5R6gXxEKPSW6/UlZfb8F5J4ZvRUzZm/1+5WhGL+IcCTiT7PqtvI23k4n
FdMdX9lNvy6W9KdBKVYD57ZWQGnL0WvSfx9LNoRALyIH4vAntf78ImPLy2JFtCLv
v/R7x8rnHiIKI/iOcGuLCVHCXLxp5VfVtKOdVsIUAXLKOzj0i6/jvJQSAiU+u+fY
dPS/a7uojCLwVKHdfYE3RM6u5fIrwm8NHf0Cs3sGYpJP0xq2gw7FSmx0pJIFDDHP
qg5M/FrtIJHqTdbiNeunjXkepKOjGYglIFTOVJVGsev3Lfn2UYNn/CGQPXpJdq3f
fE+Vl4Cc/6tLfhfASgcQu/habsc6y7bRl5rNm0p2w30+cChNuUNUR/2hxQidHnhN
ND0d+iqhYTJmSHlCASlELVxkFMg+V6OMmEm0EaM2yq2Kvn/HOBb0Pnv7Gty/UXM+
RgnYzqAeUZqngzY83jPZn90yvRdJh1JDDy5gqnKuyNr3F2digbCmXLxFDaYnJMxo
rE3XC0k9xVQvB55tIx3p4vW7IXRVrCouc+gGoEGteyOFEpnWB9RcTnCg8CS04lFG
H+mqKoaZGy+hauQ48kPAcwipkiVpZBSLNuLq90g4ZRzZFk3FigIJjQRltv/TaUol
8s6dWgFWOW4tPM3x9nVEyB5TWePzQp9MlDgyEGKzRtWLUMiWa4Q+ZpPAsKt7MnuP
S+0sXEcIHoLjADBLlfEb1LCB7GpQo50IMdVlcODg5IsxhsYT8CdQBGmTGLipRQty
vN+jAIIJUhcWvzegNNbsQlhV+MGxCRr/SJh+22wa08XpESreQMGbx+zu+5WK11Bz
8MqI5/fwZWJDsjQnUAxBzsTszz2K8yPNxZK6vHe23gVSLB+KANyphWPRPoN+m0yA
rW8dGdpLpPy1Zx5zJj5KcekpK9F5zYJBSwE+X2SPoxi+oi7S4zkxpUqV4DuZyPFM
N/wc505lWmEvP10TNDfoC29kqQBRlTcGDSw6Wg5eQ4r8LU5VDu3Eb9UDwznykOyY
i3hie2NHmhXW1XOYzeGcjDhQQoVZsJJZilgDpsBIJg8129B2yiUY+Nh8ZakZ4CSC
CFYQTd3BvSbtW518lk0hI9oSieB4nM0Qxvq1AzlG2L1kB0DU37+I6mzH5CeYDUsI
+k/+/PlddBMRdgHCg/r00WCaOJMDn+lNfStn+Wq1FBY9iLoaTxgsj29vwsYL3a0S
REigVtsrfCwMlfDD/Q8NCgo6CJdSPNoo81LFvPP0CGvRV/LNyTdNBpaMXBaONFG2
eZVS+ohBKTSpzQqRd7QBkgNoILak/3veaBR4E2jaJYZKvEGP+Xpe9vLB6h5CBImC
FMpD4Ta22aksky3DbLFlffnWwBiKDYn49mP/OEU6qc49teo/q9F/u9++LTnrPyYl
8yhVDI3SNG3per8ltvSkfnnmbyT8fuMI77mV375iGOKTifugifV8vgz2dN0HG/L1
d1XAFwyGkAWFJ/PSG1ld8Z4QcW0FX2+2Rc/AiZbjfaQqUh68w6rWi6Xxx1QdPkkl
9ssXMc+yjw2IQzooLD3Ytyz/xpxOmzBvNmANkiXTHedZzmg0JYhXhCKIsGiUdjvL
j48a0+mpEoHihQ/206zVLwzqqy7cBkGQne2OhGPziDd6pvjMcYrACbcoScBH+RTO
vXGB82VDyJ0YFgwsix+u7yn936TCkHBEE0eA/V2UZsnKJD8MFDte/L/QAxxSuB6c
fBMQ+BWiFFrF+3fNj0HVuCUpt5eNEe/RrsRp8MGa4cBgps7/YHq/rbwxeUJH9kZ/
ZaepqmvleJE1ACStJSK4ZtsCh5GK2Qq668gjap3REIg63ehijVocW/n/0JWwlVr5
eyt3WKavPw6Kofwts4qkGFhiMv8Bqqs83vPBpA4ewPKSfwQkoAXl3ox25nF5VPwK
SGQ7BvKL5Bg5L+fO1rIRhXZGip9jOhftG1FJZ/VdIAILrdMyPkPiOpuYhb0rlJ2s
TLFh02FEyun8nmwWCAPC44AA+ns+/BISl1R4JAtZ2toAB+W7itaPbIvZmmjAN7Yh
8SyTraWHJdfuc57tHZv8y1YO0WRbztvZiiKVV66zKJUuyI+FLcHDc3eXzXNEQ9cl
oMcZY6N8cfDQEQ8kC09EQywIPtztsg+4pmhmBQixL731IQ+/YxPTBIr/Jhg10HCp
ko4IlNyeAEMYZoUf7snch/rT5haD1V4upIKVE1c/QEzVqh3+fhNIlTzZlBsG2pVK
QCnZOZOSGORgFWrj1xaWX/tBBSY7LJzW5FMgxTSmBelRjyDFuZO8mUtSq9wG5Eoc
tcHsj/SuhU+D6KLPcIuywUsWNK2OdcYjjPJ/fxpGjkKJiXcCnDdauUqb4YmkS9JQ
Nps4URcaEme7hnTtzZwiN4neMxdLnP463wc5xzCnu5sW5G6hubWYgB2X6++ahwpL
vi5beDjyaxXcXZa5LoaEBu7ITcFq2AV8TkNaZxOr7rGtHL/HLetLhANtvCBxEpfN
10vE2j1GhWHrd3y2y1Ijvgko+CuXn/04SOkE+WzG/o7ewxcsGWIIINWoG3kqANUV
wDBXzzoJuBme9QQHOPPOA2pvQYimeXklysUUNhwHMUKRqRbCcDTlbS06sYPQ6kBb
o+vev3NK5VreUqNL+dMIzfwlE853ubJGKW1TiYOt+gA9u1jvqSRe/3X0vt5w+T7v
A54ZXXbMaJe6EuG/3av15HbuXDaCiSs725JX8QX1VJLIP9MjY99svZ8BJ02nmV5n
N4cPfOZlHx8WLH4rUo4S24SdnOxv2TXfpao4R1jcUpPaz8ZTen6O8PJsEVGU+uVn
2YLXqdVBsKWmYoCroqvvnXU/DuSqJeJzCNjSDPdS4LVq5+9rexC4pC2JaYS1S4tz
CznLPbxbL5B9SsrGAbkPcChA1cw45YlRMTdtINoR0NyqcQuUBzMKZqe40bK4pZYG
y6XnKKjNwwVSbyanZaQZLbm1bnnErLJ2UZhsAvyMA2jTgPi59H9jDfhRTRSMub6c
Pi6LMf1HZ2eJPpVy5POsrxJvG+Xp4pgjttwA+GiTZXadgdPvu1rIZ4feCDAwWt0V
9a50G+yK2tda1rUX3W3D1WAmNup2MoU7718N16EX0B6Y8flEgmRWqMMB6zQAicXP
yBP4R7A3ri/axxPHoKaumK6LhFXYvg7tbg0rWnTU2Y8wcrzPxgca5c8RYkwQ/nbF
xgzlcp45TL5mpCcIdE6+22TME6QTaVVtYPU350W1K5bC+SprB59hK2xh1tULzDVG
vOlD115wxbVHAiZgUi4w5Azo7xqRve+nNTDwOIxXhQdZqAPGw+HHdI/tiVHBaBpt
pXcE2NszlfP9/+3jGXaYJ36ERMp9ibNktfhVBDuKA+v9mmSXOUL5KJwt3ttXDQqu
tbGfehhpemzBCVfS+tKM4QX+MAKdIqsDAl5ro4hBSexYFlbSJat1dwCfHxZsQWTL
IFhHXKd7oHTgkVgP4/A18xu+X8QgGGzC5A1nCajtLOwtR0nqD4Fn4bgOfx1sQmxS
xF2TmF/xEGHXvvO+oh8wMdBNNf1/ecXZKlYxyiuKDXR1/VC0Dwa3mUW/z/G9yzA3
RSUw+43uMLZgacgcqr2i84GM66RwyYWdVN29d/S4XQDraHJb98a6e+1rEjO0cJx4
qdqyydrr4171SJW1ol/1QPGosl1bYb8ID9WfcgH+0W5gJKvFtetVNZdWGSr1janx
DC3Larso32O7tvh10xWu86a0ru27HspLr5sj2Ph+wRiZgLElD8IRmIx7tDUOnQaj
N7VVVrP6ohLXWl8zEU+GrJ7RcvYxsRDGgusq9NTZx9ZF3JTeb2aNWetJrwtVTOFb
JNu5ChNMZIIp0PeOBy+t6mC3WA6qDmfQSJZkCiHRJTGCn+XFjyQKUqrXEIPSIQHX
f/BCq65Sb+hdm8TTVZoenEobSay7lWtKo42O4XwKT8NhLR6tpPJdt3BxXUvrWrYt
taARrtDs8cgkFtpgdgvbBDzaaCebKBbifUMXFW/lZ7wLv6T8R+zja5g0GEvqIqjg
URpP3z+mG3XUhLpm/e7gx5xK+2FDJwVNIpgEDZZbY4REgV+Ewr9yI1YwDXMQd/ef
rJV2vPqJoOqalmiwclUFCBY7NBD1vFXtXhWRiXSMyCV1dBnWHtuD/TDs4+5uAnFY
IBXAbwnaWQNvwCCuJQ153JiDT8R/CWUSLMeiUTSQZAG7cxpQDZxLPELRMuIFTlEU
nJ5eDQ9VkHaEjakDIkIrCkUPvMyhnudd/GwDrBTjSP0Vm97UqSVWluF4GI04yDeP
syQIXI/Azr7PGKASbRU04nTxIXDM9wyKSdaKHxe+7jabq4RwHTpyHDQQWwjykq7M
jnPa66sC5SWk51jt68tvdjKtclW0HyLz9yToOkm32CLjWPTVAgTZJM5McoJrkGT7
Swc3rophpdKW007E6kU82sTQUzRslZCob3eXySDOl2MqrQCRk/i5bXjPrMqRodY7
M7Iki5WYM7EGSlrRHjjwGxKIvbKkwbQCVJKumx+YOteHyZa2XGuT9BRnc7PyrYUd
vw2qtFhrMbvnTBcjPAPgUrUcApkgSI8R0YWrPXcIyrEyajv9loUrJfJMF6xRMsAg
OioiB/twMHQ3EdjRvd4SAWNLS0HFxN1uWHyhJs85Ctlh3KqpWfmK8xoM7aHmsoSw
4VjuLlPaIrOsYXnJuqdL2jHn1M4uswoBHez220pyHpPAmSz0+gorHZ4cPjIaPiA7
mqMyFGvqV33YVAIohRSepGZMVWp3nlUD9rZ1qywCxyv6NqVgVWlUKt+Zd3LURVnd
/aP/WbSahz/Ydefxl2bMx/UJ54MYY3gdhBWEOzL8AIe+L84iBybnuceTdrUiksNu
/lL1RVih5hhzyew5Mjk4dcoKyeQp0ckFrnDwidz4aB7ZByyclQNg/xBsJA5+HG91
Ab98AJ/CB6h0eOzS56D+NrpXvMQ8ZVF5G7L1RTSev6Yu7mG8JO9nWKPDto40sp7l
IPSzAmMjktWrtHe442hlqArlGTRt+E00I6/Cqg2fd41D6nlHV2jdP2bJILwYeg9l
I3VRRhY3UPpYyY6n9jdhPqNRcEoZtjgfs+dr2ZYdLrvoEi9inb9EdG+FFiffbguc
2QTn5iRPyTXuqrDSIT/PLP86+1qs1uPeSmUtRDCj6+37nHMz9Tw2UNoSe9myCkEv
jZlGpcS5NNs14b1+xRy7z9lz7J9iVXsCOl60Z7nELaDmizzvG/rcUYJuDSgWXjl+
yI832vyiauH1/zyUHeelg4m9sV0O0CxESDKllCLzecIJ+8MK5rsstaLkxx1YArFZ
Szcwf+GqEiT5AClL4hECQHbNAZnqBXTRvkxPQ6vE4n0gq3mghbZvaaD17RGIywNP
DqLCByP1aJqMArPo28og2+vrCu+rGW8PZ13Jz95SZ8JV0t+27E72MxNZ+dXpXkCX
3h/KMFFTBS2i1UG4c20rt7NNBA1C9OoMEarSmIVi4qwG1CAxFu9jzk44DV0FNdet
xAeVjBPxnvqkqkYpaEnb8Uuzx6mXQKZcFFfDQi192UtWAyaxYeNmsa6WbpdFF8t7
qiSJPK5LKwSPkUcMxt+O5Hq/u/aZzprhdbV3zkuGFHwFU5AjA8LXwU7hwL27dRva
hr8FvT+GPIJl50ION9daFevmCxCOv0V892Qdic1npdfV++jWbPm7Au0dcbCiUvK/
9mmLSQnRT+IaOmuAKqwhP3LJ37HIi8aUHf8hRKPoQccNYUe4q3O05H4OtkSsddCk
bAaXpFQwoyOe8KCE2Z6GudqIL+Cz5mZ19/luUa9t869tWziCx84VWdcRvHV+bZec
3hEvte79r71YvXTjknQq/jGiSqiPPls5s3YXl7lOTNf/jXhl5OiO8bBsDyYbc9b6
OFCjEmc0ylhKwS4c2HiqKKIPWWT60WEoEo8C6rFdNIQfrgz9T6gPEH8hmc0K7P92
07XXXql5jmKI3VC6GND/X59FcLXyA3wzYxz2mePWcH+kGQ1Nc9ZMDacK4HBptg2E
kCDkByfc23Bm7yzwCk8NiGZY0sJoAmI329h2RHuSvtLnptoP0tlLrVi7kztsL1CU
n9f4cvfMgAe9T0emohI2p1TzQfu1yL41fW+YpGpBal2pVZBxnih7eUcinijF+qoD
HPCmrxLS97/CpjE8oy1nfQQyWGBHM60jjWuAKOA2KySb3OQ857p245wvis3KtyMy
7gXqD40GWX9hMUe605k/Ewr/FoCSn3yo2uVeC6wEVcMly2IqfHLnJ/5lHLOKd7JO
HYFwDgBuxlY+LTMe/H8MgJgcZDqoWvtgmLwkGRiVV1/qsg2DNU5OT7ako6Q6rg8x
V701aP8b/C4dLy4zi+bYwGO5cNKuYz//Fblq7gsnwcCXSbpxiEvZ0AMtcUDHhSGS
2KpMP382ywvTn+N60LeJmAwuUyWi4RhQboRp92sK7jwKwe9xxUwXP/l7lSJHM/6J
M9/VUUjaUFrQNlRHauprCtXa1GM51iHGmeIDsK9kkzIrYb7EdLdnpQnHspfuN8F3
MgHM4drkWbYNXdgym3QFbdF8eSnsAHTD8lo/jknl1wkDnBzZeDYkxud/LCBCfYXx
6G8SazsufFxezQkNtP9PSnmVqBH/0X8SiVBo7A7vpQ+PfHvxNFQ4XKI1DqucKP9g
w06QkBCdkh1gty3Jvn+oGQP3j5AXB6COdSJcnSs5tzobYtMhXgbjaW+uKIMK7n2y
CmX2ojmmB2JzRlfu8CY/bb022iM64JkTPRfTHHVzjabD6OAAE0Ahv9FTCxa8e4ch
XMI8EMSdIUusncs3y2Qh01PsIf1Uk2aPMEYaKvdxfXodi+xl0436OK2p7RhrXsV/
qTQz1uRieQ0ZOJ4qN6k1GW0cdp8N5uHxN2/TgzJOiKGFEP6h5fND+DKOu2iRjrKg
bSml1ANp5QdqcAsBjeD/09gfsE91zf4pHWP17JWJbsooeIt2xcxCGqThpgPGrx0P
wdKomkPDYbAwFUbRmK+yHddncSk9wv4hbGlkJAAPuo/J6vQS5eYd8Ri1KvXNzzRn
VQUv7xO0Av1DRVr1I2U30eKx6kZ+11rJCFPgG6eR/sgQUXHzDo2vYHSuuciyOEDG
a+v7/DQOQsazX2zVxQvZLgVVj8+3U0B35OztS5SsGz3mjKkiMHRBlvWI4svzWg7f
TK2Cce26BDnhvaQ4wBLtU21QMikH/uW5i0x9WP21CACzyBufaETppuKM67uzIst+
0ewBKhjdikpNXJ6jSqe0Z2ElwOMt81neD4IW++nIQLK2zHVld4oZzFxLTTbwfwPk
6ILLblzANOt5DUq8xrCsm5q1jyY5MbQWpH/eUTfWJuychO07IIfrw+VqcKBLxSuK
aNCE4SGawoStAR382P3yulG9cxZ5hFwNySpSEnJdBKPuzzJfRtlxVZzHRhOk/UCA
rK3SSFZBiElvUHdqcpdXoTflXTAzpGP4QDJ/9nzzOL1toM7RgiCVezF5NIkZ8GVt
GZCjgDBltk1iUc9+Kb13JWhY5T7nIkfGvqykGcVpBn/QISsnZgX5AUvwTHVwmXlo
glLfq4RNNjzaNYhBRjFcBYXf+qccp/wqA0H5lsTKBr/XGtu8lVtfmIf09/kCwjy/
gVGI7TdIqf0UHl7HbyDXjc5/pI0uEILxmovT+NwUngSb9ciLKLYCL2GAHFFN+ikU
tbTClz5ellwz1E0dD5amBbM7v4fAo9rlDi0wALJVRi1tUO0zB6N0mn8n3QvfwHJY
xEDd3TeH5K6AwWHk/+NphXWYbiRep1VeqdumDSjFm5e0aZbyBm/pzWH/TTuqFDkP
lKNDjv7V14bcH7dBwES0pCjLETYR0fPkxaP7Sk1MvsyRtHXSQvmkSSoJhmccGQtb
ipd6hPpO02iAlzrWPBOV7lektRCJ4Xhd1ZSsdxks8POvSBX3D0zaBhDByV2SXiE2
3xdQXx0HkU/uDAT/PqC7v4XRSSqLxR7p/fossBqzUua2qvTY2xSN4NHm0oGh8H95
QBJ6eFk2y3zpQz+iCQqRbmiLBhoWyjZBkapDDWKiUieCxvvvLM75Ylg5+i7M52Qb
jDWs0hUhqqXjmVkk7Eg/YHKCT/jTyFeWNLXYHyiroBO+FNpiejg/2+2b+Zw9gHSe
w0U/WUIA3goYTM3OXdg3BkPeZHbW57Rdn5PpTnsQmH9d6Wz3Y8wVycx2aDisvB5l
jgvi8y7o/BCPlRzIX3Dau/fmpksJBJ07SyjJ61okEJ/IqQ+E/H1Z39ZsEOyPaGvX
LOtz/oK8D430nMzKpR/LUaG4+viXkGRhPenvVVax5K8LQYWmbV7lpub4TQapgyYq
BDFyVtlGVemhvTvXNMEWoKnrvzdd7+gT1MuGBfyQg9waKBOssKKzRces51XnvaMg
Kgco2CInU3hpg6BWT8PBL6Nji5+TvB9Su/s6r1uBM2G/BY7+NyFKICL6ai8vpY5V
Yg3QS0mRIiZu9ICVo2NEaU+Dl7TR9Upj2zgm984sWO0ThPiKCXs1J3bBSLMYggN+
vwwRHXxzc5UQ04MG7tibBGC/fgCB1MWVe6D/Td+3VcYRKKWBUk5aQNjJhyLDsF30
w3K66kwdUs6kgqO6SDZi3P+UF/Qsw674QDHUkD9Nz7UvEcsx3p1wuzFNqfFzpnMA
wTjPJGawAum56YVNcZl60+ZCnMcY9W7Y9pnOGm6A4zMp/d8dgUlhJBmpWG8YYqcu
41xAOe38VD2rv9w2qLpBV6IE3MJAN3dyzDW+k4DQi+us+arKdJibMuFgWV9Qrjr1
suVQL8niUIR2uYDYGqsYC/E0YEgHx3i63LXzIQRZTu7N4t10SE0o7MniDbIZscrc
kN7wdzYYO2yGOd6qyJto/xmKaDnuFFv8hrsoXMWpfd71wuaQli5n92r08ofj+qVh
NQ74eUPos+sEl4UaZFSa4xolXQeESQONd9S8/UoQdyVH7t6us0MUSaisbK1VnB4a
ieKXG07RP1wA0EborNRuX27FkPzaDNP2xJwc4Z78jrN0fkgHsBRxCpkjH8dvKb5z
bG+LCv2RZgMvUZ3arGKhIuhlIvGUJnjoSgb7If4bKKYMfs7R2nls0D9VGKSBQKjg
N0Xbnl9BfV1hULtYgFc3Yrtw4FUKTbkVdTmSwzqQFIrTjGQ3wQ1v4QTIbE+Bp9a2
5NMTdFv/dtvivqELvjl5sqtK+45Ot50YGHzz2xRGBT4XTI+WHAGtS55P/o5EEzWP
7x5T/u0ry1EBlkt6d7oKh3dWPtvA2ZGnvHeSpiFAw+gL+/MYv14jV1L/20cJKjdC
0xaWAcqmWizHTxF3PWQ6in23Qbp7c0sK8Mpgf4M+CqLqOHVftgOqIuI0hggIdXao
YCmgTa5Dj28aEKf4ul8P5eS4qGyz6/rnCoIesSPLL+RtqDhE1kbl1P1okEPRgmlD
g0LGuqPhUY8oLOCRi0lGFWJ5KitLfhfQ5A9kE3EwmdZcMflRm+jZel5lnRelKqy3
eAcy/Hq5KQ8AuFrdWudTu+ca5x7udJ2lLSXTlPKsRcmkrpkw7cK16M6PDE5IjnGd
ea3z0/r8ayShc6vDu4cZVMsuKnL0Udw/OqQqHAeWlJ7kznVqNOjhXDPHUuXN8OKq
5qD3c0kdNwBcHGfT899Fd+v3xk3RTt3JiTHq3OSLyMQWGps0wR5Mo7ZXQSz+AoFc
bChcFptxPPyau+ODsUPNtYGGCOBuG1PY+xe9AlhEuYPvbRxuEjb1gqOh4/C04wCD
w6VoieFDESXmycNG9Q/DhQUP1xjjQunGOKjDCv4r7ivTSQnkNH1nksFj/nEnymoJ
K5OhhTos55390kIkHVy+KA8M8cA2aei/+X3BA4MR1IyQwhP7C4y5KupgLMgg0ViP
yz4VPiu28DBsEDoEzZbG3ELI1dwtlC5m1jzcbacVj27lTymfduaOY3LhtxlTwvmV
Uz4DDvyBCJD7IOmiuD8Hjd5Jo40GguX9buhqC3peMEtGr8h/SgNyANxDdSmCKgHQ
9sBrMUCvwmVRLDEJMHKRJSwOnhp4P1U1F28/h/QE2jxD+mR5OTKFbpnRuuBjzYNA
7VIR7j0Vi+Tv7Vm/a0U3QzaTKFGMmdotmyNeSX0jwQeueZsvfa17U/Im0YPPREcp
d1JP7VwFD7+pQvdWsX5kAP92pBWmOLizJvs9xrNaVt1Ik2DxKoJO8MPr6KEv58jw
3Lcqk/9gaNMjMvsrik4xkJ3njXH14SGdnkY6EI7ncDsq/cU9c6vmL28l7nSlJj0h
R+J9iKSUh7/T0RmrWvK8NYzp1xrURfpeHFAHdDOqS14jmAFhWmb2Msu4gdRQJOMZ
dBSBPNqDk4mXYrHbo0GgJppUrdsfcw3C3a8GiPiWiBicnNJSf84/u3pKefxTGb4q
8+VSvXD4Oo9CYlKhChu+LXIJjMKEkB01ya5bagE9Ut0BHp524uc2ezNGK/LRWSic
pp9ZkaoDsN/Ld0TOv0iJygrBFdjN1Hk9zihCmruAaer0mhHCnd5y5PwYbiUSIUhQ
GT8xUxdFa82YGk0j9E1xK9w6GnhQKDI2YatsyF2pIXpQmkbYmtG0v8KzhUALGlyx
waWiM5QRwRdlAcmuQsnMeQ/GYqPMCzjnf9FUJ7d5f6/1fs2qeuxTzOoj+X3hHgIA
M0DgPW3FVA7WwD8pZJ5aLmEOriRcHRN1RJSi2jZ6E7QtIOnDB1gNmTn1n7r5gj4v
mqMQR9cMDVNuFqHnA5aF5J8ZZvKFIy8gqqPFW+5gZLJMgdn7wtkxYnq2qa9bdsnB
XIbXPsYOTfmuqKoONhOdJSqDLoAoQrl7jqv+tR+BiR43x85rmBaaA4NdS9Jt/MTe
aQy/yCCTlpHXDGgaeIqkIX73DsOsu7r6EA4uv5KO8HNL/XgszuNY8hOPnfaB4PEw
sgNKiQjlHgwZwho1Fo7Z/TYTeaWzrxfGc01vEoEUFilQCEbeMsQtYpq57OfNh4AO
H63wXbD4vXoq663R88KNbF01O8kRTFj+wT5AEXwQAyIFB8chCZkqyj37QBzGlAF3
rrE9q3wXTQP/ZsZe7AJdKjBt2/y1aHcHBCcLs97FED0/X5dMuhe44AVMttb309V4
mQDgHbD16XGtWthBaLqwwOzR/9iGQVp107hLS2aNPi9RL1BO6LvOWJzsa0AikWWP
oYYDzwwoak5bLuTCOrqDk6QSZlAg2iJOvLuNdgVEop+aNlvFa8/yGo6vQLGEc3Vl
nI2uAnTNNZJD/fenGir7z+JdEy93ru+Pvr2PerzdD5l++rnbVrN0wzfe1LzbgRBM
hqB8c9PZH4EW+QIYD2ViZZMfs5sbZaYcfafoUV6WLuhKf+t427EavEw3bnioiw1Q
xhFEl6iOE49fJ2m/g5TCl7Nqe738tzCZJSAC45qdvjk5OaskISZGaV4Nzz/gSDwD
7+eeLtwxaf5J0uYJtBr0pzeBbToh1kEvD+EHR5G5Hs+d7t4wsA2Y27/2vVN5PYJ9
uDbkPGtdrQZcO6Z01uhYp0unT9/mNyMzt4/7q8vW4qnZPkYUtFWBYl/nPhAi1GQV
uOBAT9z7YEBS8QP4Nji1RE2Z3V79Wm7jnvn+9fBVRGs32Jyoj8LPqTCmx5OUeJ8v
5AQbBamUVqQMy1aCEAZkYWRcfvhytbKp8mPFhs26rpYpKOBR4mCo0YELVDbDE+Cj
GVMxdMm34TKVPvLKIAiifPmF+58+kdjUGQpXZ5GVOjuielMF5VflfakPAC47RJAJ
9eZXrqceDQ5/Sxfk4GxPomW5PUgfknUJigU2lC6SMCxv6Wh9s4OGNvb9TRM6lMbv
JlZqh6esuo7JzEPSzF1IJ//MwIMaCSkhhqnDb/FUqH7/OWhHJzyaJzaPMenlLC95
zW3WC2OPPSnWM4hPqU+T6Uir2ZYBj/HVssBrJNdEA9wMNOerokuuj/HkYiJgRZg8
2Ff0KZm9b4t6Z22VE6qJmHAN0aSm8ca5lsaqqlgdkzaNWrYcBkaXgivF7+/1WK8a
ascRc8pQIK7uDVtvaV+wMMpinorgiFoCMraqLhma0KjoPSGJu3LmzK9IlKeNC0Ah
dyzlbCbraWVbPXEqcheJHf3M9/Q5Skhabs+9ZpPz9j5v90gLP2W1RK3coWrHJOtO
UwNbIhXtbmYHIWZvkdr2pF/ifwQYB7sieffHelmroIRFVPkkSG6W8kJCpREaMkCn
iV+ehzKBOQeq8jtd5sg6LXKbVKlhQXJYALKMMk0IfHZ5XMeCnSI16IVJFgEJIYHP
dXqA5p+jlf4j5XIOYFpCixxF58SuzgYR/ujtCnv9OyDL6IG41IWr1NF14T/VDPcc
7VzUdj0y91OTwEbEJo4EzBaFkxED3WubjxRGIiHbi7IYz/7oOPi5E/4/l3EVDoU6
tmwBrSESzdYOagYNOZhFIOY1u1V+HtmuapVO2Zu2Q9mzgo9KwMEirYjBTnrTQIhk
XS0bHhMSHokHj/hrukKs/v9EVBg2Fwbwf8yvOjp6wUT5DbZlEiKCoo8UKdgcB5VN
8yeVI0XGj7R14DT2sKDaM09l7hl1tPxVR2yzaka8S0YX/qhLq5rMykRl481jDdOP
5ylKgBsnN5BxZAqkimXxUF5iP+wKpR6TxcHy2QsoL99+oMWff8feuWhJvyBmcP8o
aiM3Yb6hkWVqgGe0NB2DjYlkK8cAEdxb2yrIBWU43aUVGTo9Ytw7hoSCXihfzLE2
GN3ksJbC4X3DylMqpqz0D2kF5CPaNatQU72W4NXqhA4fDh9TiE1J+/Lx3rRMPaCT
iSdKmhyaEBTR6jSRiG0mCLpbjb5X6bdB0JAYwJpIr7Lbn90w7uXzswoMOTYkHh7N
sx154KtBOGIJW5lEgy5SL/uNBKiI+NmqBitsxbSe97UI2yidy52537/jJCruLTcd
An90OGq3VHsCWh4M5hVvVYeorbQ3SIXrx70tA0A5CKZIOxT1moXMxe5+suIaesfB
LCq/njnJMpeZtUYX+iOZD6Uk1faolOg+c1Pb4H2tiG/PKwQe+lC+e4kptvYd2Drs
QZ367rb8u4J3ueAe4TbgwWYCAVQW2ngbMiN4+gAN3R8/ksGtz9UZaxXCTil9Gpxz
CvKGLO7yYQOwTaTAg6i8Ycj1vI38Ps+xJSQiNQgtxFmBlWhMi3AckNyPLZQOjvfe
QmD676HEIC6cxMOZm2tnF1W4WntUyUGGSF+t/bNBBF0v6/E0lXth4/KQc2Gbxm8q
LoamyS2FO5Mmhbyv0MegpOdose4o0+QqipQdhufiq4YMLINnp2Jzv3Iih7yywnnv
K82ZwhGgqYMYYwt2PARncIcOsrtjH+IawgKyo87/tLZ4xslxMNMgOJ7lLcd09CR7
Bhb//09Hwx/K7kLB2bmmyftgp2HsYdCMfHpMSkGc4wExcnX9DDKXie3mVeuQKahE
garUM9u5iIympyGy3Eq2vSzXzr9YrPOKza2o05S1iubOSCoOjM2jEDuKj96jALE7
tqXKoOjRrf7NPxUSiTjH8Ke89QNVC0o+PevRp8Q5LUb7mvra5MXw2Fo27M4lA5Fa
4QIyI7fN/Mb1VV4KOMkh074220YZus4acIRKN8pRqRTcTm6X7jh6HMiNQAsnmiRr
7P+0aCsLslJJX4feb7aVgNUahassnr8yhX37Ll39J4J2LBNwsyJk1DApwy4IdbZH
VdxPd5MO638poQVKisvdK1LFeo82hBy85boMbnrrTcnypA+3PKrNg/AzubtSpPQI
AORprOI4TQdCWsb4TBlhyiFHs7yhv0nVWS0z9qG6+6lL/sVWzYyLHvo9gqa+6H+H
p1i3BEqvibAeiYI8y86FTp2u8eUze2C4bkKt4yOSv1FnM3fUIOz5+B9PaG3jw0FZ
LnJlnDnK/dnLBgtj30jHCMlcK9CFSMC1Z8O7nNfjv8jlygaKTB6LCyRRNqOcRgV2
knQjZk8n4k64GbMZ/l1CIbDd6erQPaIPTRvpZ6ttM/LK3cR27f21nRrrGayKdRjV
9ZXbsmrFwSMJvsIOHt8XDdQOqsXPXjw1iPkum+Qqc0WZH/5pWFMxPIIHWZugy/Cr
PvGfMaBE/5q4o3I4f+6Ew8kkgAoiLkOxTd8bH9B7tgzVt/w+FeVRU6u9aEVFogm9
qScwj48O7qGheLLskoIXfas03Ht0PSJlQFkZwmqfWWXdET7vGJM8ebPapI54oKHZ
r3ry65bnPEKdjz61BynClxIzDijOE+W6CHo30HwzyDBBI4aQJ4rGsvA6QeQK96u3
ioygr/P5dVIVhwPoV7rOvhIe/chHfBxdYodGOGl5Xvj0dXaVl7AMejhubk3lc63B
qLndzHNG8c1YViKNGCV67v8/847iny2MchXhruwThq+XiMwiDn34I08aMJm6qPKm
yzU5leo2MaG4znCIm0vPO7SVVyIE17rbG9LLGEdVpvUZLYbIYQ+4nBPrhsPCJcmI
kdGr6gS/LT2v0GY3S48oeUlSkyIx5p8DGfCSXP+9bgI6o+NnG6ytcQNcdZJJxJpW
bKA5U6GK7aAwW7Ou6zcsW58va+L16iNyYsf3E4OWUP0daU+oc5918RZ1fUqziWrI
kJ3NK4dzjmV5rDSj0kAk/lmlF2YUZeBvkPhEaegaWgKSLyadmivLNslekv+U9y24
iH00udo/tI4sWLwR9MJjRJj2UFfePxlahQXkazxg8Xk9E7eVFQCyIWMcP7a8cACy
UnGeEjAdmFDAQV69YWl94Xkh8119hXh7bB3KhzGbx01gfLHwn5/+foLFt1Km8qci
qJoFRycX2gUHjxD7saEHBtU4RhNTga642abUbqgD9qgfi9PlqITrZU8tVhbzX0j9
78GSb+w3lrNbq7/t1TU1yilPNHV/hXzzVf0CIPpqo0San+74f6L/Khl2omlLtOmL
MhJZT7xMGhqlRJdwEKY77S/uE2FseT4l8REwbq5ACyu2yodn5e8JD3QbnR04dNqb
nT1GWsvodTE8RFwMusOFZwCMJOT53CdAzol6dWLfSNQqWDKsCQUR6Rz1mENLEDwO
uHBWDZAl9wclqRAHor1lTGilcx5nWfRi3bJQLueJTVQb9sDnj6e8bNBZ3cdG2lK+
OpbCoKd33pNmCzmOcrZm5Nk9aF2Vr39j+hecpkqP2nSzYLvGi0hgfOXIkZeJT8z8
Ks13NDRS7+yDfaLzr5EEzIF4nN05BbagJCaQbx4/yCkIrW5fKhAOgylLEJ6lgVdr
DJlB8LS2FrUl+9i0ISwNYDnBT87rIHtWDDvUQicwobS2xsYH6DA2eLzeZ4M4LdhZ
n2T3yQYLcx3cI7I1jlhDa57kjB8qlITh8kEqjVoHeZmIQgPlxajHaGzlIQQOC5Ee
wQKaJDc9HKr3C4ktqMufVAzKY7hGjuE2kiNJDnuTUqSSUrfvt9AqgIkIZDbpBQWH
7jO3++REJIZId/CgOFkhGeqZ0RIA6aIs38G8GfXZSOifeY9197iFcjH2wsFD0vez
kEaQ0/Cv6JZNvo6vLcDbCjUiSuWFeFoxv0yWnRmewfg241XvILOzLgRfdo/F8exa
TF9CoKWfqSD2TfruH6YamIXVS3r+I2kgx2ciOQ1rM9zcyP9ZjPYIZenj5rfdSilw
zk/nngR7KzeGL2DcLD5FgRgynNUsGi2xTBDgywP9Z5hi3mnYO+WysNzyjFU3omni
XrKRMZ6O5IeLbNyiUqbE/Kuud/fGQ/kSFt7v626YuEf0Uv7mqImgDzxjiat7QK2v
7RPG6jiEZE3yRKmlkuLf5Uvg6gfmckhBgYb+fmlpqvRu9EsipYExoGlHEIeZyHKB
1Q/9+uU8uwDvFzEea4eYumdN9uewULN8Gwaq+7eiy1r2W58aLlXtD1bLhRpvotZF
oDFeG99JRqvSLDEcTv1yI6YImkOfoehaytskow8sAHsw6qVERB7L1sV04A2qZrYa
0C9u6rQ0xGHYlUowehUVcE7xluaBTTwxQ43RhV8ulLSRrwnRLQMisPP73y4kDMOp
9ISpZtV2wRKraVqJJkxoRLyd2U97R/s3R8urGqzy+UhWpq0quCyNbsmicRb4JnjT
9eJVrp3xyKUEMWSY9rfuc9t+BPkgs0v1C+6BtXZjdKPuMmdtAMF4ueF6aaRRoosb
mRgwNO1zxFK6dX84wk628+4jro70ls7buHaHVEmx/Sc44/2j5QIH94BnWSUBSiXg
WM0aFpDkWRXob/fHQlDdsS/UcwDJ1VU1UjnmvOfdL9nACYSt4pugLS8aei5KhVi/
qLsY5lO0RKoEeysnCqL+PbW56dk08gNJsYc5zHv/NDUS1Od2st3oqzZ0lbftcTA2
JGign8D0PLJZeowboTBTG77ji4F3IgtiNE2GOf73D+1fa6SlZcHT/xX7Pyf05c7l
pB9XSVxbPBzGCw29h98cFsi11IJqrFYjp0K5QPc4g53VIcYMH/P31XY02KZi4glC
jYg/SmsniY6oOwDJJeKqkIFFV749MtALcgmZHqptiGT7fyQdt8EVJIQuh8v0XHKG
to853znAxu2mDe75kFxvaQG35HjndWqq5xDAbYEpeAbcWJAEWBcwj3EsEIj3mv08
dLv98Xy0Wf+5FtyYhw37fT2hBgNZzjMUn3f8hIcgizLBLYrRLeB5RSofPHncYVWl
qXHqIRoVLSi0dhK8DU+LYjCM64ADMwVUCOWWLPYZbtaOPwMP1xcCtAIxDbtzpIr8
fGbwOoowRPzPH6MNc2SPM8f1l7sumo64mL/F2/fA5n7FDSlZCWjA/JEV01wur9qq
9+9a/M6NtFTVbX2548kUewKK9XEgeILyVEfS1pBoXtPiV8MALSKDtZiQpPnj0sDA
GR1HdYAwCFLxJDkaEwL2PYQlh/ZcXWJzNeUN1upopq+n1h+RW81JkBj7xRZjBNWt
05sxvmdKFAuEHJ1D7j38sEGDWlpqiTT6s6RYJfLJ7CuEiiZJ7ROI6OoW0zK2aCmT
acp/seHo9Nuv+D4POswLBkKxKMOFv77M/2sWP7c0fS7aOj6WwIsghKGRUZM25DBI
BWoPum5dTWtj1x/KYEQiPEyGDu84XgVM1Rsc6OaincgsNqxFMciUnc6iLKqEdK46
QPZwvkDwgjrK7ym5igKWfTqV1tuLy66FIvv3RgszxN46ZEUnQH1U+LfEudffJxqk
GdxNhmp8aMUn0akSYu+pJaG+FYd2MyMYDjdSitYMivLOFH/40VoZPc5eDY3MQa4u
ehk/M/Zl9FV/otTK2rIp1CSl4icuMOn3g7ucmrlT1PZr65Jck4bnO8IIjtz5LTVx
pCVdcj1aI9lDiKGmc9uw9UnOOoIVw1Yfb5qJND6rkrsIWd/HbDMHjbdwavp1PANT
+phCDl7bP8Ty9crMMA8ZG/th3GZohbuzZaLPjkScKMrJLPbSDwLaXz2a9+meAVB4
brgeToN3ZlLEbF94qPu40r7y9JIGBmRPoqDvv6dylPrdKHbXKo6r8V8C+0n/MVY5
s9umlojhSLG2Oh5x5w1JDvXaL9IiNDcdCtdumpvChT0zyi4r8tNahzyyuBkpxh0Q
Lv+3p2aFLTr4wIk/QjXx+Aj0uUwuw0QVSi/V07q0AnRew60sJElQcRT9qcaK8NAQ
BpS7wLLywjc3Icfpl2wi8xBdxFwwhdZDbl/92Zn1ff1bPyw0rCchnOwNybKWrq+7
k26k0WTtV9wOycBLtsQk8k13F4rx3USZ4HULe9lA2t7hiMW7rp2rPiCWcIueLnez
o98vSYw4OGcA+FQxf6uE1rQ59yLe0PKT60E0k/e42JsjjPJ+xgJ+ya8rCq/orqfY
/j9RRj/SQhdbuKKwd0IXSvQ+uqwWnop95Osh4uZ+Rwv53XwZOateRc1gxq8ms6yY
Xb0dngkZrCc6mZYBh1uo3SWf0Cme630xTj+cZpTRVGUW5cv5h4wi4mrAb83MdFAu
GVZMIC1WxVDa2EfT2Qg4E0c+2k8xM6BmTvuvIZNPCwzf/q6YkNnukfHgNAk7aaCw
PdJw0i4C0zsA51lZ08nttzdH3UPCIrysV+TuoGA9pH31YMYeFeEyOd6glty2yxB6
3WrjD2REqXzg8BUebMfCIEHJjZJ8UXg6LfNJN61VuX4oswbO4a218cwJxXZwhop5
SRtS1yq5BUaaUivwJlZKnvtCHog+vFpvbHODcMLY9ta+Anmu+1Igd+0l75NzJ141
IRIkDcAz1nn9Bqda6hBJP+U4bm5k8n9mFo2yX5TM0iSIZqu5SsAfrgbU8Hg/5d70
PrJhlyOD+PQIcqGguoRSZRtTScY7Z2GE/auCeEwuUzyS+TToLa0cru6xgauOo99l
v+cLyDx9ftf1RbBdMTuTDRZtaka/QbIEA/Zdilp8BAKe7bCrilfjpXKnt8uAlpRC
fuJxiqbtiYJa7z2vw9ToK1n7gV7prZzclkDxe8uQSa6Nr4q3EC/xyFE3WkgV7fZE
psXDQ8yVy5JSxK2wgG3kiXxicrWoeBqQPT5lL3kjj9GTfw98XLHAijvZoi0ZkdmZ
mUYrju63PqmcOv1PhlQXsXce32i/QNnn1IFHq/tRphwprS2G13you9u8DWoMh/QB
Umh4ZHe4NJ7STecokW0wWnU/N27hmgd40Ut5ucZSb1qsWWcLMCx5F/jjFwvUQ0sI
+a4BxGCqsJg+P+AzrZYV8vz2eK+e5xqWgnoTs3LQI98zQx/ON3Oxx8N1cHO587pv
0OkVJByKbuNFjb23pLhCkZWTzCSusIDzshoB1NaX06xpUDRl2K+fltFC6dqcRbi1
/NVfp5hRJt1k6JE/Mr+l6IXpzG/y9T8lbyU+mx4u99VSwwmdL6gQYb1xbxyQfIUe
Z6bTuLKQKp4ypaECDLZxLAv7WirIBheoaigByRR2CCn4LZ2GTNZSOZonXufdpp9N
LrOCJdU0vBsMNAbHEoSavQORlTSCBvSVeM8Bb9ynQubreRSNG5i1+GwtIXUTPis4
1dDN/j7oGIaKA8mgsqumYusGuasiMxLAGrr5HCway0I/3wluS+L/7QqqAvxdI26a
/uqouozR1o/C9PCjXV5ebrU3qwDvlRCzJKVLthMX/pLamcBUClzv7iT13xLnbb6v
ai+3f7QXy4mcVgooCh2fwV9rnMRLRfBOfahyM7CRPqizvBzrYufbo7E7FEPrxmef
sEtZOKqKXZ95nLrgVQKx7Cr+zO+VGqT6xGNiYo1KFNDEu7XwivOS/sX6nEHRDRCq
ue7nu5ZSocB7c2tash5R0EMFDoDjcJ2U0SnxneaP3X7qyEMAQKf7GKkZw7/Z8MiF
t+DNO1p6fk1mY/Qm7r05Xm2usy5uktWpH+dUzhaigLkslnGrYWkX0I273zQw6DMd
UoUa18AXAIl8ZkBZOOJxsI2Z7Nxg/uGk43YYzKqdmrXMcRJdYM5aBWS20IaiuYea
hll+E/E3WHVg3zFJG0QPZk48feYkM+5lMaKUcqbUhGOA8IE6ghf710yweSqlExZ9
gndfM3RyYA5ZKE8+9PFYv5AgZFMLyAYglDpG+PxwdlbWKUi6Y14Q+KYlq6OXm8qC
oGXHHGRiOyIJI6ZkFvAyIglMw+HFl/l0GaLg1e+oPG7bokY7ImbGTbPG3/h9I7aC
PSEci+KE3RJozSTPEim1WLfXXzwuitt4JVNvfhWL/0+jtHJZQvdGCEtgRAMR33dd
KaNcgc41HVgH9H1mtvoMIEpq34DITE2XpLDmfJ5p0ypgYafLFAa0GXYoxRbTaq/l
wJq/L6iAkaryaAxIe77g9hB01xNdt1C6+XFBVVvhBvfK99CZWrDoCILDV4pLv8ze
/Yk3vfIV61RD56RqYmzokWKbZzM2BRRXUcN9XRvy6s9KJ2BJqgxLm/yP2Co11LKS
l59uWvFFyYA+aUpKpjjY9MObg/ngaC4dnwdocrv/q5iE2nh066mepA2VFSY6v4t2
7Mos1r/ps+6DyQYmnveHQA8GkLADmoaINK+hQmNgfJF5q9xhtAZ7XWLumIMbEDqe
yUgmn4PWUMGS70QrW15RwoowT9ecj6bTadwO/K2yYxEpEHUck00R7kMp2t4JVBTA
cvPAf5zNWy4Dwct8huTnbjexAwDzUHZu89xjG5RoRCke3LeO7hJC05fGQwtQmNJN
ZMy3G9MG+jMSsuq8/P6TAR+twArBWvIMNPsQXZrYkdfarmg2FklDHB8GZUZ9nYYO
HMGEZkuPJYP9BTJ8jSmY8D4DZj2Ts+o33w8YnpnTg1btz64aRh9QqcTaE1Pm73Cc
tj+37l2TNlzQFEKB2u5cJQ4hjJduX9sfqnX3ICuQDEItMSh7f6pFE7A7a3tv5+gp
err4tC0ScCCQh0/bs4TxzCNMGR5Nnt5PM75QzG+BAiTWOBv5V8fP7kz5gvx3s6hA
Z938X/Y154SYWN37f3BCHhlQRJjhnpEXi2JNyXRN6e+Zy9qYzIpsPyXhItCEVowy
C060WxREdIUxaSLS3209+pM34n18sFgttZKUM7AW/N6jYsuLHOPMYZ03fi74xuqb
LYaM4OA8ifSOqzsF6ChOPwb9loyvr9JaEZog5wEcExizuk4KOSKsMVhqwXmcUhKR
HVrKUGld/QC+dWZFpiv9pMBHnGnRIvD1sXJXVfH7wWwuICisfKCKSTLjc9UvkSzV
dg5LPgmmEYTOGxEx79e5J7QAvAZNAg1CT4kABOVQUuXLHSYQKiSI0f4XjeFluj80
U4a16/XFGCkFtd6r97pLYH5ZDmE0mBUW+LM/gsezgLL/RLYL0quTRSdUUOIjLM8L
Tcg+sG/pBAs+xMuVtNkGueQIfHYKat6x58ytvw+sGTTN+UWeVTrgXxRwHdPu0bwr
aGdebq4k/Mg+B1zS34LNTz/k+HREEvHf6uqwQXHCDQDVsJXC3K+q/yoynJv/kqGd
ZTRmJEmORcG4R+sveM4pV76Dc6+BxirMCOH7nwCu8foz6Dhq/vMCcHIxEDvu0SZk
joythgbgLNzQZFQGwKeg+eakX6epvvlfXwo0a8kidwCiqYQkIjfLb4MdZp82dYD8
he3Q8BRavrrxh2GQd9V7YxRL1MiHBOjKwGgXn4G7H1820v/ahw6fKLd1P9ft3rEy
k+4ITvCpyGstBUT8HQaihWWGg2Y6ueaAPKuuxWyU3IsYvCMNiUAnaHJkiXPsXeY5
TMMHcxe5BBb1XkEdD66UUgRs4CFnXH1DTzv2gaJUjQchIKQm4h4hf4Mo9rX8nr8R
Y8kAurvGS1BrGzFMdfzZqSwM3XwD3I+wRP/Omfog36cBhzBx0Ok5oYPRLJFaEhbt
eFDPp50FGu+N/vkRhCR4zmJwycRUNDk12QWd0Wykv5vNk+ENCmoCkfzUSzcgr8y/
Fm8NgPYhNg+S1YXAkMN7VsLoc4fOo070QG/wp9ggoCSg2GsRKx9N3gSrXYoRl4vx
8vO73Fxl5NsLJshktjYqy1WakmKZ0EPtpuGcOlL9epNmcKcteFyDZluzZz3SRRYx
azP5DpSRtIAdT1o4UQz3EIwTVXZJXV1Ye/ojurFF4UvNQWZhuE5n5qub8CPo93+r
Ps65A0rr/Ll+ozjjSh99zU5Gl6GWHepI162maZ9NUr49sSctty+6pt1CRpVEA9uI
mffyX1CPijZ7A+IGEAmaKX4PV0y7K5Lxv8CjvIcbt81Hl4Z/SOgALvz01a5zgsVk
Lo7pE+N0ZEbuUgmwX51sZulK7pztF4I1N/P5DH+Rc/D3LVpmSwDltFdJixxlLYJ0
QRSXaQLKV9IYT/4Kcqwsb1uEBZqR9SKDmyje/KYd9mL7ZocRFlJSrELeOvQisGGO
Rp2TTYglL2GHxQRw0lkfpSL7RvS3MmlFZYKmVMHa1hk1FhSW+4gGRyTQPDLy02K5
3EblnsmiiXa8D5pNDOGXLqzUMo28Z1XgTXz3Hoy2tckEoDAo+O1ESL4hHW/g5v2M
o1mRoMjHj/ESK9bH7+8IgCEPbfYFmdayNlUGPCPYvlWhHHukfw6wscx13v2lHrGO
NeKWay0CzD84DK37pwnTWwGllDTGlIQpG1j1OxpBSPCm6YQmBDysSis4O4vAfw54
+DZ2mA8amKYhiCZaCyZHL5KNTy5Rtf0VAO2VEo0iBjMXjBrJn+oZaoKvRzQtxGWe
rkb/5Kk6/IdhM3OEQNIMiBTugym1kdE5RpWcUHn83vZm0YuIwkwUnz8W8GYEHU/r
F+IO75T3gjtN2JT4hbE63RMfd7cWB5YgVRpAEKxp3/tSDl5ylqg4XqPdH38J+qk/
trmHS23COBjHcokKNiOB56BBVRypWl3VtJiCHFlJx2wBDhfnFTD5lEfq15fJ8sGw
tsAnGI22bSmfRlde8os5+IdlIv9nt750uwEM99yH/StW3RZvYYDdMp4WG4NNK+RP
nkAlmHXCTIC3+z9ja+57bqTRJmHYKgubNVbqZuIDJhELy6FZ30yHstMdniqP8POa
hy1vhtrHbGCYOq+Wad5CSXcugesbsj0WlIDF2i0SiO3bs42MWed1mU5lhX9pIf3P
A3n95ApEXtaTXK4GOTFHLdCT7V+uLOxLpWUQ2mUtOFRHEtcPah3SiqPR6Id//lWr
KY5uyaOINq/Kl52uGhfFi02F7Kze17urk1vRvb4wNgKK1Syf257zqi73dX83cYZT
BhYsC8vs2oiTUFbZYJkZh6Yaxn7JS+Hxc5pthTcHwg2hkuioI7qUpTngY5+kyXzF
7j6b8Hh6NpLl8IniMl4vyey6oXXZJUU7mldL6a9+kwtF/p0EdXrxCIGCDoHX2aGT
PFbEh84aSr1UFd6jVJKg2OAEY0jdV6m/nMn/d8elBKBlK0URVUCJB8/N4eFPZsga
8bAKvOFQOD1a+le7Oloueflh02gHGOlQ64vd/KtsXLDgOWzShzrkpgPqJvEGAV2t
OdUpfK6hx66ejrara+vOcCZjZh62FsrdaKo5oCvHNuKOE2jZiigff91IEqStIoKm
Kz3P+Tiv51h5JnBPxWUt1XLkDx7zMYgjgZdIzKYVuBVbggEpvb4fmDtmc446ndBz
fSC6qZWBwhCivTftNCmABr7UKgehhqroVRpgjoXjD6TcjjXtINHSGMM7k9udIB3X
e4txjzvKU5FFLHUlHdPCKk5CXnvYtNmZNKFsXPyeART33jo0wa3BQCrDWjcq0n2V
Fgw2IuAvKeOegK146gAvj3ZQDTCF5mGwVC3fS9Z+JuGi4oKEbhYQECjfNsxhEkev
elrT8/7mKjbwE/p1h0WrmxS6rj3+dB2bsKTHfU+80g1qeEvOl1SjQ8c9OPueyPpe
kjCZFTcxCJinuG2asoVt91qFrCkmC4ZJ+lcNlD2tjNzLybDLYCQ5ThtHpVdSwixg
W885k8WeisvAh50SIsQSm+i5MgAERLXODREXpNw66zD67fk0JyEWZuDnGiqk7WMw
KIXjm0iYAtzBWMXRZ3AvXQBdouOFpavmEe4xG124Gymh6QO6Vend4GKZ/noLODgu
sdXkH2CqF3RYk+IbARrD6UrLXe79cLCDXWW1O8Em1zMl07QsNwrJz9eEN6kvGwih
mSw98pMrBRXHN5ZXALq9GUf3/WlPkW8BPv0iOdYYxqOcPM3N5J2OULU8Jpjz9fHb
U0LnLBkJrHLaMER+GzF57iq2QRflyQHJYIo8jukwO31fShlksG6HTTFsj3fJQ213
6PYKOiJGibn+bZIsWLpcV6y6GcotR9UdcJcetWVbj+XXDhexKePjgDJ/sdSXZPGE
xEaaiiNSdVkuNRIIZ5n6F22kE8h7yrnqlJQeft8QSQXx/iMaZFpQVMr0zp6IGUKh
phMMa0JmM0oeMIsOoCG0igbcCf7t3Ar7l9qlC87Em5zm5L4ZPtcbo91+OKw9Qejv
fxkRKzUO1AE1ZA22WfhAbLPPoDTM/clRvRbN4+eG5fYYuioDPCu373L5NwCGxbEv
91cYq7YtOkeqF4EcelHQfM9CmQcgbAnIXq9FP/EvTGYbu+WvhE0de73gtQoOCyFq
Z9QHiXGf/gc9FXdyh6oHq6XkLmL4BZfSlVruLH/R2+py9BAMui3D3HCuRSONxVop
ckRyQyiMTyWpz7yYrGKWBcgcZOxuLO9zYD1sT5D/DVbIAwbCaaI9yWnVG64P9cUv
RA645wJFaEMsLt4ytqFn2KQV4FbwRyZpMV+5fuf7dt/OTIaLa6DcUoSNzD4S7mdp
emYELATqjYjYfNZEx/+vmKorct/ni6GbxqY2I+DTfbS/XL5+gq3WhYpWyilTEwa1
bZyI6DLX1s25TA3d7AHJv31YY13f+RW7jFuZCUtouI8iqjTxbzji6OUMp2RdVcgQ
xO8XngpS4F8H2Zmv9NrHNpA6RfKgGku58CmJBkVSZDhgiKEhykN43npFntEwmS8Q
N/9sQFx99dwHTZEAFNYD25pxJNMqKcYdHltg3C+YmQlJcpQGPbJg9KxnlZC2J4ua
qlg5dI58h7U9r4Lrp0z+HXXeDZ5+klHRjEI5DYzUJrDgScvHWyr7R2xGMNkOwlFl
nMdfkPFausd3izzq/WdJJeZcHNTrSDhj30XkcN6O7pXIxd9WLTStikYe1scB5ceP
sMDp50n87jCJaPh3hyVO9xN3132scpTkwkuJFf6WNf6LzFBD/wAnpDv5UwontFsA
ZhEiKBr2m5e7oh9v346h7MDzrp5Py4I3TqcD+y2UJh3nVWVMuiaRpqtaCAkUKUJi
VyUhGtOVgXOzw5/DIlSncqRkMx45tyX2GN2hoM9XUw7lSKgObr2Zf6nF7xoldZNh
BeLVLgo0qlfVf+OITMH1HUX8XoQHagYJ9IcFt8Ko7EtqIOo9/D911cjCAby8KevP
7bcJ5JYNIpFg/1yhNNxCZXYT3eL6gav9Fsoz2NgVHpuNGgZQaezJvoF1uKjEWTSN
kGF7B6YMw+GJt+rx63949q8Hn2ortYUIycOCNz1Z29rCJVAt4UcVbiOpj2Xelg9G
n2fAmanpT2rQ7Ecdgi4frswWbLAGLOtkC58HfPOb3MNZsxE26pBZkfgT/lRwfzP2
wRkv3QiMes2ptrikk/e3WuwOKW8vDMdTRBU1NwmpmN+IcYQYXoCGTqSvgt+Vw/BJ
1m6JNmvpSSvNn2RbH2TQoSCl40ajtMb5fC08ZDGN8Sg5UKXUDP43gmsNHqkCdsBx
6zmCnwTZf7nBj0WKQUjDnRGDDn82qMhqzxot6dz6tDSs1rbQrLNuq7nEhhSQWLAr
3OKN7Vjt4mjC4piw8linAWJ8ip6Mq34AiGVCRxDLHTVKASSkGLXJPwARHaVGCsmg
sVGs9aqjgVJZ09198aSJOoEFjiHOqNvEl2HE8FIeNKaTM6xguE/SZlp/OdtYvmaH
5oIPNzq7EMJkIQ2VK+humjQFCkyHqG2CWi5tR9oia1H3x9woo+BTKSlM40Lf3jAu
rGDa5UiBtkKczkyH99qMuDf2+uei/nQBnCDTp3ZZk4Uwr6Y5yx4iKBWA5blCZsEY
9e14hWYJOhI4ixNSt8AbaN7C0JXCQwEP70s3RoNcl1vXHvwddJ9XFh6Fif/qgKNe
yqwJrC7Vwb88F0bTZDHOdMw8c90SfaaQnEkUoCkTtASH8i5UbSEPAay2Phw8DsAB
nRNMTMYUJHT0y6pb2AJ508qmyK6f/vqiwTbNfzNscso+QQL/A/Ud/pJOo3rBEl1D
hxuyYkWYnsFQvzP0JJYPSgzkt52AZZQxqscuHCFokIiQyz3gbs/v+WMyYBCKHTpM
37wgXoSr6wRW6zaQw+UZy71KbjxfnWl0ZkEFZYhNrfaek3HiJqfK7VxKYzaUREuM
zmcnuLbUKRo1sMLFGA6dkceeRjlwO8V1QoJXbfif81m36xcP4XebWAkZbdQvgRsp
f0SakQoIZ2MusmRmT3teXYo3j8q56wmZLC8WVu2dYrq6MqBtczOLZ2a3o68Cm8M+
Egy5tC/3loAuCaOo0MzGdPiJ9jPnprOjhV8lIK2W374+16tl2AS70AqRgnd+I76t
67+4yqIFrY56Q1FjuctcRUyoNMGj0gq7XudCto8na6punEJheb4ml1+XPVAADOpa
EB8uaIKHP/vm0Ho2lvmbnxJdhM69SpTBFHEFL2mEle+6EPTNwgP2vKGEtzIdqag+
jtOsxFTbHIPii7CxwMQIUW/XLi1rMaUlxrYwL1idveeaKbETVxW5uTfCl/cM/yU0
hHKcgHB/+LtyCYseBcxYt/EFnxbDS1vSf1GRqacB0YBbcAe1g8slZeTcnDNnFptk
zISllTxmdArFkujaHQsw1vWA7Kzy03fkhXA9QGGGiLC7IhjZLrPA8Y0+F44Hy+yb
7wvMeHNB4S6lTBn3OsL3xdD/fiaADw8oEP0h2TPGKGfQmggnr5BVfxk7YQHRYa4L
ah+asxjZiWwg1OpihQ2yUWKYm68/OCqtiDGoymxo+ZD0zWGoQazo4Il+6qUVUrpi
18TCkuKWehAiOmIsxGlmqrOwz+SI3/gkoQe+5C2YcWTZ0yLLSLwf4FboaQcmnJ11
b5csbXR5ocs6ZIcrRsK0A4yDPrvQNw1457i4lLI01AWtE1O0p+jMCBcKEjAskqNw
VKUmsQHdQN3T9lsxpwTFkCPiN6byy0+PmJUhOLN16xKDGW76JVgW7AXO9JdeV9GL
izmeR1O+0HcWQmh4rYeYf6br7HaQ/lY2PwK3Hm9Rryd+eGhqumzo5UfepSUirbOP
LWV7T7MkqPzsb8c+vdzrWIyiQLGq7kDvuJE10trhMV8el3plK01rOAFRpYUv/bPK
agPen9PTNoQa+fjA2vxLNwODA8KezZjQCHo4DmlJoOa2nxWdV5fqvng0y9kEvYxH
q5xWC3KT7rVrAQolnCLa6i34lSNybvyEmOZKhACjXPV+J/ViP4NbrGPY2dB9P1eZ
0nR5oZS3di+L12w7OsMulp/4ttyC1uOlChExtWpByDie33c3WqqTb+rT3O1mhwFG
g7rPPz8j4FRYp0/rwmfT3RbGlyK2pY+k2UQXZd9FZE4rNvt5bG/r1rdSjnAAadbr
3i/pySKNp6iWxHTyD5A7S4a+P8eN++imalUjBdPgs9NArF5UUYNDflHuNh93bXl0
+KVxDtYRCg2XtdFTJm5fYGs7KaJfQZ2nsBdQN7FntSmPoRvOIuqheVICaHMfK81y
G8uiqggyahhMZwy1hKfgmVkguRV4LaDOx+BRtbj8Q37o6zGzqVGCiGjeelwEYn4g
d68K5II67JO5WYmRfdSupZ7c7eEw+7rJgZ21JmSK0ZznJQK54ZDR81kRacKdGAG6
hBC7qFZTqsz6CSmIbtvHHwHZO8Jhr8GtqyVb0J19A6N+tSZJdxpdFerp8fZRP/lx
tDdNu6ds4u1wnRs0ITezY6+LRJrWBmlvBXr1d0JebU9bncfojHSYFaCy4zybyMB+
RLY78OqCPp+/yNJmgq/5RoCDfNPJNp9DassEc6BCvegK9A3nh02xpmgcqIKHazGb
ZcIbf+X58xcS3bvfk0HbIr5fmNONTxlKault+UISvaW7ck0mbhWiRpuad66l4VKG
8H/umksFtDLaqzRjA0181MAhRxRbA/ObKFC4vd4wuNWAZhahmrvbvNOgQiuA28Y8
Z8J1f2YfPmQaLq1wQqbF/CM1RAvxhIZHU2Ub6WP4GhkDti7Fu6axStQgyuvVbr/u
m0roWmfTq8Jog0Gj3uS49GNI9NJ4hDV5UkUfIfNPVJDM0NcCJHxwrlP5twT1W7WS
2wvryp2DpzvUn2Y8H8inmElFAsSJa7ZGbUGx7fMOHV+MrvIg/bf+Wx4sbfH3pUJC
EbQVROg/32moJBbvkmTF8otwL21HzELA8jnFBpfGhKGKJuR4g8n0gqhryHImdv0+
cBOa72WATkxyir+Dp1SgtArPiCyBT8QOK5SEbHcedrAYkfnOQGXglSBzoxdwoP3O
pL67mGVAYZ5FX1qLuVU2PNAVs9UycWz2IcTtIBWzkK8rKrre/NlOwTzQEZHWGZ7B
SRLRttYQt+xxahKyb1P9EIlQEqJV/yMrmqDFF7AWBxKPSTrxyARAxJfS2v6s95GK
IqgR1oH1NOJUU7/l2I6+OVMeIWVn0avQ3mLi48NYyjHM7BoYuHqTVwe0Dwnhhequ
nMm3nh+blMzMK3129xP102vKl7Fh/wBKwsUKHbR7Balh99vIN2CUDKXt7QB7BJTP
Rahk1jEoKO7LXww9xzrbP2iHI8PVxMiBHXp5h2+zS3du2RuuCxj5DNf52d1JLhYk
PlApQvrPTnTmP8mT1A4qe8Kp4gp3TDdCBMipdGlplq93rP/2kQ7Xn+THe/ILGGfo
cmva0YdB9VOIcCBVCs1TiEZXh/2MDwapTcnWJs5netH8zusnGmhP859BCOCjUDma
yXtDkLeUGTW7Ur3Y/zJb6VA9QJyZSbxUCSxY3UkZqsJ/3GbxYVfeP6P74lyBQqbI
6cSJ/PerLUJ3l/KCv7e/q3dTygNIxAAm0RARdVFlA4Szy/Xh4jcR5xfq6yVEYwI0
1x9XI1x8yZwD+yD3ep2wVroF95tdq5xVJuoyF1BV8jN3bpP/VTVRkofCYnGdFiHN
TibuwSndeV1dg/uHj3LyDJ/kkeh+tjqj8qEXnHt6P/tjJlySIHE9Mjgv9pe3ERcP
NobpFOo0GgY48PiGhv/gxs0xcQ+NeaHreQvBH6msSUvMN7wSIxx60HBynHb6DzFB
wKgqjIRzeztXBgBeDlphzzGnStwReh86x1PJHUure94hOKPDJL5V+C0Y+eXW7f97
VHAJjtXHq09u+qlG0o/rKwLrFQ2dNj8JUC5dXSo14soZUtrcGA+bxgZcGMkNwFa4
4EJ+TumCYAlpSQZRF8h5kN8gXuzzJ16FQUqA9j1/UAhV4v515kHWp67whCLIX9vf
OKdYsBs3cPDFdhGLCp3fDN/h2cFbua/7jE81eOlIu9wGIGR/iBiy5qKzqalaB5w4
oBl5/8H3kUC4+I3tHJoYWYVdDk7Cr0AMIXOEulXXARjEj8kDG3kZVZPaSvrfI7ld
BSfjUFTb8F9acmYjxi5DPLLDlHQsjEBCR+itsVVTmHLPF3iBwaiCuzCn2ICa1tMQ
xWmFxmXfR+98odVNi6G4rRdMKVEobC5zEXKXXorNxDO5+m+H3jqQIR+lltU23bEZ
NlY+32gAlGC0CnaRo9a81FjPDnlkYzKuBdnCKAIMCeKG7wu0VfANrpuGtel2GeIO
gsY9dxIwuLgTK3y6xyBpY1EX+tIv7GSLjQANLCbJZPHXv6ZpC03TFTdqTmelPN14
7z3IaHv9MpEyunbRbxtrYjn8xV1shVpoFfK5teFseorR/MVrVb7uRPFKglVid+vW
0BpWKu2Yl66wnCro5vJxGbK0uehC2ubXl15Li4QtFq8GGCPKigSG+Y+YluvB5C0a
dxw6P7IdqgNHBt0ExRXK6vfFk+Afwqgd+7nWUh1R/K/eFhM5wLzgJz4pEg7ofhGa
AYw5+MrtoIWXFao6Vw2uRj5VQZDeNVDnYp3UqPLSJIa7K2FruCnyU+2K277wZM/P
NSU7F0yV/Nv95c29K/H5bXuy990+0pEqsPLZUWVxiSH/fzKH3ivEWSUXXxFhmv6U
YIq3CpprDzWsDaxFgq0c1r63Pncz5KH4dEczMt5pvB/OAA64GVjpoCGAWW2ITaD6
gsf/mq70UQRQFRFbRlObLV4x0+uPv/qeoFJRqkKg5KGTtYR/flOfEW3dk/XCkkWa
RD9TCUwNv2OqgctZyJknKMi4m8liACxUdRyP0XzgQkGlFD0RCb99u9aEpZ1Fmudj
l+gpancAM1Bk3CjQT+xme89JCKvlzOZihm61b6XTkDXbPWHPr1xBG+De8Q3qqS5y
VPr5ca1uW1RJ/vQckXsVv989xcA6PGSD0HjTjbx+5BgLd9Ancvk6UKZBYfGQgTME
ZmNUZkxijsWosoYDshlrt7EUmjYxsvk6eJLQX7j45rKh9ZsJg0mwlAlmQvbl8fhg
z4fNz0wgJdSl0+qQzQifwzsYInhFld7y4ffj3EIU4EGzivfTPwl2k9OmR+geQQ9A
rBJzPB3KPay0tBbx2ycby1HpZkTLh+1rrqi//AfGwaNvsFof1+zV3NsIe36ZDILA
zqDuQsQ8zm8tOMkFsPKafWF9srp6wWPUaE/xLEwHAEcQaxcnyP0Oh/2P3XY7Ao2/
v9ee8rlAsY1QOS1ftm0+iwQ+0OF0QptMX2eVetji/dfc3ueg2rHRnNAsUoFqLJNu
4N38pFY4nMrBDow62Zo3IOFWNWZhNIntE7lU9rv1ROPLRUl7CFRFQMNGVpJ8FhIe
ZhwAt5WqIlszFy8VZWrAHUCPrPvNRDJS/gZld/IQpOV5S/wmtqtJd3R2/EOxxwiR
TxULzs+mbbMWFr7z8XssbUma0vMFxYsP9WSe1ZMrO6s+a76SlWxDJ4k2+KPBUdLD
s0HPfxR4nabkcTBd2uN4i4nR/kmJN8eWkT/G6I9W7OWmeCgTnmPzZcMLQnpP9wg7
gMsVOntNcWdgCeXztGq1blereKQBx7H3NhTKPovv50sorrNiiSofPC+rGO6jrrCv
UNQyD4wfUlSeRojrfxtZ8axy/jLStWfkYmQOecaxQXvGjqDIS3f2RSon7l5gYtV1
9HPM6F+lLngwcYZJpWIEDONV88zpwKHJbYtJQW4bQ4BylQmMsTaX5Y6J2HQE754f
wUSD67ZA96kThhBMz9KVXDhu7NbzAz4GolrtsbHUlqLeo9KcvEFJFnYPtXd/8ULR
DaeyfEPW8QLvpJuV0feKmdJ9F+N8LozQ3OA8YyGqigygU95RLjLGXQ9x13TP3ctf
OzFDaYCrtALXDP1JSk6jHZD//bFiRvfCLzYHhHeyG/3DS+Zv5/rnaLXdVsqWdGw1
q9eq1f7cZGpXyFvJKo6pRgyFMyEnioM5at+s8pVzDlGMUKdkISo7AmrRsi/sYzbx
fEoUQ4kXfm3DFNR4MhSnZizVelKsvdbW7qFb9W9oR0RQznmlr63L3BU4kSSWnW5Z
1Y3ZQZp9HwmFDFmsLi7qJvLEv2Tr/AOcUhsRApZXW6j43lR/4uXXpXY9noSEAJ/3
BhIyESmkS6qZ7NexuNhR1Oxf7DaiZujKLRJ4/RwY+x9DCLNXM7zJnJPWmV96NmPa
Noht40vLR5ADC6R/uPbNudLU65i1AaOdFhep6gOcC5veRHd2v0uem9ZMx07suwmt
NwpDmljo1NMpNr5mIGvipu9HcxF1tF09kUFucuk5bI0VtrUN9AwPnv9T2sr+aaJR
0CSINtT+3Vn31Vk0A3PKkurQxk0KX2SUXUuANehqQbJEY88ruFXJX59KYzBYISpi
NZR1z4DPziGyAIFVsbRSgsEf3z7T23Y7s8FAkufLTD4try3sGrgQqKK2763YPmC5
ijfn0rPc7oXVtH2pTrqT+GL6d4DIl75zw29WXwwilx/Q1a5bGPJ+97WTSWhVYwSA
n7C6CvQ+4AoRxxOE8TqDJ19r6mLfWVEhkLNfrLu2fEHAb91A7g5DMQX+EdEKly7m
ZPVwFpb6ExF/85xVW1vpqriFSD7CDiqj660kdaLTDy3k7MwN5MI0/0gxy68a2c4k
FWnIvzU0ym9R6nTN5QJ07ffaIo9UHXCCHUdpP3Nwwb+npAa93NGdBwRjiVURobf6
Z+A1vmkT8y4uEcUkyT4+vu7wFejlMrmJ00XldmKvgh9UZuY0eyUAVltujmDWOmNq
TrCNseogsNDoTSW3iIQ4zTO1773sVBmNmWcNEXVCLhn/PVvR7JLKJE+3It7LGJ8V
8k8o9CrixJHQIkp07r+bjzF6gI9LivumD6fI/KsCID3bFBoo32obRi8lDWxUHjyq
71kuIZ6RAROQZQtaG6LXW2fjJFnOaGFmmJA5I1k1VgVcrzYxAw7g+NQEknNyU0BB
tEA3AWk/pbhmqUib8WTC/aQpvxOjNj2/GFGLq+Afbf6+exNcIF3W0aKoPwQnmFvh
wjS1qD74hf9zNNOAm0SmWuTFBDE0z89I3meL+YkkqJa640c9GYKc1ZlCg0KzdE8y
gA9OgTYtfwb3MzbrWoQ/8senk4RU9N2R8DxoQp5wXZYfC3nbOiB9jY9ZADbtSalb
WfGnLyxlims3KmmwQzplFif7swJn1jgszcY6BYy1gJAb2FmVcPBRroCTEWCUT9se
pPV8hkDLcQN3ocwVzRGc11Yc5x2YBrdREu8reBNFtq37WQ7RlG81vZu0fZouLoh5
2OhkoFgbtUXXiCKf2lJvLg/VwpxIPawpBxURnLLHuhaUzEhyIZXVW01eLFj9lRPO
RdO3aYDq0Af/mFDGnSMTGrXPZDF9LhCLJRsXhLx+A4aTtppsR4yBqi08rtp0FArb
cBvqsJRVZzG/pEwF+yLZgC8zVAluK/oi8ihZMSCgU9YWF09ztuujgykikiO1dHP5
uMQD8xE/RBbaUb2nBdFiNvStr4ux08zMJaCAVi6EfQuB3eMJ6oT3b3C5WpM3goy/
4LfcfJHX4fTlF4yqvD+Ye3PuL2D6eFMkhL5Rb7irePqY9cc74/WLpIMayGa0GJo0
LI5MscY4IIY6DReTJIyT5Iba8RnJtBakZfIWG10QFOD/5/a+BYGkNcxTYono+BIO
FW1CHiYvoiFlb8mz6dyV5hc+ud39QBI0IxhLf0npKFslshm8SpUq49gCFNs5nbhP
DLFOxb5Z6S4FEm+7DLTIbXt67/85bbJCzAdjdxTar0aDC3qvBtmLJghBGdBv+ruR
sUwTfSP6efunMtw2Jc3iyXrmpGBTTBeg5h9fqK6IXtG+snvs7HmD/0KnEkUZZ9kJ
/l2D/8rWJ+HZKGpZibeAy3m2ggcTh9nL7FN/k6CQVim1R8Gj8jyOs1TyOyt0A7Lv
qzDzzisFt73ItF3gK7fHCyYYdkA2ixe4fYii1h8YivAekSJRcKfg5EJYCgwnvT71
grit6yKL8CqF89VXGy+u4WJqO84M44Uuadip8AQTT1iKR6PuPGM5c4EAB4nCdaVD
ByzQfnfaO6QfHov5f0kbtiC0oBbHdWQG8SzhkxlvXIcyfxrC29rtsDor0F+xMdCl
gXjBxurW68fp6fvRoDKMcyMLIUW4ySLoHhz2KqzQ+NR1QLSnp/nRC2VJ6QqkSBp2
YhWPmSwHK1AxDKZ/v4QEXIt6pcba+tDmLy8QYH3eccEgVLQXnW45/NZ9ebmkgTnM
yz1/XKY8SY3SDS47+e8mviKMxt7FaD3AlHK7tA88gAISYGSUQMxPC+IuovxeAe43
j5GxpheaenByICMwioo45kwSW/DSYe7uVfDkZBU56lLR9x9J5e8LcP1lY6n75nvP
hsYpD1RnzDUcKlm/oeKXucf4s9bMpTl4pL+xyHZ0FWXvRUjXON2/Y6OiRawUXp3i
POH080Q+WySyYjKTTix6FiaoUOGcZTl8A9scfI7BP5rBXYqAyUSPKxOaOOBcH22E
8sE7omir9C4y/XNTSDi3aT8feWF9EHnoAb8mHR/kX+QDnseDnyd3tG8q4ZSXRPGr
vzc50GvWqKjhDB2xzBBwU9HezzOQEnASTbmM0sc0MCgF3Bg2LMX0RB9Kzk1tTYR6
cORcM9d8S+iTXA2xzBsfmeVN6z8H5pB0TVfQXhpnFHU2hb+ZGgrhuGJqvTLbswFg
Eg5Fw/fatcmonR75HY4kosbp+haLn/QMVevNSFqVvRLatyt17oCfealybNlZzTqr
EdEJnqGPaJiFbC1w0yH5BL9fIygcK28z4wn88hEjIEUNi200o5tzmfhB3QOE/Qhh
EzoJUptSeUTrKnqpFrPiOIqdVsWS8C5yG31RF1Hvrv3qmgjrv0ueT54PLrK3mvXg
X65RFQvkoZ+xgHKZ5HkT5kybDRhYJjLLDQrENqP4u4KajtgHpEQQx1JVYSD0Jfh5
x4kHQgAhDDnMSi+J92ahgtAhs8qkj41IOrV0iRg8qJAgCYgxVv2E7BQ/kUhs5Hdh
kqMpURVmwZUH0gAdyYSB2OtA+rRX1KxwdYkWqzUj36ckQx7bGUhLn/HoQaXrEaJI
byIrGcJn3M+64xrtExgAJi2Q/OtNM4h4sD7JaEj+XkIeSY8Pv+D8tBc3mkfWuNAv
PyeldN91AY+sW7a+tMtcrSBcCEMeDUK6DQJ2Sh+Oi0WFk4eoo/PqhxmOuWT9+S8O
N2mjpVJyZI6c+H94qqNNGIe5wz7wTvOmrfozSbaKU98s15LFQ/NfvwfuJrO/lRY8
0VpVtpqD4n8rlTniKPi5+SzD6H+IfSKpkVahm9orFPnlnwJjdOvCRY2yJN3CUdoa
6/7iII3Ybnu834n2dv8LnLEyLPaa9x30T3SC+FEph3KMTrSGfGSZ3KOtwJjUxi+f
Wn73dmpi7j/RfN3hEFl4xca0cnOT2XiQyhltjWqf9SRPB8RwPZSVQGb6TGOspeR6
PYA5YMLVjY1KPb9ZCeHQF56rGBLcCIvxpr+Vxttd5BnT1NNqpLBk0Iy5Ddgwiz/Y
qwQt7wOs6HN4prwgOTo3VMinHYx3qElp1eOuwYtFrCh0lInEHcteyPgbrLI5bxE3
Z7pvWwHFO9lXt/DWjZrGUe5GptGEvfm9cMjI9cibrcHTvUjKtTzUMknaif6IFyO0
9WkwRbp35h0V1hvTB5ErQyv3O/gSjE6g/zy+9lUc1hnFBol/MSvAVC7iIEYqLWWw
6+pXO8IzDxXx2L8R0n/pq8kTpYy+owUpaN6MI9fjr+QXDHC5sJdYknrZFh/3UoDA
J64gPeB1ZX0mkodhXrfrMTbpFVu4hYVwXIKrdhJ+WN/cmMQKU+pQKFEuU8/Vsl1j
ZSKASoiD07Yd69WvgPdKik7kET0OdqfCjD/SsLA1QvsMNkMAc6+rRz+hiq8cwY1Y
FMXSShnslkdx3TfClm8kUesZRYrqMxBuQ2mt9nRfRrkAPfwOaFfu1bHg4F87sMBx
pIs5lCWUJsCqHC4iHrTO2NGjAPdiTyggXUgQ6JZ1743I0M+pRZLOS9EPxjFHiKxS
LMTFoci8jrlFOtI7BzhvqXgDHuvuvSJ9aQye6vQr1He9i2YIxMLkuwds3Zq+CP4a
9d4NlB/XpWi8HVUX4+W6idZbyeo0IFyEjwi7W+yF+s0sDOXxz1CgOk712g0eSFo8
+6BzImNpbyy7NTz4itujiRNr6UHTfkX90dFcKetrpqaO4Uz1gygPpe2+q4fSbjnt
crNZgl0ZwziKfE/uCan4NqUULvmTsi/S/JEoLrMozu9SYeEolp6nCuAM3enIEhUR
JPzo6V7jXs2TKiUd9LhqMMLrpy2zRBRh7o3Zo6uzPKs+ZVvHQxARi9FksPxwob8M
AURzOueyVORfqIn7Mbf1boRso3vwosS931xi3iLGaHdG1FucEBJvtq4nDF5d5xOJ
07yYe3b7JoFskcfNxmIy+mJABsfuA1xkeI36SxTCrAkb8rIqGas/btuQHhHl5TuK
gYSHftci9uzdag4bbrikAFKzwltjDYRtP7skqt/UDvN1esisCuWN2PR7vjK84RYl
la8EaKo0J4kDH4pensEZo86f4C4uw7Yuw6dYmI3t2Q+myzYEepdy8VNHEbXJ+kAj
mEjTpZyoTY8djsWsE4v+h06MJE4e3WqNeJHLIc3R/hZiHQ09NxhuBW8bI5LpHYpq
Ay3v/YckvM0YqnWuoR2AvTV7dIVTV5b6G6rcDcbwekaQ25PdBBR4A6wRcIAJK5eC
r/yaR7Thb1lXmxXjb/yKd1Flr8s89LDzW3KU0OnQJHzsHJ0F/bfbzJ8a4aR9zKQj
B1wIbIL9bTT69QVB+dLXH/ah6i5ol2OrLaY/1Hhhu1ib7CjMWC0lhHX8Fjr/KEES
y5Cqff5oMFgMzsljQc6NrzcpxHZ5fld1MqbWHKRvcsXDyAdmoOs5LKPs5uzTzinb
4Sois3gBChJB2uItBvqXl+k3jNcJeW6pwj7Y0OewmLzT4I+1ztijpT7i15X923nK
UlhGWaP9ZzDHfBkxKDRZrck54t/K/rb/2MGWGm8YAWljE+dqrs0rBYJfK3lGYQjf
yMfS3NW9u+cuYRZKKFHM4jBrUuu/mqw3RJVNSTwsgWhvAgeFneHOdF8cAuGXbICJ
+aewkv7rYZOFnobg3dVvCpknwbBM/os4OQZoQ0ax+2Fsdn46XL/T9B5Wc8TOo5Rj
ST19VIu0ZlCtoRLVxCoRPaGR2zvJNdSupEbEXxVoCJtZ75LWjzIZnrtmFKMunOFj
S7r+yuDWZA7K7EL9f9u1xOQEK69tlEiPl2REzHs7DiKL9B0IiZ3AvF25rUaq4Q+L
E9uhbJUf6p4mawXGaCtcW6RVTEmta9TnTW0FKwLO1VpoLAxIx8Ihy8uAkKRHomx3
72QpAmylZPoSZb1MU0qiMl/8Wm9ujn+VmzVCnpnZTRcHs6dW4B4voF1TLoS2/w/n
qKvUCI0jsBbbjFD5FGLuHVxKbq5BMadqJ/orDfw7WazrTeT2jOHw+QOmcS4pn8/C
AhnmT9zKaGwfw/G17xe0MH7HoVckpBWyexPCHV10yuAPrYjsC13WiOHRK7j4WewI
ih1KYA62+u21/y1DinmfXzJ6pSVbBJ7YTlac/THMddVcc8wtoo8Nh5YUB8BzLvEH
lqAgpoh3pZ5DIVvq0IbSJLm7mP0pC5I3JxE1hBcTXzd77nSUyyjS/jgWP8RZw9gX
CHdiOiZyiBsEu6T8BsC4bb4mZpFoYCA94HOh8Q3Cxd9IHvCGTWbLhHaUorNU1tVe
A2bat3eFg0laK/3OSZiXalMUjU18+6p8RiMDJDN1FVpGrlxrhjXBCoA6Fp6tiM0l
r6c4cdzRsFusm4lXnwVvHOJS4en5mn8BEjQCazEgE8zfqf038K9BqmQzlPjommSJ
C6CyAAy4DdXxq6BAR46Vkwq4Ugx4GoxnhfvNhmP0YDVho1W4nJDg/nRpIIUgM4qT
IXoZiaWh6Ed3JEzP8yGvWYKfHkOcvO2yAaqsb27ZLBtaB8azBq/lfQfHZLqWTxqS
Reqr83bWPyYMY98YG/E+35SfT0ftOUHClU34OdUG+CclWY+/xYZSxjlNliLEKqNE
0g4l+T4A0ED8g73H0En7vDh1/9xQjZzUT8DvPW5TnaLxyyyKgTi92XWVCg2wIt3C
+f2VowSZUilSAs9GYGOGCLN8qfONJuKzIBQF0IVj+KPt1vWU+j86NCT70DxTbzjm
FmrGydgc78IekT2VYOwXeqellM2+e29Cqgsn48o0fRGpD9vkZJskmvsyPILIHOTx
Vq39Kw7LMZlgOzXm5YYEE7ZwS/HcSxMwdg3KPIU7p6VE/gX5S4klD0H8fuqpKnhs
5ERWnZbIfCEN8vAF9FpnAai1gABJZq1IdJE0YaKbjLwoE59oiHepL6JrVBFqbK4w
Th+9J72/NXUcJBd7ekBa22MsIAmLkZOVkJLy+xS6vXeigiU46gHrtTadVOLIyhdo
6XSAAByHlxMb2+p1Qb0NDmmzOeWeGSy3XxrXAw1GYaSfaPC9i9mAQL0ch4m9/P9r
nQUXE+kuKpR0TUCMF+aPMKVor3GV67SPDlC2F4BO4C8c7FJatNn6PmWson/Hzek+
jAYxQehI/9ks83PeReR6XJGa1iqZ90WpbonsfCHljHYfso1GJR4EJ4OPtHD63+7Q
mjFms29JtKtUiSxKqu8Pc3btjTrCSptUvDgVEyw3crSi/GWWdW+8hTQ1b0pGd0YI
x9xfYgBcSMDd+IsMS6FbMNW2URW4w/UD2GIRSHwityaBtm2rMx3jXdBC6NTjaFpP
Vk0bVmwsY4MR8EnRO2e7cBKlOttNBOUj+nU/im5qenhCSnI9p5c6q4j5caz6UOU8
QSC9BL5M0vy1Wk7s15laIATJmrihUVBQ9ClIhRnxkrdqh/hHlvumYsXk4eh7ZJdL
TXev5b7sSBTACCl55Kt7pHp2wxn4KZbiVOlNUREv1ci7yJ/RF59V9n5m8KAwBKg+
ld5fopHCemTc5JRDoynwrh0BQSZBTIsEQ2SsdtBtnPwUqCNpMSO8uSMgKnCZj9CO
mYGRVWIS9UlD+gJNivkW2frGrPrfOrJd3CfwExTueN5v9a0Qhbrr3UqmBBBFI3Gr
lEOrbClZZ5CFYFHJto8Q2jcFjagxt8TIfEJ/q+MI0BeoJyfzc+BwhM4lqlRXZ5Ps
hXVvMaTqwfHOnu8X0JbKR1Ybi5yoMCiSezCfkBdyVw6NT5tlmfH0lhwQGfEcb+ar
2ZME4teq00kuvaS0ZNOODj4G8wyYMazLW7PLn1mISqHgnNvbv8WWpqJn+AHcY3+x
o2XrsGItpbZj+w9/ODcWHmmCSTiTETt9gW/G1fZk/FpaqJ0mhvq+t49RnJinlHFv
gmFn4EmltENu+J0NFIXiL4QFBrz77vwNF5FXVabI6gPl7DNdGTEtA7amXOoVuDGT
gE3TvveUyelm7hujAA/J0tpMDtJa7+4DVHBU3qZ/yFk1s8/3vc8DTtwjYiEYmQtS
zdq1rCeSFLdA78ZZmn2dCWcNGcZFfsF7Do1WWbJhbSkaoSPkpU+W/fjf4kzQ+Msu
4us56lNUAns9HqPcq8GP/cpNXx88ypYqc/FvYxrIyEqWGMbiZJvHY97Gk3hX1DqA
8FmwkyH8iNFHEZTMq9ZDkKRBjIBKISi4b+b2DmlsQb2WTPqWE7jeSlFwjl3Ee7XB
j5luKv5u/wpu4xQt7DMpsnboni/E8OBPrsjEHjXWI5+j5lqtpljRZdb6YSJHSgfw
XDwkwDquZpUIpUdeoJ/EchZVEcaWkIuhWRVCjGXEcVKFqy/mjHZvSXhf1+2pCd5Z
5KMsPZpI/xY4LHm+ZuD6OptVEf1iVbXWpA19XWeNsLEShXIDJW6Z/dJRswSr+qkN
aK2IR6q8OLEeJ98CJigAgiKNXNYKVtlntiNiu2PQO/iX4Yi9V7aPy2U1+gUMUf6s
Y57BXPEGfQmKdzUqcyokTbGSBGAs+TBWsUxbwGBCFbk+jvsOtnjfBBt+/VAOtff1
KWgx7GBkqX6fYqTkYgXKqA0Wq7S8EKUswhS+A1ofoaOjtT22soKMZjlOE9IM2phH
ZtyD5RPX2chinqzNlZvIXbuWMvieQ2mffA55Zbw6GGDnGOVxsJR6oltYv7B3eLlP
TZnJRJfOP4EWaCB0URNrW5sl/lx3p4g1Gp5kj3zvwjYn/IEEKxu1NfzcFxbKV/3o
C/px2FNkSEtlzxCvei1G9QY3klwL1PGFz/f79f7WLOiNPevIaX6KyxxVjVOWF1u6
0clBUt1QnNjfxfeo8dzpdkLGtjNCSc+yB4JDrtTuDw7ZwwsldYNQodHEkzElsv7F
Bl/XUfZ/7TLkcPURo17gaMNFsP4FqR0FW3be6C8pd9vPxSpLr+3y5VmYY06sW9SS
2U/vE6VHr1FeNK6BBs487dwoSxuIqRk1vPxVj0u9GN/P2NjoGkc3osA4OmsqYGig
vjRM01DpMoXSTulTMJ27VrdOfpiDLmeeOKoxOzUYwY+//RO8qg2ViuZIlgMtREPX
oBGmRJQZisIxjx5j4MXXtrs3IXBF5v8/BaaNoK/87a4pPlHMc0S8jZjOMeSBsCV4
UqPuHs21za9mJQaKecvz53tHnMJ27yeVaK6NGEtP99hS+5XojH3i9XPRe7QeUZ+x
XJu/JlJSouonf/7N+ih6NIOcAOrUv5bAulJwBTspw33PWhDRM+KFUFHCvb8jNUBZ
e8px79VMzFR/jyY9GNuVeZlkyLR67SLRudZf4Zp1iFGcYGpMFs1CVwVhHaNpdgdC
HRsCkSsTWX673dQ3MNEcwvQw5+YNQsPxC6g37U+Ber8beEHLI5zA/52KRTgW9+LP
vq8L+z/K8hSDb8tf/lVeDV04Y8smPWf6eLVUuaQpPlbn8rq2Jegn7Z8arka+otvY
eCPb2FTD4ImdFFL5N6S8d+L7GxbNbg6tAxMsDgEiaDZDkbOoDJ59JJbR3nnSPAmf
1wqN8W7/uXo0Yw3QBRLWSJ8nGAQdeeVyF4DCDvpL/t8e21hdMdNsI/EBUCtylvZT
dJ1U8Cr0VZkAfOmgHjYow0uiUSWzkjA+JWzyQag+MdphbtK2HHdct90gYkWOBbUV
F6uEBYkcUB3HDJhwCvUqFibysWtJzTaMfbm4ui3bYh4/oKFGiFsPNX2yExN/X88t
UA/grXmRiSys7LMVMVJ91ojq40+GK+wShOTPfs3dj1pKcizFkOD0EZ+lMmv8jTnn
/+fyrOuDc6aUkD8UGwOrNuxMgUaxuerEawiJlFlTAsaphvmhV6zob+8Q1Ct7NQoy
nbRYMYSgXoo8eWOe+3AHjnmi5J1zjfyPyXwjDX6+4Ib29XxCDkmwEKDVCgRlsY7O
N6HvI9j+HiPdGA8sb6jSzKtdFW3eb3fvdML5SUl3uOswCGHRn3l7Dk1PKfvhtdrM
Gcsr7nhw+RFLEEURnt4+LJEK4jX3ShvKAy8fX8ibfPSA8hPGMqr9SBvBMNuM6sw3
I1b5P1htxXcmms5D2gp+UHUEw3cWsSPnxSftd1i3cJLw0plE9l06eG9i1sZEgpF9
jGYKVQIuv6KNmsjpklw4E06y/LlB+4RO/tJtskgSBIwW7scA9CLikuXuPTYgYKjf
AeT7j0Zorw8At4IZ6MV9Zfkj+5EkK5+qf02ZkyPibjK2iYhLc78AXXaPc13ZSRFy
j9utnJK0JnuKDiwtRvkQ50QJ3RXR858rjFy2eL+hAMpXFGJTMNggrXEIXUevlfiR
7SuajC3iSljBJSmpdCbaz9/vuZr27gn+9oSYVtaItQqkfqIPLjc8/OOBK0X+kdbm
jUsjLuEwmd5KJKhjMyfsRunVmAPfAWfocfoFq9UtASTcDOh20CchlDWM6vjOfTML
Bao1u71nU3I2oeji8agO1+DcsphRo85PLwwG5qMU9tJcu7r73zZ/pI1hE8vv6KdD
OnV0czbuPhmaJPqhYcPN2BIC+IRYfM7gN/E5AC5HUfAXF5M5LIsv+YZzeWSBkv5H
QnnRyGzrUd+zM7UAVcAMITU7Ijg1NugzbfFfDqNpKQLHlCkxIovZGZKnS0IUUQls
mTyOMn6kxDNyyY3w+Yx6ewyJ7ZCure13pCbYrJF3VpRC4cNryBKPm5NU+wvQz6Qz
of9JLhe1AUZ59AIJ3Rl+Fnp8BBpgqZ8bJ9gPB3LNuOQtWXKKfuY75ehHIRfa8EB7
ltmDeuGtz7jRi96v3us8TUHc+qqaznsBwCcIg5BHgNZnLt6VCqeT6ddeDluE9mHz
OGKa0YJzQn3KvEvar6idy13sV2X1vSKwQ+1BeqkjZEQFUyGsSAdPRPtPeq68lX7u
1Ay2oGtoEb5IIOyX459X20o2HeKC/yS21bbcFfiowj54tEBM7+7CLeaaMdGb0lLb
E8m90is1EqTRJ271e98LqIWc6amfesWvzyyBjHXvKFo0ff5UPCzX14eg+wRqMjVn
/ygrEQy7RdW3tU3bYAhIjVPeAeDD89D21NUe0KdCs0Feeju8muUzT1MKNUVn4j+i
mya/3vBw0jNrfBdHXitEUsddftO4G1vFdCptoY+HxPTXHT9z4JHGix7PbwNAzqkW
rcyrlW1sdSGyeBb83GtMTtsjq/XyWdFyzyodcihTPWUOvSFwPDt5WASyMxEgmkph
RNFfVqjrmRoe/Kn+yDRWDUE5EUdSIrHVQAxFONSs22xIniGBS5Ot1vrSvTADEFct
qcTlTjjh++CoK88trUNRv4ia5ASDbVJ6hsqTLInOcZzoByFYmw0dJE1yrlGBzfEe
4/XfSCiBe9mdnfP6tyqhPIlldPusBd0yuznYPRPn6qf426o90Fac3Li2sFbapCQB
mBdUI21MTZ21yZYfxYQ5Cxs8drTDD/LNzIDc940uYvtjNabQpbmfy9ODByedQMyQ
UiPgFQeLDKuQ8f/zd4+nZpJeWZN5nF9oGn2x9QVj8q+vDL3KNLv+aXGeN4G/Ugfu
h7bZau8jDLl3hMqrLXg3A/vW3pyITBhkUTqKZruRbFnK0oNSFnwNuBKvs+iOlgkg
pQddbCTTVnPysd8wTHQ4VHtITgNhqc25Ki1CAu85HuORzWDrEcCdF36JWpwMNzh6
0hy3gvWTINzw8JT74+29880XQ4lA18rYG6qnNn21+LWWGiF0vUiPWqlOrA9S7y7S
nRKO5kkeUGUv3nXYmmcFP8hgcShnPH9/EM25JwzJeJiaLG11b/Dcs8wR4u0zpwXZ
JW/NquIoDo21Atvo3hawrAd7oPfZ7KjbaSwPwXJlMuxie2okXUU6OgGS2l4ZsV09
ZyKeEaLR1Y3iUOM6/FLV6YicHU1lgXVNK+TXDN12KBghPbZAdAFVzBGyekBvENlU
2FDkpbjRhl4gqDj4DlLitMmMRQhjQVAPLjYYQns8J1Nkg2lo0US1CxSCjcKwaWmK
KbzRHGGT9WeQQ+KKPAjNxPNXnmpddbrPwyq+row/mN8A2iDD8sZeMDfHUBEogHZQ
TsDGl8h+5PHLsWKuURVIPaHboprYMD1zSURn969KK7ln5qimRHRSABB4hYRIBakx
sh4Z7qmcH9pgwTY5RsiWBfwdvv2mzm3A9I1rDdWLnUC3+o73hlTAMgzWB1wH2smq
uFtO8pnFLklsXaazHIBOoBZkJ+gesinvu8lc5eNbjNhZ33DzDVVAcFHzHV9D14Kz
875XlcVypqzRsd2TWAXAsXxD5uOOiwLFsW/2U/29N9nyz3fOA0fDiRFbcJEaAhug
05KWs/p4Vs+uEBvdAegdhkJsBJ0X64EV71v+x09aDXX9rcOS2fwkSKNWu7Hq+fpn
E1ALskw84eaK/Wb4DvGLDObEcQvLbYlrqg1knX4KRcRilYuFdVdxTJokTwD31ceM
FqXkzDxw05FFV+ptymwRQ42CNsMsWrFyt/FDiwthHm5QktLCJ9peOGHBbF9Yj3wN
CU8QzJsN1Rjlvg0qV3PPWpl7AZbUZ7zREINgrR4qRvGgfLC8s6uK6+OJuCYVTjwj
kKszsL+82puoYVE+fyJyYPaXegb0CU3I8yeWhTx0c83jAWaHRGvwvLdwYbA3E5cY
8y/GX/AENsDpVM88VXuSqPe6JFJt1jtVNaPt6cmn1eBJ7URpL6C2B5hEpEAV4ibo
ygCIOFBBURvK1YuIoGNhECQsKmcGdyrhkxaZwmsUA78dZasL37lBlDAWuDtZKfCr
o6ITSshyYERHXGI5+yF5nAVZlEEWp4rFvhsvuy1NcSu0eBrMlQIS23SOowlSdvEY
VvqlvxA58ViNC5rRVGN0sNNjyvTrkQkpm5i+PzPlsp8c6gPPHq283fDbgQTh0aon
eZxCROK/4WY17I9xlW1j8DD2DrJgLsjBR3kmggogoNCkcHvB1CTiAiyc7Luxo/U4
SSPmEcTVZ4IInSaCHNDOXJPPVtB+2bMKvb/AmSefIGO+RLOr6o813Sk3JmmZD2n7
cvmV7Uzp1CMoCsY3x5QV0jkEobY3PLvF2rGjn6UcnAc5ALuVUCxkKC94OG8qcKxO
XG9Wd1Ox6CwjgOFc9q457xPiRuPVUggiFJ3mS48tRd5cWUQJdAxuhJvdcj0Eqxoa
jHVtrp7kJEOb6M7fEyiaYwnrutZknSC1C9SQBdpHqfloHW8tUwvCt0AHGdYdS6Wh
Pq6uOcJG+945daDm0pvRFr1wmyRg4SbhcCJfDoYl8pPBs5K5YX4myheEQdU1IbgT
QZyPGheMMiE37XYD1OykfJsH2SoNsP2JY6gOQHm3BcpsldXiuyglLqxqfPVGefZn
2vCHc+e/5h80IkG08qN5V1E3r8ULbX2ZuOhDEaLWneV/3YohFo1ujHVoMhGjiCYb
6UmNSPExMkRvRvPXQOT6/aCVO29Df6BpLkr/Kd19M3QNOnMUyNZIjH0HzeMSE4MA
zwEXJWK9szuVDn4ZTT8RumY/jblU69ne03fEcMqzEQJ2AH4ahLCPmF87hJ4Jc6eu
V5bPrLiVDsC18Jm07+GIcWJzRWQTbdmQAqjJNdEBLa7U8FMayjQETBtzNRL6Smv8
EhwWbQ0pObT5BkduiYzUaWT9Cr4uMSCqH2fswvX6Th7FjZ9MkUupdW9Cumkq/Y3L
SJoPqcFQIiy+77Eq6yPM7vJQdbDni+0z47Qs3Ds01BB7tyV823O4jKIobhUvpV40
rgUVJQKLYa7xfyBCrDO900tDnIpSWOvWOkEYA/NVDJ4XL03upG5zAoLgPjSkj9cv
irek8jgkStN4jy5RPcaxgDS58xFXGDKOBuArfvL3vHmM6i4qKWZkv0Rr8EYiO6Qi
565dtgX95QtufOjwseg0L3Z5WLDmYAMp3mob/0ClpYy40lvbAmKUfFWyKW/Fdmzl
L5GjGuJlihX79DaS0IzqnWDdSK5OZVdGbYVTlk8togXh2ST8JBRRmFdUfEImFYSN
DAdar8rTvD0rjKGlTu5GEWnFfv5VnPqvkiNajJWgGUNehE+N2/geunHRENZLqCSn
KTasSY7XPY8Y/m4TzVryt8gqAaT2KGbosGK3GrSuyCa7MTa0b6FUJL+lQwyGSEcp
de86F4F8vgpArV0mR4E6FoYov3PgJo4h5tzsCBKyMpFbP7MolPDAgLVa1qPuAa9U
jKEm3EaQnR4KGmDj7NSG/brdZE4Z+MG6SIKNPM0qNpoj0v4k6Qx+onXkzQRUfoX9
bE/IFQdrmx5Mb6uM/Qj0oy+theaAiy5Sq7TN8+MXRis8tR/+v5J4T85O6Jz+dT+2
QhtY/8w/OwNfpvLKo6fXLnpPnxayzzsIOm6n20aZOWz6u6/RG6Q2ukrmEHbL+hBX
M/ajaWb7t5B5jKzEKg6IxawRN07CVJq7QyK+avnFPVktgjSw/CnbZJ8iwzdm82RI
67qvRt3kl1cWCzcaCz65dF4eqbSDtmePwWZFc2Z4XnjiMS4ivTZhmFzI7LkW8FtK
+FMrc3oa+I43xlE6CEyzR6HRKdLro+NThOqee2pmP+LV71PT30RzAqEr30GHzUV9
Bs3VFgK2pIp0/8Cu85FGYM4u26MRmd4JehVfwN2l9uSzXmo4uE5JDwle21FdVnCP
d9Of5XwNVg6pScKQY5fY/cbiJpL9xGyKMrVxP60BlMmb4WPdT8oVU90FomuxZ3S9
upqJfClevXYW731Ym4yoCU6BTle5RBz/s25xiMno/qlZxw5hE/j3q3gz/6RGZv57
yqmX0VGNs3P3QPhbt6HW+EsEr1f8FEEYRVtrAZBYa+DBM7clwbtVdYhyXNGWWMU8
+eTJQLWOcSTiIUvRm7mEDWL/3OxMS6N2nXfb+JMEiI4QRsdnmYaw7eOk7o/e0POZ
zap0qCYrBoRbfVw6CX2pF/Lb3xvqJ9+S/7/CA8I8IU1kAcd7POZCYa5FV+n/CzS0
5beHittt9GHRRxhvzGT2sGYXcRFeEYyeeT6Mu58hdLmvrV159n7QOV4fl7j6nt9z
8L7rl30OfVwhTzMFGdBidxXTiLkrFC8kxUzacjXfi6Ltoc6ksQ1uCciZcmxCnS0Y
589DtNRNJPkPjsJyNdGV2zvt3X7z+0NRuu9UiY+ZfvpYJOlVvwvmFxlxPLZz2Loy
akVfCokwbsYKg/uoAz/VltymYx9gFS39RvH0WtzoWI9Peell15EpEjOfzn1YkHEa
ksq7ewoBSBlaUQ3OHroS+XByzyURtEeuo80T6cx8xP1YFSETz72kwV11YMCPiWgJ
k7XSRybLL3F0wQZ22QjQefmaSMYssDGNy1p/9d8wqwGhwyDROMxjAPw9ag3uqk9v
HyhTgeqfbLybJJSHMJ3uM4XxiexCjEfC0biyqpzBZyf6wxEKqRX0wKlz13xgLYAc
xjHkW3eYvtV7k1Y+AGFa4Wlf/GlXlZdTY5iOLEgjRqIHOzl5Naa+PthBOvQ9Ve8x
ANAKjNQ4RknY7Q7A/ppoNBYeOR7mIZGBODcL/YbJeHY/WAYfjuKsrbGUaI32w2fx
JOeZE1+XgvO43gdtU2fO6Cs3zT2GvGzr8mWt3II8cpiX/XN16Tx60N9fulwe1Zv/
zCNgapgu8mId5jKqaxe9zqsmRBQHT5h78rAFrtMGCPh8R+rkXeOvTZFcrQyhlhGh
YrhxGjRwbJqh0cTcMXnqGFBL/TXRyhyXOmMvja0mYbnERPQScVuz7vPid3B+v9jV
nrkyXFvlIGZnc0GBcN/g/fDvc0LVBwUopi/5eoRUngrGTjIj/WPWMFaEd8qgl0tr
A+4evhrKHk6EzFiepgN8XxTXxXt8gdiP8fnAnQH2TphCYkw+aU1RaXLds5ua1l2H
Zg/4spc2RY03XIPY7LSTRL7DebY5QoLuTQAACDey9J43bjMwvcOon+4yeKjuWt0r
lTZoPYoqP9z9Q+lN13kwV7G3Uj3nMaB9qlkblqr/9fMhaRPwZM08jWcuq5rXkxP9
XzMe+3+R1SMDYu/g8ELiyHMSczw/1qY6tOxz3ucLxlrAzcmEVQLk1IcVY3aSN3Fd
LYRPqRJ7IwJjPT7hmbR/Dt2V3NnRHQjfKTy9Hlo2ASzT1HDwK09LqrCyNeBSlW0p
tpg/RXG9mKoh/JlkD/6Gpse7ng0MEP7J0cfn/rbZVRASTkKqyfZ//QcZWaxSlFvP
LcQflIwVUZDNk6/kiqS0fqxIq/+vtcHRjXShWmtRdxkLchJUXxBkYAZKsC2dK5wd
syjY/F34qcwem9rv6+tJx2lYXFQDBh/a1D6MqSk5r6TzmphXpwdmCV4Ebesku9nn
GmEohilwjZD8iyAnwsWdxRPJpKHX/oxgSUFuOor8lBFfvm86rHYtfobQEepE3+OF
M6owDQswRJDjWh+Ibfl/YTBkVr0Pt+PJqMDc7Pr+7X2nd5mLNoC9eCs1W0re1j4k
LVzWjF0PU5ehuhSzltkHAfv9M8j+9GDevbg/CuoArkZXzISVDzJTiWsPdgynSqWl
57f37BUsLnDXZ+7q5+w4ojJ5dXDxYyyz2UmuvGp1jpAQlJb1yZrJ69MxWb9OwTR9
Y1LwSVUdNpX+aAvD/Vbd6TbeFcqVReM+6mar1xxFFCBK6yEUqAfG0qUZ6c3v91kO
e8CgCvAaoeRSDZPe+UseCjbX92OI7Bcve3N0URP8JcLokxvnckqhkstO3I1Tc1Fn
LaRKMiWWzvPaklBqP7qy4rT33RrPmzJoHNmsDosDujnmRIkqeRl8F8PBCmMANxDW
hQLN+CF8InsV6JKMd9XMAhCwkErjU5IyQl6yPGl1PhmUPUq+VpGQpFPEDDsEFQVM
JcVnOjADeykyiwZu5qJTv8Ct/L+RQIUss5S4cKcqnRu19yi3xIsQb+zGa4c0zTao
sndcQYf21d6tcR1HnRPGeHSRYHEmUF1+YFeVjEaSsJC+AYG9ZfxpPml/96VVqXdn
NWYQpa6fZm3IfK0js3UAf9c7hBzoUKiQZTs+yq0iUr+xg0ZtZSFsvd2KK8XSHHmc
Y0i7K/DWlGwg0iCprEhp63MJnvG4FJDymHtuAOlGWvpaZ/MhmB3U5tDHdohFBFV9
lCWvqcZMt6cpdoDeuN6WOtVaolxYTF3KS2h2D2Jf168Shj2VWNCe8hfefzM2eRes
u3NRhLqa0YpHMgjrmFrGso1PjBiRztz/AV+/lAFmbJr58dx8LS4oo5HFXySnXaXY
ocAvp6oE8bZbHt9zMllGLpLZ+IAK4MCszBmjtDp/xUV85He0W1NLJ9+dPY+cDBHB
9c+VYSpddtoXRZYnleEmyi2KTbF1TZTDOwyaMbJ+txus/cPF0XfyXyM9QiUKMTTb
2tLNzOjjZveMhONb2guo7ZJXj0XqI6tOoYVrrEs9QOM/9XMtdsAqlpqPQ7xv6IvK
jPZr/T/p2GiTbBtNcxA2aJ6RZAIJ7lH4vYFZsjp3/m30KaczU7Wk0IPozm/T++DX
/Em1b2TdzoqvwpHmvj4r7KaiZW2Zjg4L9vTmscWWPuLTehiXswLqibDUwahgs4co
7Tv6BlFl5vHecXXSgMO0EOwyJ5Lb/VHw2oX4EdRZePZ0Fb19IU5e1im7Beb++fou
4oO5y2iKKZtjELlfHsQ/j3WzA9cCtB1jSR4kGemiH3UXWEwB13PW6swzVBbLbzfT
+H8Z/z6RGIEDvtKwF4WDecQRE0rhkXgr01km7esf1OIXkZAhzBAVICu5cckZcwmc
Eo4kp41FryU2CPuddji0x+LELc5EEjJzHqPMzsRTVEAWx3Ess3BSjjOAEjCcGHQI
gdIMNEgbCYMDLc+cQS1177c4pAN4uS67s42/HWY/EhC/1ep0DEuV4dsNlL88kOC8
g2s5hY5F8vRa72ZA4X/smXW6BSaEJYfXoXdv56adDUhCI8MGiqqaihN1VsWRIDMO
IhYBlO90DSm6UzCd/Dt9PxisRDhbDzNU+YgvPdSnaasqHtCBtsHO0ZO5/z1/rLip
QZqUXNZ4sk6ra9kBriZqh77dtEGDI/h5FuFWgfOtzAZYfVSdbZpsaCrQs4FiL37J
RTszPVWCkFwFH4VXGsssDr5srtiaIOqo16wjuseGsDR0Sp2qd+hesmE4Q4/FdZv8
TGrIqZJBdBjjdRvSTNNLJFu6HO1pyl6xt2FBu9sZXkS3WRXr7+lu0LAZ6RmRr7Dg
2Q+qff4UreIo20w8bgCUComobBtRgu2Jz2z2UmTsliv91lebQjq3jScXgNne0uf8
h1fZcGJTkqJXjx3zK+jBhVGjmcAqFVOU+nNBYIJ3fPBSn3CB3/Nkzob0NNDrX9uI
dODnUzJNHH7iWcoWcf41fImZ3Hy5AKayp0fpYpUPW4deHfFAqy/mIir+ivdo8dMk
houXYciDQ0gQ9uSVU5AON5W9/9OF6ewT2holcc2XSW2F2lRT0bz1GnIkzaH/ZdVq
tSNct7LJvvakrqcaTqS0KnjScEEpnFbJ6+mgmcTvc/nSXnmT9PXCkSLcKNcB2Qht
blIS4CzpSsjC7oBh3mpEdmBpQmJxAp4zfC48STnJupupLr4R+DfGdWdYqOUiaZno
kWsvDOo3Aps/qnit4ERGhQcLKRlh3u8gzAnmqEZdmuwEz5D2r1Gt2TlJZ7UBUpZX
f1RwRBuKCcpQ98Rr2+hzmmY2pRrI+Cl7JApHFYho4Pmv3NJAW97TDnmgbOZsd02g
4vFwjDplqD13gV3evWoaW5Sd0ixsn87wzFQyPtUIIAXqjtDZfiQQC1cM3ie1VWlv
ufkOPYw6KubNioM5WNJc8jen8YoyMDzhOnz9uc6ygJfEy+3EWlRVpu2Olf4h7Qsv
yY5uGqK8ShYqtjtyS6JP30OuXMSmPleL7xRC7jpBebLPMXapQB9tkxNm5OxE+fzN
SSOa6AgEKRMB/Lx+Tv8BBiC9VUqMAQeoLpJN4s99lxsU3NML2ua4ME+r5uXOwbaB
eDjDpOgltF5RaIkzpNngsFjugz4YKt+aWclbOig8roRu2HaUJkYxKLMfYT1biXCC
8wYD8ACEZNAqv1ggqCb2wC//Qvgl8vF/G0iCTaaG/ofVCDLkhRl+QHanIiKQUFmr
JpyxiFV7o9vxSnE6/+h/9w3mYojfKyVB07HLqQEqwbhDxDT5n1tyak+5e7nMYAuJ
DS60IGwvxtRDPtC5nxXQsnIN5uBTmP63/sjsQ56vUBsOU4gRWystq58T5XIyctOA
YEnAj9QbaJW2NzE3TAhTykXLofwv+qqGGK356AOPZy5oXy2azFLWCDkSa2AgWg/b
RxjrtKUKtALiVrJWcM56v9Kd7hwH65I8w4sSdWN2NP0OUX/Ks5wOi4DnJsqnqDDQ
KvRXXN1eza8CBDHvhGnbgsm5HGPUZvfimSaavsUXDJmNXLd2ci4O1GTVZzA9UXvS
HWcZZYiZJprYB+/ELb8qaTsCqfPu00ABjJxvah/+S09cc0HlSg73YiQv7NEgKFAK
xvHDVM5SMyb5DUwIHvdC3xzEbrcPbtoQ2cj/a8GSw8eBC+Q0i410wRek2wezj/42
/8wtBUlDx5+33gSZ7Y4c0cVhcyNRgDGuJMetfKBjo6BScQOn2D92PoXeXQO5ZCm5
2o0ZkdXTejtyfgczZE6ckGgl2JyoExNC0KX6dbvg7HPJIRQBkLgPw5MKRU5Rsj6f
Ae0GlZZvZRMtZl3oU2uDwFPrYf59EqQXV52cniTaCw3HpHNGN1ZEM2AodDElqXO6
OFivT/cHWrwYdzyhlNu75tm/VqxJpigjUrWgZnuqNETXmhqy62yQcwz8AO6s1gdj
Ajpa5BslxuCHwhyFCrCTn4MnRccujTQ0CDDVbU6vxujpi1hgf1GA/lzoTcU/lJb2
7F+qc1dOK+xZhygRqF5buTe+XHnU9iXUiG0kRQwA1gduD8s6TCV6MWP9mCDq6+VN
Ayyp9bajMji5qh0AAUtdaET2daaaPlsZ26TcGu2B900P5/Ajw86Jf67vjHX5ZTh4
aTMtSgCOo8ZBz5jWVTUYgcq6Iq+l8QePfquwJvm2EYyP2zxnEfmjxmXdczG/oW0X
Dr5GbjwyleMhUg5bgw/ugWv8NpMSSUtKYbqAPtW5nhF2Qlnscuhs8GyLzR2jE7gj
y/r2Hp6BpaKNovNlLqx/DNW8uttj2IplT1D/v1I2fjWEEe4ZOrdUy+J/pzbKs06n
GEVaTcoC2kJOK6S6N/uGmn/aFhlRVB1c8WdHvHQuLJepB2mfmnlzSQ90XeliAkF5
Mlp1D4IV8ilfvPvh5dOfrGOFgryppaopJanKq2b+qZk3O8TqMTJmHQmAWJVtXcaD
GL3+9rDSOwSeCh9xA+TwL4RSTjHp4T97Ik0F0CT8BXxUq/UcJ64VnxHSvTwE8jac
oqVYKBeDli36DJv7PJF8KULaJ/WqFkXOL0SHLaUtMuZ19Svphrh2HdN/5WMGNZzQ
Z2p5Ib15nNWbGY5JINskqlfmnylfwpgauPpTQ6UgHeblja5Yxt2dtaKmb+lSZSSD
/F7yeHTVVuuXEu718XjQZI2qU7oZuJjn4bKtSIGH+DSAoP2wrQmoXoGfZEiyvzAm
lHfztz3C7Mqsen2FUvzSV9wcFFLcqEBc6yrtKDJU9RaqlMS6Mi585EFYeiCecQ2I
PHMuum43ZFNHTotFFexJsbnRJn+JHLRRDB0bMfPX3xreoNf1OVN9RhNoADZ9IHyf
Rbz0v1MB7lzZDadkbdgNN2yqahAEGomM4iyqUaJlJecm4WdJbRDqkUdnz+fgtoeG
ZT5MnEUEnmSm6nXmw74jq41w8yDHlKthsOaVDgcxwprGCQJzES33nwmc6zFkayne
cdI1NsWni3004keg+VpljsDDRWP5aIryx2owVTdVFBgIl+D0Q8/8o3gBvC1FzQN6
BE12LN3npMV/xcMoNw4ukXMmBkEPaiyew3153bnF+M1z8Att7ywocUDhCLIU9nzT
zx1YAmSnD3HdLTeHY7XeIT5ru8ltAe7LODskfK/lgB0zAww7ZQyvpwLHrk25Z5m6
XEG2624O1m91yVGX3ekAWDkY/gCXeXTova70+bZzl7EpBXpAXFKYeDUTMmYjJycF
48Pydpc2uN8d7nJvvZ809yrFnAkpo8z3T5ceoAf6R/S30sI+sV3QuxVIv0JzEiAt
/r+FVkzRZ4prqi1rsQedIqBplserWEVnAN17DPWIQuIRcYflHwvKr4KQROXfj6hK
cr/uE7zFU86A/VKfN4m08RX1/vfikko2cShmSaA9gSV9PBC7Jveo3oq055d0gW4x
sKQUD0Sirt8ZesJyCTXo42SNrFanGy382q8Uo5Llxl/QMArjqDfy1fwlViVQNJWE
VyYu/1iSfnXJ4TEIeipHDyMjk09FfWx1aUmnfCDyUnSaobJC4v0/l4L9B6UBsKeJ
8Hx0qSn3QjmRTgX93AsCQjAN81iUuEe8P6kIjWgPbMBoKo8DCKdlpNbzSNbXws7D
64Ksdy+6QlpWnoGfnVYqqgDhjMZFAjYEBdTRIrsYKKU24Wq16o+S1XRllyvXRerK
ywTzbzsoAJsRbfexEMv2uB+N/2+ncvt4RdmTrWcyA9GcDoSk/2zNTgiWTjgwv2z3
1xCB+Gh+vza7s+tJzfYABDwu9iRJkWV9J9T3cGuxAZNXNmftGpHSXIPNSN6qC+si
4Xb4ooHVSM6xEgkhbOOkPejGr6YROY0t5V0VFvyFspKWljXUqURzDfvxRBcKh6sQ
c9q48TACO8Y3ImS/tRxj67LrNYlWETBbr9I6jkvvDpGo+55U6zGH/nZdLzoKHx1/
1VcLch1MI9xjijpPxPyFv2qGdcS23fbxgzsDEgwJgTB3dj7gqxsvMvafHvNrI0FB
qPxPUXnOVWzdzXlaejdnc3WFNxM6zX2nOVTj6DkVt6aC2ssXY4WGu9rkQvPOoe/T
YJ+uYkIcuQYNP5SZXxwkckLVEjvM/kai/vCp/JFubpUB72I2KmwfTeoESXzugrNx
SefQUkxfre/HzYoL78n6v37CpiOgXqgP4nzjhUnggcqSJWOCcqWAh11LTKLrf3Aj
oKyjCEvWS/e3pTX5YrvtTlxlmJpOiDYh5lVlwPneSso7+UMxvCfzLrGK7ZfQCOSt
ckIQoR8FHl2/R0hdgcNm0ke+4bY1oN11SuvoAsjMjVwAiqaA5eDbc9bfnb6vHT4U
zaACOq7ugpc8Dy30OmmwqJDO9TzX0E5nEYtt1zzaJ77QewwzMxF/c8RpnR83q+5p
7/NMCsGZdjYdN4wNuKH6vqwSqzF3hsnRc34HdNKqyJLmje+p4gyIRdGvvjXewoWq
I8EIGKgELHiEg17YhXxp0N9lMuQUQZQjIww1NVXIXaFkXXPIICPEqoO0piKYBMFS
6n8NnoYOmO5jhma3fPNDVmooR4lYcJMO7AnJrlx4WdOS9VTRa0jsp4KQ+VlAV2aj
D4aF3Y66P2v0ZYP21KlUyDV+xRuS54UQ4QKlg8cS8dOTDuNcOh0BgnRkUG29n9ZV
QRzGS7jGJ1jp1Z4WXJmONpLQKbAKTvQHaPV15K2V/Ryu5f5Hnu53yfJWU9AGqhjM
CXEQZufQN3WhvWsPOx8kAHJALY1VW+UBiEKhRBVOTUVBFgKD8pq4aoMvVl4mhpyR
rwexmF0IKS47rybv1FHXdw33M5qcuggmesAMlLXW1WJO9ZjreUiB4jEiEPxJQOXd
ZWqYEGDtQbPPUfplljcUkXa8Tp1fWp+KrIrpMDZiZiCfgdtICjuYtnthYSpVXf8R
cZVbydeMINv5+Iti+hf8jUt77q/+bImRxJYo3dIgon3rmCF3oRPl+YRTu2qvWuio
hPX0rUgQJ1hRJ8Cn4Rhfdrf7TQBb6JJhCqEH6JLY1QeSGPhoL0TQgmPhRar3Dm8W
f7emBxqOMAttyZ3K82tzHlpDALG2/Yveoc1EO8aw6k2WXHnRIKkDP9bBbH1KGZX+
TGbLvxIYVGHnEJ3cvRs5oIbDz3aaeDt7gVOABbmZjfbQWKoeZW0fbuKWBMEEmekJ
8SarUIe3qf3wZRgUjd8C96Iergr/hhf30CBKED0/enygc2fVPiBbAAd7B9zYvjX4
usOnhAXUAchyIPBfTKKOoTrlcJlZlLVa5rZHpZmKITvgfT7j85HZYS+zvM13YBr1
QQA6YNEWkgHmyd7aQ3hrcGV1l5ufHUuAwtWfv8eI0zZr1rcArM2E95I4HQGhzlBh
qUDMp9+j3+RrmVcM5NWCPp/LUO/5Nsim1jdDCMlH+I9QC7e8iFeCw9RqCkRqBN3k
tBic5whnCRvtFuZtRQZDm5Ao/7lbUSXit20w0fOwx/7NS2KCvb/S55X1jR5uuQxX
+3924zxc7sdXu69JHhf2cZqh8vluTMvmNaLqoglMAI7KBNLpPMJ0AcmWQHDTlj4B
rYBvnMtrYqOB+46QQ/NjXziVCg7yYcvzfkd9oXlAf5iigTr1DaNt9em2TUsl61ZZ
id/zijPW216xw9lrE5U96qoSVktZwWUgkqEIn8cQxcJvPopxPZl23uZoeGPbn/qg
4SAofhsotJfpOuK0kW68NYK7szLhqAc3vSEGnXi+o5CkXX1zFcJ4NhIsj6dIA8YW
XBUzrozvnX2Gw9lRW3WQWFh4Z9l3BVRnpXm9zywEWLV2E+JX4voxB6g9iy9vc9rr
z9gi/0WMVKRlA1RzgivlsN47ZdEz70OdOjwlK/oPAW32ypD2wLeVwjpD1Zikv/hG
GHVts3DmsercvzkSio5lCTYzPv2i6OHVLjb82aq6ZmqE2cAinsTjxqYvjBHd4SEt
2nq7ZZmY3vScaDHcgZkVgNKCXjoCPGow5GANKnviWcvL/3xUalf0iKI/8ll0Xxmw
j66nppZ8HAqNcdedCHR2oKFYDwy3bu5oM8XEcuuhJr2+3xR/7tLOV6u8SKB7dqNg
/Nii3myt0nrhZRT74FQnm/oSZfHy1z299iWrHJ1cFMWLO4d7CgF3frp12JLZT0/B
QYXaBlrl7eGMyOf9q5VU6AOtmWOvzNdN9LqJEwtndk7gJVA4OmTdnVjdOV4BO6QF
T7S74svskD6kHq2CMpH3FDlyE4fv6e/vemBdZRLw3/1A2xh4YFYSASopSNxTKP+L
h4sSO/udRVHzt3YvDwUJ0d0ns+9UH2vV6SY3ANApw62PLOE8RGW8mYKu0QBQi3Lx
zDFI5JIb0TLRnQKN9Jbx6200Y+Z4ElIaWwu/ojCG+LXJmeDjubDY+0rJUgCctWtS
p6hXQszEV3N5Ce2oiPKBNI1IFmESEHr5+WGQ3ll+b6ub/o71o5HcYV8tEu23FXZa
HrLdr+WcvT8u+UiKe1X6ChpZ3DuWZRtp+Cjvq+CR9JhOidZEDTzRuCDP/5ZpJa9o
qXaC2h5u3GzbF63L6XUHDXqJ7n/4MCt9PJimNeWIzB5Y+T1iZLaamWMcI3bDQuFE
BXs3Pm+SwitY159MwEJqG9JfmeASaBXu6N+9MEDbDRvyqthSp6mJZTXj0aGqtp0P
/gwRV6PmsAUcZY8H7wHOkpwN7zxTgeyDlUEQ4by458KwjRtKjn5S8cLLxGL48FUl
dviWVB3Z8gOEJYKFJaXNaZWZ2FuxjSyCOkGxKmsYIqKAgLZivzQOq980I28HjG1D
WqGcPzUdO824zgd3HZOj2WmZDdqL4B6Dl0MXkMFpXqesuUbZ2ysTk5e1RKspAeQh
EuZ88ncec4jKLI93atS2pgaswq+f88BAHxyonMNI8ubL8TCGIEVzOTpgQtVhTePA
q8QBksP0FAy0fgeVAIXupDNnBKATSIYS/HSgLhL2j8GlA6s+iVae+0O0zzaBt7oA
4djbD3PWeFkL1ODcV1O3cxZjgHA4bOFtp+6Y97ZhXkSL+ZnRDRzhtmM/X2X+AfeF
OBu8uhwL3BJcHH/iS/Y92lLTfYSGOCgaB3iJexn2SybcoNCUSPQdB/VP0E+v/Etk
c4mDar4RajwvWkLoNBJB79N250QnYcVwAIdYXhIar1FWbcmhkzfwhfujaW/L5PbL
qDf6j/Yh5EdDL39rs0HUoJNocSXGK/8PdNo0Dd1ADcmOJNYpuR1SHyJOw+BeDmac
JxHuzGjZXbro5vGhE6JM7IEwocmM2w3E8GnGVOI3KNCUVRRooSC/1q4urZd+xOMr
vUS3OuuTBJxFK9d8cDoAWFikLLZX73YqWu1H9v0zmZW4TOSUTY3nl5NAGWc6xLPh
I1Hd78U1a7WYwi3nGzM/hcgINA6NjJpGO5ClSLGkPAYE+X/GQ2hP5oArPXFUCrin
6gxDwgUrv5ptjRB65YpDvnLm990Om3+02RCe08KfVs3/4a4JZbik2WaDFnSJvXLg
JEIItzNH9+9ldDDZRj82ZDgc2XddpaTYGEVxz/6qcjlLsl7eMiUdFnLlOeY7MICm
fj1a3GTZB+RaQ7ejRhCfzG7L3KcDXVRDDFLgOFeKgKpP0paeABKugjHeyU3nkqQD
JC+eKC1STSxAWa5TuErqvRyrzOR41G+u76dvqDtsbpm4njAAA/fUn7j6P9yRBKUE
UYmSrTT087y/c6XYKR+06Q6u2zPqIMxEX6SowW/MTk0FmXLNGA9csBmAsIomj2Wy
ir34xsvqLDV/7UgGpkfXBoigGWMthTFArS5wJ1jg9qRrfQbKY0tJFYfci9jPhf6Y
OZyS1kFEAZJB70k5Ewkboy96vwGc99XV7YpbtuwPR5/mpmgwnptChcPAPbbH/X68
+reHPOMaTeva4a2rQKcfUrbC64HDbGUiBD3XA6s0cGPA4geE9cWRSKyy0v8fPafj
MozIcq6r2oKXd05hPZp440IbMyyYp5qNHIrb/9Ty+mNrSaxiox/KAQVW5NVl9Ln1
zDMRsb3LMojVl2JTc+ABjNOY3bYCSQbI35jI4+1S4zU7v/uM8uKKlJV+uXKbotXI
592k5lboZCJHVtoTJC319VKGlaaBBw4i0Uvmfxlvh/b2npNapVrowAOjt/1h2NfU
6mWroyihfkEfTR80EE7OsT5Jedj/q/325Si2RKdlxtfmLyK5lTo1+vTJmxsN79wP
eiDYlg1Wt9EyV1NIeQ3SycmQ5jsG0OTCx+wLlHudOPFZGVj1WBKeO6fDyM/XzBdF
T5a5Zxj1COIumay0mCb2ogl2RNkRhrTjRstsCguxw3pXUkmGHMpgh1DQ5eyGPar5
EUVy3NvxvP00PwJrZ42EOda115hWA5NG4wuR3bmChR+U/Ua0WLCGfnoNJyeQDLw0
TTod0hkG5J/g5VtdSJ6jp3t8fxlLEBY5gy1eqedZZgxQYZLcrnyGWxd6GLuaqC/F
iVn+0pwa/uXweBbNK/XBEF139TEUDFuih493p5pW5/2gNmYgaXUnyra+4hKOn6Qd
uxTRJaXFKE3hKBfdXWCtBuY3Im3+ud8O7Vuql7WId8DSMs3IWHMGoRJSSyUS3S/H
Zc/1v0/uOwoL6xTZ/vcSGUkwkFlIhLkcLi0CzsrnZAB0CnBSO4Uo5M1XQBqW8N26
R7QcRbPhcRngFpeBzako0Dgu0NMsn8IGuYPLa5wEmWkRjA/BSWX9PUiqnoqNXGI6
Dyk2L9R6mnO7NT2VchwnO3sq5AAfUsto+7xHQ3olFYjP7Px45mys2jfiM0JEMYAc
U3H0TXWKQtvybgW3ByRHIVw+0Df+Lqr3vGQW5hbqTPTF3fWA3jQQblWtazdF7wdL
0IqjzWZfUru+W4YjKMGJP9uO2ImtgbFa8ND0jfU4X70aSD4/1h+pR01zwyqAq+2I
xjAToc9LhsepGcge20p9/fp0AXE99LWadY8ZnoAxKX2RJLYkHttqeErR7kSxbhJp
gQ/9cBIx3dReU7xgdGI0QY8YbaMdib/lzihvP0JPBS5reHp7CPIYDliiHGd1/iu0
zr22WzQs01Et13r4tKODYvrkadxZh6TQWWU0dXBJhwalBkOV+NpKJYgRxzXrxn6Q
QF1nXIuwy0tYxcrCwRADXC9pZHA5PwgARPYTNSh1dW4cvch12CIijxbkrUA3uRTy
H6uzx+QuAlRmjhvyHKKfBcZBrCZHHYi1IxyYiY3nT1bsjn3ktg9es5HQj63dQseL
e5gtSnC621KWj1+sW6MNYCnijv1fouV3Z1NofnO7tmVsidFAUJfh0mNMPOsoyBKt
k5BUSwpByp+pbF2cM7V/aVW3+ymv5aIsHWNEJhChgaehOaAW1ArdoyAT4jONcm9N
gbsKq256NsT3HLevGsv0+vPVn7k9Gg4S383VTz94HMyNkYAqelkt09B5DLfp7oip
uLHuoqaGMXOb6vju/ZEvlcSw/WCuPcgtut7PF+CLZXxi7ByL3OPmAZVcVeBA6Moi
B6kbBsCx/MDLIzN8M2Xhyd7NH/AlnPinZBDVBlvadxl97aK9t1pJBsf+qv/+zXZN
PwjLLGCRkFhVL55Cl58wgejvjdIlgvR9ETBaAQ1ejuEhR0Gs2RD+yA5wFm+28LTM
L5xI/bDmR5imh5uJdRZrIIveAMDssYmVCbzEoCfFz17F8HOOM/+C+HdTFCggDEKP
JZ2/bGsuzLPbcS+OTRMUVH45ofAeUGh0bRaotWXzyd4lQ/aQi+I6UlYkD/VQDPSs
6LFFJmcBZ8YzEwgKRbMveNQLCL/mdkJgovfqYX4QgP5HFkZEJM4WXoimBpfZHNHb
fjFktw6XS2EtFSxVK69eXHlnyW/xBIEg8KixL7oquFNXNXBB+40EFfi9EkqpIqew
gIu7AHqdYhUCk+uU/otx85kP6QhK+iRjUdJ+teI4a3QZi1dk4+U8s4fA8MQwuNzN
B2kiZkg5QeTEUrIZszNPzGtDhZeSYDZ1UXUS9NZ5/IWFO3w58tXtEBP5OgRStr4Z
/C89AcHglBudEECJp+7DCgGo6vruhGwhEj6t193P/mUCUCBZ9RR2QonFM6974J85
OQ//FumqyLHmtIg1QNXYWu/KtlEumBDEILWjOIrQ0kseqO4vqGdd7X2+0158RWoH
sda0yU8NzGQqrX0LT1di25lzvgkw6EJiibFHkDJyQMA19dQ+xJ9acpf2Xfp+eWKS
yXwcp4ubMDqSBvIj1/rYEDkkz+veE6yGJCq2VDoBnmGG5J4bKFsalsdsubp+Tl2A
tXgu/R54zA0TGaQ/D4ZfIB59aNJVpVvxTQjkSTHxpe4Lcz6ULFwxwSduR8KFMWAZ
IXwZrGgTNyjMhrAjGcNQOL7o3wFf44K0zkRkZtkBn8YZi/6MOyHjYM9IgW55+RR7
IiwxCKtzeyp70RuzvBdYtFgFBRssb1pnt5417cFj7K1weteBweQCVvZZtG/jZm0d
M0fx5HBPSgqgjLapBr8qBSxgloxtjkDOFgpFsYLH7jL+Ah2TeJXO9vb54lAWf+Fe
f9K7sRBRuL504KKFiPYSFbwqpWDNSSv1/Fym56yC2Vc1ipjEiMYy7UXIyFkOAHyq
Sy+82lSp4ek+4ctNE2FtnXo2Ktjp60PhUOxBrRB5qi+XRP4c+sxIhTiA7vgoVFq4
96R4zBrmn0bIUucCqm/fjXojAGL0LTVL8Cjj9QB3Ksy4AX+TitBmV23dEhQ6Tjzz
Vs2C2InvJS4ycCcBqvYMndH5bn2nciSHJDEjGYtn7r45plw5V+ElQqaXPzT/odEV
AdWh+iM07/lx33Ao4HXo7hI06DKSejZoa9nf6VXfZ/pWjsqgVbolmlPkULRe1AZw
Q4RQoU8xPZHI4PZig6I4DfwIakJaDRWFP1sUUG45L3ALYLg3XThv2Vu9U5zX8Bz+
UE5m62uWqZRbc+cY+vMKC6PXUUvcdHBUuh7WLPsyGNgLkil8xrgbXhhUdWJuEli5
SROSKjLNSyqhSlSb7YZ9hmWKJb1YPO7L6u6wrkgJyIg9i7j0XJc7ZVBWSAsePcSt
n7Sf2yXyuB3pKUtd9inQ5UR3fGHw8TiZDoSCLpajyd1eDlJlZ0RzL1L+L4CTEVAq
k0Zs+Ja0RNZx08by6Fw6uz/unF5/V2dGUa5M3/wbdbl6RPMSvXTv5/JTbMJYy3kC
mr8KfQMOy1VwLhuHGZahQ/AoEoiWG5psxChzx9etWrx84240G6NV+w35ROVFwz4l
ih8hiRkE5xk/aiV64vfJyPWoOZ1Xyh0elsaB5iujMMlsA7deLF4RUOBMcJ6uVf5z
sKeK5NIj9MqLdIm6bnOWy3SBk7YdmuOtUt/MZDbDHk63mOF62nQA0qTJj6HWNmPq
RBsFA0Qm2b9P3W67DaqmqhRxzxx2/Cv+mE/IEJTP2ThsXOQHfND3WGrca+pPTVhJ
n62uQgZDI0Ns0rRLspgVujeczIALBM8RlEhcSir8y2tnnnuhr1N7D+k4mDJV8Noj
DxGLnNASCfu2nSfF/EJAkNUqdQy3DVf2XCx7zUfqRA2d0VPugqs44UQjfAW6TXYE
vtiYRsonOruEzm2xHnEsAkYzeJ6CmUs8vC03cxgtJ954HHXiW6szWt9UtUyuz9SW
HuB+AxlN2Keuqfc8TPV648OZJMb9l9bCrRAgoDH+jP5zOQDFQ1fHQlrhHrBhTlWv
+PKGOaYIw75e7uykGdroSw69SB9Gt1qR5nnufp+1tV6U4rzETfyKrJ6KPBPLVipz
3rnbIAjxyzJKEufiAB1v7jjTyWtekfzvnJ4rRYxqcxednG7h8069T1QPSAuIBoPR
18Zk4V+i+KAasrKegOIb9U5dyOqMmF2UWmEfVHRz9V0WFk8SiuTab4pLNA7uMxpu
TtEdFGkP/bTIJFwM13+b3YOngOhTNoVYdNhfTLPdTUgHJwS6cVi+3J7MVooW1hvV
soOZhM2h0hqh8kQm4IaeIBqXQ8dWTlHWbCuYwRzLMfmsSmmGUl2bAMggv/Rm7kNm
gLnx8u8MCeRC7DXUZGvaK0g/XWN+L5ASrQlITfID77/j4t0L1epbbEMUbO66sy/q
eeqyoJazi7Vrg5libk2bZzNq1uAng8s73APWPnmz6n+PAJBSBjz8RjNdMdZRr9Ei
9UuV/nS8z2S3ybrVejxyJ5Hyo1weC8KULbsBuoxSGwBOSCErvaJj9JvWjVbLrcXg
pVBh6iJ6xsP+81vza8LmX/ZkgGkTbqFld03IkW5TrE85pMzpDoxintjbMmZlMY92
stWXURzrSK7CLHuqDwdUkp50Ha/uM6nkj4wZcsNmSfOui9Oz8yXyo8Xd4+JgGNNk
S8lv+3YZTuWT+1EYgTSoQ3h2h1ECSoxJZv/MzhH2Qzhz+eGiPiAluUbqJdJ0ZVAq
oV8QM9TMaQ1B9wa/ILgxzQG78jE5oVQPO04JQ2AfzTlbRvkIuCyEK9wFrM3qzgYt
JOaH3WiAN4h15VHNesX7avC4a1a71k2LRqj/uGAsS9apcHWHFKcbt0IWKNcgD0BX
VGORzIcjH3PaXVDO6CGfsHiGobSz6ActUlrjel2m3mgECnJDs1KA3DlieoEn1Vn2
NodTZgSnoFB0rs6qbtRTthjn223jcBNgdCpJurqS9BLjEzWDBu8IW8xixepldvq8
Nwf/KwMmeUPjU6mT/MWnH7tnRLZjfn60bKJa72UYpkksFOPi/ywVmZgGNC+LTz9N
LUxfYlIH98LAjT9PjNhv1kOuo10LOeUliOW4qY35qJvEhKQ6UrIXWGtC1S89JCsp
aneUaLPahOrw+1m83uzQtO25d9A6WMO9+onKXH6CRe3uHa7flThtSGosjJdgiEac
DCX7oB/A32qWU6mWpXJdDqk3R+9q0z/fcPjr+m621Sm5Y2VYuXoed9agW+RL4f2B
kLuODa5YXHMyMB8LnT52rx03oQ/zE0ZCCcDT82uU1mfZYzEjbijZlmhxS6TOe9Ry
zrolxqYcxTRyMmd7SaXT3JSfTxaYXf/h13yDm4KFGRa3fGrlhxsgnv0v+MZv1jwk
95ZvkAezYMx9nJsvfL271fbvQZsZdI41mVBzqDbbZf9M+igPrlAuh4Uhke5DEkVN
55PY/35ckodA1ZRckGD/hQtMzW8qjpd1Qioq6luUQ3iO+qPCv4lUeouFFUKORX7Q
+XlUcb0PdQSbwZkBNCB1d0m5eGKJGig+m298DUqvjwRYIHoLSb/2UyKka+rJePvn
n8tuh9pYMNhEOqvUa35mUDBJh5KgDWlgUDoChE7jT3059AjXDsDqfVbcht2+1eEJ
cad72Bn3n1afz2ZAhc7VtQegoOh99uAtHwIQARqs9ETT8W/ZtC8U4CE6+0sSdo0v
HAeQDOe5VgmIiZMP9lkZKhcU4NyLHqm9iZaqB0Xd184cjPgyCNVy5T4lsq+VJpPr
Kkg9q4gC/ApOfpsWBVDY0T5mzEtBeG76XX0bDtDJ3cP9uQWmSzLmV/K8HbeRmLer
9IFk51M9pBgfGWwCogrJ7cJrRzRGGhUzsbDEA7egg1RYlLtoy4ukPCbDpExaaC3a
TATg3T8gUtNdpy5UOpCFA8pe8bf6RvFxQIB5v1vuAEMBN6Di+wMRVrShZptGwkx0
UFA3o1NtNzvOwngOKGdrh2v0XVthBt7f3XGPpIkPIiJHjKAKikSeZ1mrMLN+NlHW
/cD9KDsi8qynlGEoFYcMYJOqv86HY+BBPEZO5H3V4B6sTrti/+iAERQJOIMkPF9z
TyCs/p4R6ZvZ3h1wlREkKzNXAK5pi2Fj8pdUPx0RzB1YJXfy99vlpR/YK2LaLNYt
01fLxLAjt5hPmnM0nhSx6wvTdrMRZfrrAkrc9YkXmBhyBZ8DW5SSDRkGOls6RjVX
10yIN025pxYCsiHdOumfWFzB+p25wfTE+HN1UmsnOgCsrhdn1WIfREdR2yqQcV4K
PUEMUDYo2WJTdcaJy+JiPUR0dB//LsIZqqFZRWO1t+aj77vN3zNT1mQaWhTWNTIV
cCDqjHyGPhpyVeOParNeecpnYIhqHyfYD+3BZFWkzIN0+7ISpyvdiMz5n5dJVIiQ
lgnMqO3U3ZfjXRcPnSwEXnOv4XdHWzdMfm3ZvIIIGX/PJ2KUE4Jadz7bL+N9HpBc
sXvK3QkOIUPGTpJIEx7E+shAOHAIXD8cky7a6yYlY+oHWRhjKzZvy+REiuv4H4DL
upsU5ImdwkHtBCaJVMKrO9qGPfmo/dn22HSjMw1x8iHOGV7Ey/oAEODDTfbm4Mtp
ulVO0GAfjKqYpV6rdyn64UQ9rxcX2qAi9uVrDlCW9QxUuZGAUYrjxyAm6IWzGiWt
YQx+EXoPlQTctm+AjJMr9yiMwegW7erEK8wp/q3ZwCP8BDbjXG2pdymVrNopsHkx
Dfy26umhn9jibvhm9+Q5RsopCwaZeHJTsj/rlvbrqJUt4b5cJJelFlDrg543Guqp
2MWVkn4VrQgzv5gid8n17wxJnkaPbDVVqFtbm9xlobcPA2XCo4piOVjNhcWc1B3C
8s5QeXqAYz8rBHxGWJLCTmLCsAkRibkFCmJqjWcspa+ZTklyE09KJgZqQ+RDFq4V
gkpk5csXEV36G82aoyx4/C2k+oafGb5ab/keTKZvQFexcs0ea90qpBpcsjCoKk2+
fwhLlcl9kiRtUhmdCNakRmu2zlfeeUz2tmrCLLNrgffTS+BxR9DpfPPRFAoA/UFz
dW9hnKGdiZXNtQMepbZBh9egXa31vyZNbOadfskn0i0uxudy4jC4UKPR4TCiYa1g
Y7yXsd7+Ok8tFkEFbUbHV8kZcvjRMgHPvVJSAahZmQaGb2bJ9ZZky/u+meLhZhSY
fvcsbjf1jkCNy7o3lu4+g9gz+zzldA8t2QwvBcFsJiF90SpXsRzX+LOZd0kcB8f6
PeqecSZpOw/KhEuMJqV1F9Q5L+NuHm5ORMX9sOC0Bs8Xw5x1AtHUnHJHgFm/Oqj3
Voy2NDxSXB8xzoDz0767bdSL7BG+m4/xsYqdaVYJvUV9INYdKVEtY9NFreMsRcVl
y5L9AripBnuvN/C5wfG3bmtsWv7/RbFytbFLZOSjjPmIU+MKD4TLYHwcFh85vTC4
fZn2zvGo3Q6NybGj72HH/8BTBoogY5ZnMg5DRL4Bpx2f75OpKPyaTD3cS9zYBF7v
kVVhD9CJ0wWbOwK4f11ATzgFwYyH/IhzLQF9TPHCeEG0K/o5vm8KU/80/BbYp1SW
34xRoLtBENcvB3luLqrZIh1Dqpx2KZrthA/HVNB61wwDnVPeV0VqSHI0pG5kARj6
CL8wLHgJ82MbgKBEbn3bSOcDqhVYGXhVARbdD+s/eA6rTTscCPjXNZunyF6f8Wwz
eoF7YI8WgBrPuyMioEovnp59Oxezr/siFj+r/Bi/PvgZCUss0lwUtdBEd6ZS6gtu
jAs8MQDaQkgtiWHYTY2Y8CIkgexBvvsKaiT8+7Mg5InP36v8VzkiM5sryCF5skEi
HoQIumWfVf+3C/28fxh6uoRVslO+lwHWAJdi7L9/unpTVH8lYPg2keCrk5gHMFIa
+HZWH2v/Hb0CdJcttNvjCLkISpkn2+PZzdS05+WOmPhbuxG9XqvPtmj2jvDbDTO+
hFNZjqjG9QUsJBusd3LdeI5f4hYU/uApqlfT9q5iQnxzMgKDvT+llft18kaFhESa
SK/T7ujNIo/IRCis2u4FZfSoYeVZXDoLIzGlVVy+rIbmzlKwC4bj16xEhJMzzQO4
OTnV+wXDg2jz9OpCTfb3aIC5gfUmLT676QGP0vWlPXS+qFCNYWsdfKp0bkVl5fmz
yf4GUnyU8iq68XxwS0zC1Z1P+LwRXEfoih7+65maIzUv/Lzeq+OLTWApjvz786GF
vCblMc5W2yyN5yz/V7hIlMsCzCrCirq2GWoclGKso5AlAUANKU/i242fdlL45BZ0
FryBgK35CfScyVZQaM8YZggRx2bzy5Lq6u2cqNNrbTktayntXm0XCk6huwLOvgZN
fC043Fmis11giwq6fL1VDhybv2HffNRZrzTLUyJ4z14zFOFfKCmK3J6PzlU6OQyW
bpJ7c2mV39qkietaK1f6bUR9sOg79G7AOfCO26GRMsImilS+rttQXjeco1SgZeyL
yR1FUS8iF15etonfhuwPt3W9yqXNyLgvr/whhlYWQL2Rmnv1lHcLKvg9CEf7ZEwh
EWXEdHB07unU2XGtRemNTEs5NMTJHLjBxoEL6Xx9PZ3VIzU7j+sglbM21NXt/M4/
Q1Na44zq0keNFPCXlwfsjlyRLBsnw65FTKNBUW4iJc1xhGLGlHcjpim8DmHAJGXD
5+m/CBiPZ0ebqbBq8OGBmKtxo9oQaC41kjx5ntR9wpcT9kfp5EeIQh3na6nsCJLC
ftx8x1bd33RC6LWxIBgk6De0indwIFcA2bvTYUwlGHYLjaN4swzZIcVEiaC8rqMM
y1uvSmV1ST2J7mMlVRctNBNn5GbGgz2Bc8ZEZgrUS1tB37hWa0IQ2eJvn8kSgq6U
rcJs401O3i/zcMjmIfNvP+GM01lJ6boOPUPVk6tEzfoFDs28YPcqi8mjXSJ8cjdS
IPgo+vVmZJrKbFnvAoxgI3CjRCg3sBLQaaWSbiLDnEvgP2HO1rDwJ+VeGvWNqy3y
GtVV9whYloFFaJou+4tmpybnUtXMy3qv2/xgAu2PAuyJCKa3ruBba+2nK3IhWdv5
IHL4X4qL2OWV5v21GqACxYqz8FVBNoT+eIEkw4UOXpLfEV6EBazEueqFkuGjrVf4
idRh/j4WwBydmfXUCOlvY0UIr7XhSPy4OUGVd4fE/8pShFmtXcvUqDfj2yyolb0K
E2Wm6KUj8+HqmNyY76JfNSyG/dED3Xo3+X75jXXDzB2h40zbTyprdFPoIH0XuwPa
XcAdBD59L7DNtRj81WtFhv1TIZa7thYDmnqZtAQEQX/KP1iOEa7q0D4WgmptsNRl
iuTQ+s+OgSMMQP+6KVj+B8PfCxFbARJP1zrc+fQDspBWUYRVAKo3Dkjl0l1NLYzx
7hqK1mJuWXgb40TgGyRwKfF2FCXXusSou2PQJBR891kUp0ovci9Fu8AeO/2H6YsE
vByvFB4cvc99woys7viKtPms6g+RzylRGbM2F7pNjha9YA5lgXa+gp1OXgBx9txY
raF9sX9w5DXXc4Opa4T8oda+ISkM49TT7e0AebhS3RcSZ8Z+hQmTwoyEMCK2QXyY
AUKAn3sNUUzd6PwW81yMHq5khCWMREhp+Uwmb9ir2Gm+r4hBEebApHDkecV+p5gT
aiXML4XFP0Jwr0X9MdxcS+LP/kiESurefEOSPYFJE8NwVJMJ7I7jVgQAkRrCOlcq
8v2fI+oMAASSmx1+XSnbnpzVRbZvYqaSJYJAGqWupKpdM36jWXiUbaIe9jJN5wAX
4xm3+gTOT6qgKU+6HToqC0clvDvZwVbgfNRuD0rVCjAPEs/A66JrRVX86yxbHu/N
PVEJx9dR4eJtqvjFk2Fh+m8jS1+J+sD32Z0uP2PBfOfxknGWX/jliKOtYx2xG7wR
0CTuNJ0GEbTjQzm3N5KrHAhcGwJEdGOO9TLUsBFT8p6Eji8UhpGD1pTMhkMpVj0q
JxFrihDLS07jl/n+KKcpg/kY6LzD55FCXv9ZjFJwLHujxaDPwkTSKXC2OIKCgWaY
lBX1l3EBzHc/ptn+6tnIpsnJ10hTkkotZGr/qbc+wd9a4C2aZEl06gFvH8lEAc9V
gGL0GWas+p23pkyzs3ApCsLbMqVIbYLQofVI5mDvMg7BhvHLmz3uEnH3IyP7Z73M
p2Ku7JMq6tBO9faEM+fpOb0Rdc8vgu6iUTOOJkV/inbT5Euxo1kPusHUHdB0eppl
ip7Je7ozYw6hbUuMGuSET9pG2prnaCst3N8FFEpopN/v82XUpwBBc881Dj+gAdW7
hqBcPob2PqbKHFniX3bXGWAV9sx95Sj6+gtmaNBII8RZB8mmEAde4n4ZvMHiKvGl
pVr7EBctZAz7YwsGR5xJMX+Ye8OmYvR4DVxG5/P6ow3VaifTkZv6bm7rn6nwe0+4
4a4ew0Xoi4hVd9Gxn+ZJ3Eu052f1tEAOdhHo2JR9eFu/7hu6opEv9Jiat5zRsidt
6Ij5fh5ebdJPizu8weH1Dm8vIqGm3WRbQhwLPOFEmwY7C6HsqDwMlcxY5dWeB1eg
yHNFNVxnh2mxNBf0ZJ+Fp7ZCJlG8feiBRdcW36qr+gnpwCutWo4XxDK8sQiXve11
uqtqvIZuHLh1r+4f/Cn8rJ0B+FO20x9oXP5C7DL//sOCKRNKIMnDi3aGZYsrMgv9
5KsRptTJg2vrhs5P6D+iK6VWVSuqRHW4g+tipy56t2HZOlxMjFuy7ICsFk99jHem
c10CSUZIgzitx+ihHsXbnRAyOvng8WYGdu+Uhro5NQxFyKNhkTE7h0xZdSndX9fS
nVK8MS+Y3kHLTsOxbZSOR3s1pHx1B24V8UsHm/xI2oyoLUbJ4UiJfLeezsFBcE36
hoAXvby91BBGHa56ILzHgWlzit3sW7XrXNvK5x7gqdH6LOYFwY+8e+YRu5RHxgtK
3GxwiayKHQOIy6ncwzvZsxy7yvFEK6s39GwU3tmNE5A0Ck143w0Q1CVdIFQr1Fj1
if5/FThF9d83mlhR9s1Z8BWgE7is5uI7J/b/VMmuD4oPc4BhRRo0QJlXu079JNc7
05/avI/VwnNDW/eA6wJZAD4/1FVLoDSvP7LJ0UgjCdA3gtpnSaDUpreJVrZaMJaz
SkrKZEKiNRErYS868vGT8Glw/aa6ldE5nX75R/ulKksv96SlLlQZaDup4kAnj1RN
5I7XKEY6uv4FOcmgip87+Qe5tSxed+dYFzUqD28DHFi8yk6/r+rvT2w0S5sjRI1a
MgOzWHFAw5U1kXU+X2sh+QngOPnseeN2aQIiW8OAlW3Y7RzTbwZuk2XfbeWNZsQU
YYrijchUpJjOVvBM/YCDEGqlRKQ/TOa4WvTEm0GXaDgZ3N0omyUF7ZpCAEr8+QkE
iV0Bd3GsgnJubD5YZyHun0sbLP4HTO2HLg4fwZ7Y2dmrNla7uKHy80055h+Yo5Ub
JB8/1xw0yvDUKVp26DBYVfyx0PcmgL2Dlw5zP38YuY8bYw1i/UaP51axZctf+ozD
2tUGpWyhg/Vg6oypMS17QRE6InMAQG84JpjUD0brLPEAo9Hwl/gFBcJjmkcoe1ME
kRXnYi5vccZgn1vk0PpelLGWxKyhh5xCemTYfZSsB33fb9VIpinZWFb5atxCR8Z+
urKhCLypGkHhMldthHVDKzV2tXc8qWH33tbYT53al6KmV14JELneKj7HK5uaRFrU
fnAAjE0BJ9TZj6u/OHNute0UNc29kLuOi7J6X/+Ofgfg/XRM9Cl7Xv/L4zPNi4Y4
YpJ+b3ZZhx9ery6ZKI2pvy7fSN1lFXCtU7Ryi2y1xUGKQwwP7NT31jCQGtWSkeh4
iXhN6xc7AscFUlAFHjojDQ8Aea/xintdC2rguZWoIzKJu6D0pQD5QfLdw/BBtx/4
7OpM5MP1Vdxm4UV5B6ifpuGsaQPLSukBZ4YAUODC4jZnBWuuUEcVx8kQlLVuvBqu
YY/tzFevWgoGty7AzMh3SzGc0nTRgvkI5HHPdguotsP9i/IIWdHduf6Vb+vSWQnc
9zY9BduMTOxoOu29fqRQcViiSoj/7KyTYtvuI+20SJHa6Azm/GdCfV7DULsUn1V5
MS2d3O9pHU//EC+8h3IRwQgw9X6v3CO3SBP8C22mZAwrBsVsyfBFrVz6dvBVuyXv
8oaosJEwXP+DvfPGzHpf2lG1QUR0Qc2Zs30gcBAJKq3gYBVO256t5NVBeizJs9jB
CHEwIS16kI2gdkzRZCAKwLC5yPjX8wplqv+Glx06gYTFeFxsM0ZYsoLr1gKaeBad
qpdFLp0ypzNfdMsim1mOsCHa4Zmg6ANhM9SQGs/8pTVuyCmrhVkGlxs+dXY+Rza0
T6HiyiOLxD/IARUlqyPFnB4BKGesfljtrVx1hsY3kK/NcgPpEHLpKisI0nWJtLoa
BhYa2W/w23AK2s4uuTBnCMNXPcycgMmWFdwMLETVEGOcubWkXIiKVtc2vtpShTe3
3RNplV2t6zR84VdL9vcL5fVC45EPW0wjK76/FuomwP8cyEQC3GI3tIKdk+wM7WU5
ZNpsVhtX281QFfe30DL1OoGGwdEwfdLDoxVQ/V2J94pvD1L+g8NNk+olcl9xelj6
eDHYF5gX85LEZ5CyoKe6KbbSRVFHyVcSF9UfahXFHAcjUmPiJIZZN1JZ5oJAgQQ4
8wjMTTGMXk79X+3+XzLYgln8opmbux1ZqM1JKandKSPqVkyfnQsxeygppivmFMsY
4X2KC5k0klRtMgBoXcnBwUpmSV7OJhH2ChYkOEep7L0W4A9IqJyV2GXgiazMy6XJ
slVLpuyPb0dY7GxL+5sn7N9y7cTst9nUi+/z7raYiWYczegIwUu6YZRKtyXJQzp7
BfGP0Ds1mBU/NWwa/4etBx8KeZ/w14sPcu2hH0wzf2ocf6XKwDNA2gYVUwC+Hx57
K4LuGmlnfxehbcUVEGtNvhU/CNaHG7FS0+/1p+0Zwg3iHrp5m6iD3k2TXX3X4cmL
XfAOU8iasnzIpQcLtN6uDsiUDNtv5pAcFm2sescRVifI3LSsvhtFNhRFnCgSGILS
JP9O2OyMYeBiGCRJv+M8viu9+WvNfafZJ+VTlNLS0LUStoRHqa2naOg4z3DekUXT
4iOSpqllRDvrjxXsD8e9aa4J8QLz4elCPnt8JobxjVCRvv0KyJ8daPfW4A25Gn+r
ZU+ImpNSXMaUgqsTk7RqoLFa+L0cUoCFZBxbssP+0idD2hagIRdRfXEyhS7MRdBs
Wx0hPTze/mF7M1cJ1mfLpPUfABA7WLsHVjXLYKsBniOGJKPSjX6cqDDodAPeYWv6
BMJkIDzl5oGionZzGIp3Pq0ettlK0/x+YDK6p0Q3Flno7KZJRHcYZD6J30DsEtxW
G9amvRcMHO3nnEYljFqpewagDbmlisN5Bl1a+F+nlRH7PK4q4m/zrD5amOdp5UTP
Z/YfhvuP6t6CVABQhLnoHVUh66Tb58pC7gQvZpzVmMcOh3v7Yl/3xuOWHh9Ya0g0
7BrvqFqw14TDDCgHvmISaXO1HrMO1tCVNkaWowcUutM7c1ylsvyFT356fwxU0rXO
0PF7ERSygu7tTWdh6K7ZF0RyQIlOKCv5cefgDhtY5kk7I6TeWzjr4uLolv+AqPni
V7kVHnJ6jLzKCfyW1vsHXLZjLwAvkfdICGP99raZ1IdojHjoNh07by3KH1271OJa
X3glTjcLJRipqA24wZRpCfvBAQLsvswD/adnmcnOpQ1qCsSFAReZBCdW9e8US8j5
bIJcAhnwzyFy8ZaJp/qRrOw9ZRto2S/ZY41cPg3rbQ/CXMaGmMxblkS7Ar3Kfg+D
AK82fxPRIFqvtdezTWkW8KTfYjV7/eGjDBrRbaXvIfWTon/fHCswuHGOvorTRk4G
hJwo8UsdUbWxh36s07rvftMsAlmkk+fWAT4KKo08zobJS5WIk/TjhRnU7xFgiGqf
bWphUbxHsrwaIP++tKHLeUkT0hdm4x6Wxxsx4Vtq7nWhhBTjpqzoE09p8EZmhemy
xaZc4S7G9+VK4cxV5V3lfHVuQUnXmVFh1FsI6FxkhQEAYU8iwHSfxORTwsj3r3eb
iaR3WMWmPTEf2C2XURyeQXIQ5yjWLnNz3ytyOgl8uS+Dexz1qRA5DCUTQ7idJSQC
F9490x8rmT06N+Cg7D49ftZAK/9r/PcZ7hwLVJwqDn28Ax16FbpXb/hqVO5SPcP3
q4x0XF2q0fqfBck58wfc+w5dgqTYtaagpzsnEfu3e/yRzlrDE9QquDS7FDQ6WiWe
mZ+EKaSadiVI21BjAgNixNI8c7fmeqrxcCjjBJ7hRD4VZ/qAjr6cqUmumb6/nuHA
skno6T3c7teLD+e12kHqGzkgIRfpD9uQ2N06N3N8aAVt5NpL+pNH+Wm4o2dG4rfV
Uu9odfjt6XOHSDf4QrqcNGGCm4J8LlSrvqPkbwkLHijMmwGSQUrqbK9oNwvJgXCO
317Nf7hLwuhPIWLdSxgkAbOcjAhmLdA2Aq5IxVzbA0SKnoremFidtlMJemHVAM/z
nEzM0brSMAco0bbF8evqm4nClZ4DFyX8WPzYaK7E4DQ11ODmQjAYWN/aGiMSuS+e
XnGlozKsuTQo2vfC+MicCiH3zCNDt4enZ/k8E1278qgHDmJe+l8E+HQBFMQy0i2Q
FhOcEdsfTEefMwReY4WHFFsJQTOPeDLsyJlHoF6Ft/menjd5VUDvXqWqNamfW54W
yQSDsMxWTK8DHjvUFJkqxs4xuXksHInGhN+aBzUstx5FbbbQp3JNbQL8px66QhUc
UWhXy4UXt49DaWywFuMOLs2FeMBlldbTQTOQCBdA6agK5AJHupNbIW0T6lng3Xas
HKvHWxlRMdzuGQwDpIfF5vlME2Yy1sGvuKOuj7QM09N9W/a/TiVQgBhdIVHSoKSm
8BufzLUwiWfiZsTFx29fcg1c2OTjbToOgzq+tzajn7vGiyUK3tjZMJ00JMEMIhgk
ryzfZnQTqEdtkRN5s/ypaxL2Ttrp1gfCmbopGEpbrfvmlwvpP2bD16f8mDrjsBw1
ky+wJ/BnjXzlNIDTWLjS+LfkPxMFmpZ2zsdpIrFwxnOsuJ/aZ0iuwwUw6dhZ2uO3
oxgKnXXIsx2AKglagAvNP6iO8/H3c1tkFS0JvJGVc6l6Ei5kbQkgVgFB6I2a0NOJ
JGVStWFGdRz6mD5qgjheo1dYdVsfyxRHOhqKgfsgQEXuOj0f8uZbhHaRp95/vchC
zuTnFDqAjOlEbBulqHNxCZz5dbfbRyzPRjJ6RX27Rg13pR2MvuVGu+liU37ZUwHB
elwGQqjSd7nr8goA77qAAzlWKKauxB1C479aTl6rzTyOTmsgU70yvHee+y8+Yfww
2tWOo1n/7ZJ7Oaqfx+1wPSqaiOlWu1SuPLlCIXJDeFTIt+gOulH28WnnTTrgf2y4
i4/yzTun2m2PS1vvczQ/9TzyoEY3U2gJwVzzevDyFf6YCWGfb09Fi7WhbqHse+gY
9OkhM6aYTKNmyAesYBoz32UZZ0y7jLf+DjfhRhvLXw2Wjpvw/Sk1tIWGg4usnaBA
j8eparQ038EG2jK5gQgXoY2aumy8ElC2AS2qFfDvOpS37xSPdFWy2gu6r3+yW5jq
G/t5Fo6yaqOgZzfEtrm838IhX7ZAPPXN/qo7ZquE4tLDHXtkDRIppQNEMo1RdIWI
XtHX5HSH3YbQZHVcwGGz4IRhoAV7iuqg2iBD36wNfUqF3RFf52epk/OxiuU1w637
reYJ+C1XeXycIlrHsgcvV2CXPiT6HfIzJchtrIohMAKmxtf2MzEaw70dysxo/q4k
6+0K8I7cLQtWBTcPO3YlwEPRT2+jZSJKUuoP4ljusI7Mv1Ov9Yue62KFQNMGyKTN
4gsF2/SOersWuzNSHLQzHu5USX3qB2Fnqjbrj9/cLUwVs4gjLIOBc0UhnDhyMVlx
UtrIlYgD1jusmL8WcRctttH/ZuDFZIIdTMh/y/1fD9SF22sn5PrySq082kP6Hbxt
YSvQinP0Y/pcjgtoO9/nh168kNmATcQYbunqfYkOu0Ev6gWeG+lrioFjZLbL3hCX
Rcb0sa6E5kqdb7CEV8K5LWKSRiT/pp1uGEqckMd07F9c1RJGZWKIECr9utTxGwUT
RDFWVe4lfO4HYEC/l0sHmvXYMXHCm32Z0celAd7gRgnJ8XxWkoxoOG5FYcJIGJKe
+5t/LP9bwyzSkK5v7hcQOUDCFU51ZfQKOM8WlAKan5gWCC7Q2d4nhU6ium8++TbW
JqB8Q7Zr0ssd23IswOJqXtN1zxLO25PgNhhUqUZbWNWYROZojAU7bx/IDYv1LOgB
6BrLN++nSO3L0A1oJgtQlG+Zp7EERcACjpiYUCDEQLL4yhoJ2PvbyJgEMQ5ZkXO2
t40SaWow/CKgzWCm2OjvKAlmh1xf0tudDc45UPhQFHNzKlQXFXtTW99XTIEQ62l1
NCwMhC8INdB4WQOcgAOStfA5Kq27x/lbRoxs70m+qpwAx1q1nF5zzs1LAJEEIJ14
YRQggwFyApFbSdny1i+xCwl1F+hQPmIQZ5Aqaot3e7NbXAsv1Rfefm3J67KoZRkE
b5HR5I3Pv9P92NCc5yeVAilOeE039oSYRq+ieP21WeiYXeYeTv+9gRJqnKvHchHH
mWH1HBRwverEaIv0Zhw/gl4o2o04/X4ZCGuu/ji3eRk8aGsK+guFBGhrvkMfR0FZ
/VyMPnIZJRpSSl3YhcrrifF2eXwl9I8qtXo85WzYsdS1ccLFZyR6HHAJi5KgDBPF
5m/UGvpcvY4c0mRU3cPsjzVLh4a+45GW1d+fFC2ARC9u4Bpi7rWwJuM++CvGOfzP
ajd2eZDsN+A3cypJmuWFJGZuZ80oO7oNGqH1krOPDuDLQ2RLTh4susrswhx4NSM4
IHvGfoNCtuv9dz30XnLk88+8/9qCI7edRueQnBbPdGH0s+uyfQXIFhwDbKesJq89
6t5QdfBf+nAEk5o8sP1DHobTTVGzEqhRk0jEbLlAHdSp4hviNhrdxQhH0G5BqG9M
OL2Py5zKDcrU31lSYhoJEcsi18m7vxbl23F2MvR2+WR6TC98z1xzXS+TEi0O7a0D
gdySdfbM+2JzmNLtID85O3VqcMr6A2/FUnnap9wEERKb7NUnns/VbfW/wYFCvsD5
1zbhBxrSWwf3ao0vqPxqYIqYkb4EUvhdeCBvsgneCgpbJx4IU6JKmmAr7gI5jyoN
Ms3V+zUL2lBENtkBtX1EMLJ8LEwtCvybl/NpDmiEA05LDjiobutl3N/LtQ70JoEG
Nh6OoQb7EqWhM6AF92lYyLNyLJgSKPeIUIVMd19Y/Ki84XjlenXec8uFufrGXV+A
jz2oJNze8FMFNAeNFg2CcXLKKvPR8O1EHqVaCe0eqnf6gZVocpf8nTFISkuDJBsi
kFgrBP6o7+dCGiFpdZCxlUJKHUNv+eZa2e2qdgB5kpEE8lE18r1nESvunFR++Nkt
P+MheWEjvSqp/D306U09I11mKG+/drqrJtYpHewqaW2bGh0qgJ78VOovE9QvTdrr
fp8mdz1eFq1I9JKlecxhHwjDpASzqwPluq4UX6kfWaoD2zAby5eU2bHSfS0JajBK
O0blvxwybjRtUxxuOehujTyI7B47QOBZc7TzI3dgM9ZCd+1T9UXV6sDO2xFhbAPa
wzfB0sexXdNfaW7762jf7jWk+1Oz0obupfZr7GiW16T365hSgQbB/HZBPhXLs9cm
+B0qp49YI0N+MsHDWxLnCwuHl8K9dd5ghRrDivLoB0batHabmuIHf4A3i4k/gG7X
uk/8Jqox30qJF/M7ixrDjGlQPajJ9AK54SLMD5SguT7zFGdzh/Hr7hNVNnvUcUUr
C4QWo9oz75JQI7zNSdOVErekTVE9IGw5gaaTvFfNED3O4XeLqlUoMAABTwCcOT/z
J7ifKYgD6/4D2uiUXL8j9TMumcxcOzYCp0WO4H2JimQROoIxdgYOPOT+WQz2sIDx
3quYCQCx47HZyd4RoZk70V9QQ6DgFUsYZKz4M5KlSUSMAvZ7GI+punjsHvMwIjmR
Ry8j1QFfRzbVA1FTgAGQxrcAVcy/jXRyIF8ZXDc29rvpo84oW2qCsPQjkIxTy7Nr
ZwqP0FWFTIGgixr8ezwb4jR1HHzkhDB0iWEJf9VZOt73F3S3VRJzTqvQfgE7NVas
cC2N3uEIKBCpUXSSq3srSoMLyvQm/ShdeQWoIwLq8yjwYqkTUSuRsoZ58jGka3Za
lRt9xmbZ7/PjDuUmve4rpqehp4qX/g03RzJxpdkOlHXPkX7Pc+sTAntcEn0LoqH6
b1gaHCfyAfTENY0SJeM+Po5lSHlwWtgS2T6dHdlrw3oZmwXxEvb2DXLuH2xg7oco
4NyGa383rKucfgs6jah3fDRmMA9ARxhEtK7oaVy/fIKCEc+D7wyay3jkJ9+NhEcj
MELweykTIpeVgY7aSPdUw0ztROnz6LHj6lyILD2RoMwbsEdvMKLvTajuBVCU2fsr
IsrSj7XVTXCW374UUa/zjzWIh9kp4OwyBhW4cdkUud1CsY5XzcRjyNWqXcyEO9BA
XIGHefJpWkx5nVcYw952LHC4q7c7RpbPDxi6PD7SdUByx/rKtU1QctixD8FokPHr
Erl3m473F5iV8VcgtxzGp73NeI7YMLn1S4EfmcQJQgn8e2fuIVgQS3tnCgwu9Hm6
rTGiUNtN5eYN/WDDdsjBVUOwNX6lwGcqTvbIOfZSdx/nl/EKA/3JwViVPWz6jqVf
4BUt98EUMUApszJ7H8aTXVr7CPMnHIvMfHd7/X6bkb+HmBOt36rmKMOpN98w9fkb
opb4/4pcDgu00yuTj1/ZNty+7URjpmEWOm8m1JCY1ICTlgzHDLvq+rb6gjvfDJue
ypIyZ4cavXctEbtL8bAFxjX1/S4IEJFn34f2pJSORC6UTgjttBxyjfFzKlQ0Cv3S
NKJQaFRSDdeEKs5KkB6G0TpVSa1SSCT1kHs7Oimna6ZvLn+rsT1p7rmlQwxWZE7z
eASJGD5VUNm2lhBMMeiBQqy3qNEI+rhHF3rMzWcb3qzVrxu3I108NQ9toLu+cVSJ
qH+NXNuRlKowUbgNVSwuNEECRXaT1f+oEZQU8VR5VwAVUrP3EcZfZfk2zr9JqYTI
+f/viRyy5MEbAGa3wmbrVL8KK1bmfSj3i3tHnRACS6c+w6HYtGklG4PjBXcY7icm
xqcShUu0lvTj+zTDKEwGTQefeGg3WzzXoH+8096re5wz+1HBQypSbdkKBbw+6gQL
VUs6YuZWr/1/DkVy0kX2/mk1tGCqIBxYQRrGwa/Sn4dEOailAEYpk4/fMQOAdcr6
K2K7xADtgFBniCKbBR4y8otbi4Xa93ct19KgHwJfvMJ+bKgzATCVwilctsKOnI0Q
+JNNYSEFaJ+ksf/aabyluoZTC0or+3KztO5G/TZwUlHShR5nK2NGE4as7F6yQLoO
6LGrYXJe5z8/NQD5z7V+2avrLchL21Pt8avNmym9yQu3cYjxIdZDcCY62i0UvkXy
PaNVCPI+V0ocflxO3MRexrnGxEdst7TkgBsXq13WLzmmhV18vu2b/umZbuOiU8jd
UfY4uWfomh14Ib38VY/RCeZRRirDsN5eGJ3FSlVjzdTjmmaael/0eKrGWaodbTfz
U+39W8opLNJiQW+CkNW9XZDNUlhBTuYpmTuwWG5GWdf0ewWvP63pSo6Q1MrbDgot
OjeqlUz+SzBbqh+sYaP2QCcP1L6dbW/eJpo0UmX11nhlwV5dA0Wxa6QKaVONqXNP
nw5Z2+Dw8+Lk3KzKr6GW6m+LXjA13I8pk5/8nN9QliXKJMo9OAeUYpbdLgG1ZRVN
P3FyM6F+Is/6AMcsEf1nlssJPOuXcd6cyGV9DxSFY3wCQFO7tEjy97zK4vq5II9y
wAgnJ3+KwhoKV6PLxxfoMcEg5wVJya3VTTD6rOfJFjBWtV057hnyheE6owB0JhdJ
soH9zYrh17q1OamCQkOqyYg4PO1kTfTGl9ipseEStKWyXH0v0RY6bZuZQapvC31c
QVKrk8AEYnrBMKPQ0XQvKoKMEcgtta6LlvLZjqFVf74f7oL4Px1VoSOuouCyro9w
4ieQcIAi3nVEQaQ8tD2lYaIjfPOJKlAlr3NzHexrX370kbxMNQQSRgt4KE9qBP9k
zdUzRnimGyjvsXd7KOZsYrpep2dwZjhQxCcpey6suqPJJdZPVa9nR6XIVngqN49+
aGQV3sbwLyd3Nnkz0OoAjZdJO7V1y97QagH+W3nXSW4RV7Sb/TmqcspHJzr248vf
DDWDVmPK1oo+denjJUDU9TGcwE3UYrWro+0WTIGkxs3yPeGoCUhUqLJSe8ntSntx
yNglLXVUEy5l6oTxIabB4jqFagEvcOraEBG8qmKC8Zk2u7tkcoFIh0FW7ZW9t1c7
nPj5FTTNmvE5AxUGnH9SKdW+RddGeSp4rPYgFhZwc46npowN5dEfv6B50V5i1HTD
irVoQfACckLEYPKhyGnIQBp3bvl9OTArIaEzZqHaH4WnzVz9Obt8g16R6jjAyXMP
HHU+XgYkre+q+ory91biKHfHqaTEXYJQHf2aOzXmWmzeUoYTGwtE4txOLCWimqti
XIjzY1+qCUiN9NV4KToe+8/MLnV/3Bof0bs0biPiLqV+HWadHzSOozXxSLw6JKSD
A1/oXL16/157xZnj3MUuEohpmdw8dVIo/n+SvFXP2MLGNfNAKdm6tc9DJMs4BFnM
9rYXeFg7ywk5QCDAY0OAMJ+cVCsHPchAPdFetf5s+5JBcJSGQEuATsH4hwOE2V1l
s+/rNGt66ofQAI49VpMoyxlhaAYa7dAaOOMU9mT8H063FNagHFOAFZ7f3JUQKYFI
A59odHyig0WGh9eGWct4sphb7mUPfH/3Zmi2D5yIE551U+5KwdylSs/UszIw7cW2
tzJKCXNB25iYcDpWZaxFPo5yHUELgEvnRKbg2eDCbPpfpkpIwriOgHv0v1MRzeLw
s1MKBQuOjpa4hXanWziuzTaelnZzPAxj/rz0YokGLfB5mMf3sKGkWLpzhHyGI1gm
HRPLg4fqaNb0drEE0upBxkgi5IF+vIvkEmqEiAtHRPVLXxprgAUf3EDsBQFAPdNC
hJM8EmAdPEva5BHH8SIKZC2X898jmqWtRCKKHos3rv1+f7FVLnMAT5ssCTVbVdd/
ytHhBbLA3mfAbFr9dUUOT2GCSpj+SIiA7qcPhmMUeRvwZ6Xvej7XvyYeahrCzpGr
ztkNNsf2o+MAXphShZ2sHUI/WuA5hqj3/G+dAFV2ByA9nB5mdJTGOKUyz2XPx7Jr
LTmEhMY+FNnd1lU5f5vqswWAVhUDCf6T+rfK/5kA/9zDIAtMzQupI2nza/vn2fWc
vDr8c2XuGE/tgkNKqTI1Cu+yshZJwzrL4c7VFr2fP9MVMDjcZ10yYlxONHzTf0Xo
6l3uAXxzjSAmYc/nwVSP8p0tVLN1bivrRwOUQVzs3PFWh7/njMcagqb1qkcpbJHQ
HBL3FAif6SbBUIDM+uAG/2e7t/qlkXNBhiBlveQMIv1pFn1gqwDXVk8GqtbwGitu
IoQ6Cn7H/YwJOO4Ntenkv3aC50KsMaVlhG1FSfty2Z98iDUNCL21m9Mne11OG1eA
uOc55JccoBmALL6VlFNZomkauVu6bTe2EBeKiUMlCqOvuMLrRJ4HnEqxuunRWXFo
ttSkpHW4BHsaj4YOwTWGFVvPoQGjnbiEx3aokY1YTwj4aPTo6nE+XricmwfNfuM7
IWmnh8PQ9c/KFIuy2OC/vHAL5bMiORbxEzN9L3ca1+PbuRTNPDh5w1s4/hfL9SM+
h5EzCLkndqOfQovYQd2hFBzL966Mol+li3xs2YLASADhNmDznIAFE1ShuvwiaNO3
lmFxpi4RIe8+Vku6XV9Z3Yx+bTI4h0XjNKFyyRh3rk5bVPOdsqJj4AfswnAnj2Ss
qzHXfe7Ojo9ZSu6qS2Fpk2XUbGChZLG3C76OP2okLCs/Bi7RuVSZ2KlsTEjn/TEr
P1wSejv7eVJUV2TKYhFtjK44vydFtpZAZ+6NcyC5ZkV5eia+XnuVE25aOa8p4ka0
xkWa8FQKOVI8GmR+t0k81BxaYb1Dzl0MSKGiFRHk9G62FcAeLWpaC/QTkqlXfV46
3ywLMfohG5XLA3eL/KLl/zkTNH9l3YGhtj6/ZoZWgmIE8hpfqkc3VBgjuLwRTmUF
OZV6OQtVE7fgOCA1utkawQI04jJmNasGji1SVHsk3+riQfXL1UiMPlVjmOtxJEsl
8yF+5XfTC22pTiHMhv8qX/pPjyXh/hBH6bQMbHv20m95cfg3CRFyG8qyBTS99Zy/
u3IBl2EQb7lywT7lOrlhhR9NqmqP8uZ1hICR6uhHIdMj0pkLLEjcvAo6/R73AdUA
UTvomPBMJYe6diu4JCOFCeXXTcMXmw0W1aElPtsFZ8dWovmhPDlvPakZAYLo/Lbu
/sVjzvrOpXLLV9NFv8lWE+RwDx0hTNM0bc0WItrKkZi6V6/exaLcRsYi2AW0w4Lp
FBPOzK6kFmrpv+7iA9U+mA0JBLBGgCWsOe/CkCA4gppiOzfmDXkVZG0fF2IefyQr
on8MYIKkRhJ7Gp0XI2xfl3NYBEjpBRXcOhqoMVMpwuodumtGrSYs/EJIkE/yUGY4
XVv4ElApY4QUxFO+/Uf4i+zucPnkqM7gQ8aFT7H/Ql9NdYlds+3afocEn8zCA9sp
4uYGWsxQxMkAvXjcjViOAvRA+g3hoKqfcfyoY3w6aRF7SLKjYS3wPQxmsiq8Z2QL
lQiG14O3XOwJWP+CFbt8qR/HMQpHflhHzgCUhYtE+ubsz6zHQnTOLOESNfko4nIo
9AZXtM0biRbP49qZe94uaSTRiCgu1CLFDOzY70SMQcHEoYJQFwTudrMQZpyymEPY
D+yDnkbCHOYZo/dNFwgts2J89QTz9DS/XDHi6hkPAqnYpBItsvXh6RarRYzXDSE9
BydD6EHlLtJn1Cs6XosKzxOcaCwmreWoCOga85RDOkAiHYC4sKYHyGgXVJj2aYgk
KvUSf88gvTUE4BhF5euZg+cgdNSAkLGUJ6vOVLkntOwi3Vqka3+hqUCRpdz5mMTW
+BjDRGHARtWxy6XAGEwLt0pooJxH1ZPUthEsOt8Q0EUHhWwWoRww0hhaQDRjmbCl
xwMWmdWvK3SvkuzhX7/JvthlYaWiM0RPWH9+fkgpKydtjtb/okU2GyuSqecUBQVW
/ocy8z30KtPYtmvxpqy9Aq9Q62tA/WwiAz2YiUyhPwjj9YBvYa3g/xtFyGEaClSn
odWTiJcdHWt5JxbgTM09iMoEEJgqJTL53bxNKw0m8wh8nJcExUklZl+XhwTaRMfI
WBqTKscYUssRmR5pbDlenf8raqMOEHL6fW6TV8ZqCUyJAxrlO7+2Baahrfg3V1IT
09YcoqGwPn/mOsEnxWxIhD1incBzysgT3wNR2b809smHsBjjXs7MC8x1ZCNpbR+m
GFd6sV9YKzZ0UDmtVg10/ivh4vvcxqTU0pZKLCewhYtf8hUsnFrP4mqoi+2s2AOv
Xiq3GAnvK7nLqpOw1298q50kkshJNjrx3RCfBAv/PXQC1P5Fp/vBrJUVUO72JuYq
vt9pR9WH16gFZjiCvNah3aGLREMVLjjHC6P0b6UN6V3o91t0bBzBGwry4Vu0qE6w
YERKMze/8ie/XXlDx6Zs/YqpMmagBv8Kj7NFexV78AkE7HwcIMryHPLN7jh4qzjR
7dh9LGJ/C+QyjGL1UC7LaNv31t7gxotG9VRrkLlSfFCK+2Dx6IRGbS0evn3W2ZZn
9ic9e08tAvNOJbsdIO7UmXRIyNQ1Fw7zflwcAFjZFRaUpAkEwyQRZeZqbKxakNzM
o2a+Z+zZQrxRN+cvXvooPgY34OPiT2KUNw2+qNnFVD5lLqfJG7ReLIjwR3K+rOLt
uw+orKm3U2azJ3oQHmb1/9zxsQckYP4UD7r8RaHk1zDULL2TPubmUlImHyoBHOsY
RebpkNrIJ0w/9lKuymuq4DzfHnLMfLvPefYO7rmMa5SAotNt0vOc37SjvBa1p1XC
ivRoIt3QiVW63udFOf5a76NTJDtnXRQA+KABJTLfgwOgcEfcAru/3OhJX2XBjKGY
dH9FvPKIF5P5//iohJtZfThXQgnW92+IJ52i68wy1Bxd1/2wSOMCdFIcVBXbOoBc
kUOHHWE4Lo/1cUP6L2o//k/mxYOtSIvyMmkJqPVM4Ikmo+d0t5lnXlXOwpsp5pIO
cho1jSaGdw6FlGB9gz0u30+qOsOhjI5Gbfeg+G4edEcgg94mwYa/eztWiDHKrX72
+rFk19+RLq0vFpkzAYILWwBVuFydIdO5gNnwIHZNAtvRboY81CyRPGd4WaNwJRc5
cb5Th4aOrXBF6wn39KsnFxkRdSZsIwJFglYa5FdQQ+xXbFa3n4AV/grA5ELqh7Gy
m/7hZGlx0ApqlZdxlBvrISXYHWVJyKU5wSSBmV7BhKBvNpSiDy7VGNtiU9OaHjeR
zWj0t7ouw+/tCDu0kBjYhjpNqK5pHzbvggXQbu/yFXZVPBaKd37vxdXlbKsGZ8oG
YveQkrRA5Hc6YF++vI1Tnjerxufvv8EDiVfVt4kWlPd525VOxcPxFp88p74ME4jX
jsa/KdKwvtTZYnH2eWMsiW8EeV4Wds2DkW+ZTsKiB43Upz79w0CeFVWef0kyvx1o
QyN0FrOGrDjxUmkB/YPvX+SYCrVfLrvTWr1GtsWIKos76EB9awa4oSNHqWW24fbe
xviMZMl/mGWTNNJtsK+biUvKIKPB0yZ1Tt3l9kiiLMw/U4+6ILX6PbAwY1OkfWV8
YSbOOUAgGObFaqmfpzHIZqOGFXn8bqjuYypACX9AnqcoLIxvSRYc8NbbGT4/5PmC
rlaXt19WegxtO7N8rXxjkUjHtZFFKN+QUcuOQkU34Vx2X1RWwhU2M5xeYf5mdzEF
SMDT7VN7xN2KE4dzx9vEPTBsqh4IUJROYNOO3d1zBcfdw+IuLF31HBX9knBIFgi3
z50vTl7uxImxnaLUt4QPu75YkbwFOzyboYtDMdjszjVMVkVl9ZAgnDCuaJCpqJCt
LwELYXJ0XoWn+ykcBRFdkAXegljZ4g6t7wTDhBlJXcKr+8nZcgGOuKdhYutCNqGd
mL1cYqZaUqYEOUWZ5E2YX+3wAswooWeYbdsIQoiS6AGkVmyNreZ6lb7QhRBtsEfS
m43nJ+vLHVTSOXajVMkYJ/QLsxFqeXen8+0aNSWC/n20jK6JbveYRK0iW11tQyj2
mlJekFOMGI2CZ4zOyNpKIWiN9+pmVolxBvcopJiq0MZ1LxT7oZlIvtOeWH5DRuQk
L/Y5gYauBvbX9P8OTuIbLDHIzmlnDcPpPoy6Ji/n9kAJvRwQ7DyyGxhm6D0dcHzY
rEaDZOLBwtIyp43SdintfIU5f7mOmNlzT6ngsYzA7NU5NGkYRGa/0t07QX/yThg3
6rvld2oz876ZQj0+LJ2aTWWMOw7GUZPM5dCC0GpCVoAzTXQ3D1yhH/Li20MNJ6zJ
t1t7FNqHPMfP6Cam8y2RMNswpvWmKxpI0knp6KrXCTJxWNFSraEU2ghuezEw26h0
r138P6S/pbDYHPyDzzAF1HJLalsYiPUrzPWQrTOaFUVh2lZc1og/b1S7oHMHGN2P
aucaFFHTWE051YYwmLpBMb0ZfyU4sUES4ynEX2uJomK/Pf/Yg3bElir3hNmHER0n
9Q1f7KTBDspVlMSnZbDRDsf3RdwlaQQTHOswo+k4nQTUvWfgbhP/xRu+FAW3dPlz
zH76Pdd86OR/wF4EHgBguLsUKIX3rSIhI5N9xRVhT8p10eD/dxUdEV9i9pZyyMoF
y2nnugQA0gBQLQMHgIdvIwG4THRXJ5/NkEq20Qvkqm0dua4sxvZiM5+AoxABWOdu
RDN9QBsEKzKhxMhvbUj8iEAB0Knw2kJC9R/hUGR18OETEwiNYiIE3uOuYv0fPYtE
DTacm4htW3CmK4mbd4z8PY/2Ldn2P3/Bzl4Vba92xEt73WayCtNq8oZ34SELlpUL
9UhFnQYxPbmXZmySyGHE4NAMo0k+Ev8z6bjsaroiuc9mDOGCf+aJDY1l0q4awqEI
K31p3xw6+f94x1CwqfMqzslvnVIdLJO04ccj0ia31BOL1nwlQFdugQ9u5fr1sRdx
wgWMwy1yaDof6GlVUCvOjX0Cu02g8r5e4p2dT0KsQCsq8a2TmHUJVtjcQ313o+A7
N9DCQGJpaVNBv0hhO+7zSsqs+BCCbtOTplnZiDOyFZkPgneLILGIdWQvRTjPnsaV
hrr4+kbTRh7INtTtl6LvXPaWHQXy+M3/m/mlOnPcQ4YvY4aOH8fubRf4SnY6ka15
rDKy8qTGpxXlRYKmS2Nvg+jPKIhCu2beFUS5P429JuUYqT1ZyGAfkuJBq9hidxdv
VAw5JWQBPa+qNZj5s7eB0lQSG5hh/69oFrjKhuclGf/hY+C6KO+xYj3uvzqhF64r
6+jWkPUZz1l+l22Ku7CtP+dO9W8YLtLwbGnBlDu0caC09Qi70+i205XLT5+jMYoq
8sYL/GuSDdMOP0rrj6NrwdAvHkDsx+fwos3NQfDPOfMEVj/VSTvqdCn2Dmh4JnXx
EpqQoRmOGBP+mruQiqVoBA+Mm80vZKyK9Visn4y6LJQYsOzniAqNEn1tpmllhxwh
4GB06h/r+MaxEAanWeNF6c/jZxUSKsLGkDwvq4CpyxCv6bCPXMaS2eK+FDtP9duG
Tm/hhFs1Xsc7aW1UY3kuTA6vG5nkpnrXzpL/n0i7KyO40sXY1ZAI+hi0Xpp9lIh5
LirFS/kQLMDPNlXh13hxnGq4I6iJL2pZNwXe3Y2CFSbsMxkjPZuuoktlaRssW4Ke
HTilYf8k9R1blxksejn6pf2NFmwxmdlPTA+SoCYakala+wzk32tr9H9F4KXlVsVi
1rNqBFR2/BDnGIXRbt83Co4zP8rY/N6y38vPUdmm/uFS2tzKJh4w13+Ob53qcxtU
Z7Kd5F08LxmwXI/iWf/AKtsy05P/nJy5MMffxlrMRp/VoAwypjFGtimjI1DwXI9z
hgZGLxLu8QTmX7JZMTKvb3+0Ehwq7Nhn/+P04n+pYmp2c6KRTEZOahuzpB3mT0dE
7yfXQvuTRbqfc/BXT6Dm/j9j8KVSxwtv2BZWvUP1S4a7PP/sA3u6QgiqpuaFjsYh
/q3IqNENufKvdt/3SL15nNl2oCZAEsu+VdMRK59ncnMemUm0b1HSQbK1rmCKunEy
3ArFGGXNjcLIcdsZGTzzBqItDFEd1ZhfMrMxyF16f1s+JIFCEZQZlv9f9s/DdG00
xihnljuUZUH8mS8KZbjXsXTfQZb5SDB7jZSv8xILXofDzGhBGd9G1aV/dyUbn3yk
bNSzpZKpMk5rEj2TKfjRj1T2/e9FrFyR/VGxGj4oBuWw3ls1N+gQihE8emmwyk/P
izDDLaUP48rLjqKmFd7AoQ05Ua31qBg2yS7LDtlmu4IEUVgjOGEeBO0A8l5G5i0G
zO+Vk/8iQ5yOiSov+B7ta6EXrDr2k+v+BHc6yby/ucQmWUiv8nhLG4oT051xzO1M
btZFhtgil7C9Mp9vdQnTWpvRjt4joCLCq3NMPTvGwonBWnTHdvwK9mAdl26hSM51
3Efz93Zf2vhOnrrfMV9rYzUWXAXBjWmyKJNsnlXsYVRRi+3SXcF8wYhfobv0ikSj
2b6Q7Z1dS0RFllx5d0v0pd/VHdi12712r5O7xgsDP7Jz8CGAhwSxMfhl0oYaq72j
mJNKvQSdb46HXNBvpBFysWr8vYb+wLXPhzbNJbUyZwOkL9C2HZADL6gRl5WUDNNJ
rfu6EffIha4U8Xhgimvg3NTaRHo7MvhEMujXomiMzjNcpecgkD1dSc1EgmsMgJhS
pC3BQsb0wrriRItXaLbduoYDsUuzu7Hwc0LqG3HQfi53oJeJB7gpH+m3w1NhmX5I
jNkHeS3a8QYFQJ9y5ndFqGJ0LYBu19Nw685M3MGeOt1MF6Qp5dBUce8kZKIZp545
Nq2Ro9UvebOrgqAnFRUGo6lUVjRgA+61ul0bSdBOFR/8cCiBL1ZnycQVIeUNTCg7
6UmmVwCcAv6w/fFfVgHqSdzfSH6W52k5ttuZcv1GPADnzIoXyS6/xRecQlzVdA5W
GeulFJnikBsCcSbb1nbxPBbFBRrf8iPY+Mxcrqu0cXdojQcjfqZsjradyqMdRViJ
ptVCsK87aU2gLb7OQteYNAu5Hdw/dbj+ymWN2n43W/2JZbfvDhFVL4A9Nv9ir+iw
a984qCuJOS6Se3iCASaRRvZTPgjGMF1Xi8d5J+5hoko8QdFq4rqf9gfergzGxeGx
1KBbKAx1Pows8szk4v73zclU2FzJIiiWRp2evy5l+895VxAgUOxTIrtfHF7DvUhB
CttXmP0THkDi+N8dp68+O3b206xsxQZxZOfVUyxPpVku1/7ukaANCoIFm2dyZ00M
EY3SaX+hymvoQuW97tGy7Phjl/UPZiHysurG3vyqjhWjkc35VlTSYxbzxj6f/06x
IF2UeVg+x2fyEGZG+p8y9O0yGXXdZX+0ouwfRz+t+s+gNZxYNf0MOkr4dMiXxh2F
IkIqc2Gqtj22pvlLUH/eZuC31W+9N2TGUcQTLiiyIAmjMZlnKwPDt2ATxhV5G35n
489wxiqWwwYfUCpvaUDagy6RuwgQkVfbBK9c0kYwA7/UFSTHcRcfC9a3IGARg8PD
0Fb1h/IZpnPxYChkmXEtkdN64cLsyUq5zAVsV/26sDemv42CU2+PeBGisUnpIEZc
6iX5kIZ4t/GTEek7ATZ4WbqbzQzF/x8IsX0WAW/jGCHK+ZQ7AjgfVnnrmuT5Gyn+
NHwN4XOKfq5gGuTFHYdnMDk9vGjdYKmGyMPUH65lmzOBzCyDp+04CQzslUOgKdK0
hcgnM5+0hF5Perpn6JOp5kC24zTPZeRRZvSoT7NwLLFv5CH+sNZztQcQtdc4qw6h
Xfgacq+xGuwRoR6v6khCsI0nMt3TP/hVp2HMvtrYgAS18gmUIvTw2LglQ/CsPOoa
DyNtFU8y5z+csPWEKu0izKIPQocItniJAGQ5iJbYOtIpd+yQo+mMlONKH0BbPNBZ
q1oIXqBqLMIwhb/K+0n76xR1MZrXCQzSi1MSTiA0vk9eGkQq5AU66XHPDSbSafqU
Qvlj/e6SOyYHDq3RZ4XqP0mXqWO7BC2LgfINSqLlWHPYlA4fhngaz8fAELy+gyy7
LmmYkO61rNJZ1R1SV2TBcCGIScpgzi2ctQf6/z5Www+gm7/T/iRPf35HR4VAnCE3
BBSM9TDEVf9gNaqVtAh3a8C9Kk098V533YUyZVstzuiP7fZdzc6TnNYeZpttOvNN
ZZCYRs5z+F1I2n96uFX1iG5gY/NbBvflF0fARYBeR2JESti7hTJa1w4LEsMeDCtd
ONxTG13MZZRZ7ghWl2R497R26EgmOhLKdXZ8uU00EnCQyBSmcqGToZlSU9evBSWt
9WvwURAz/AnfeU8opHdsYzUc0azxgR7Gtmt/AS0q0zus/t7Tdj6Ugo3NP5UxZH+Z
jmLxm4Kwx3ZOFq4mnmfqGw8zVXVu/5IRTJUZUkhs/V6Ox3Es2IWC3+Q4v70jq8CG
oy9IkNbVBzdxjkHfMvi9VkcaXTNfC83/wUF9+YOuHm+orkmjjK8UBwIEtqbvYyqr
pJdnTYdxCZ+u3SMtDvmgoNPRVN/0TSkzvKu7fwat2qZ3tbbFR8rpDg/jIHIdyqX9
1ftADVgTTcVmLDAxE0uG1Rc5/wUZjb84iQEE8Hv+eSP/WrN3lljc1XszjZ+alNGS
UkMiSMuF9D+JBbPspyz81PcZBMDJTNn1zQmSfhImUGxIXZd42J1my4MmgwGeqqAj
lBIWApNIJsLkbPPpKHWPcIiNFFvPbVzNEArpJV32t3Cr0HrG47nM4I/bOmPDNGNR
loElxgvKKOez4UsdfI/LSSNOLCzWpm94mZDPOdDJgm9GCV1HrwPmX3FTuOaDQp7d
HvBni9vXZQSa9YPiu6xTVftsGS1MBBoJ2/ueWSNSf+CBNrw14yNyj1uauJjDMSk9
gmnsrt273FJdM+dUaEK+E4Mu7qKpWzvIJjOdWlXOtE0ph7FkrS3yOXoXKGQyO1yp
uJoY72sECLC5ik7Zbe6rwQeROSazlwKkhzpBscHu9cIV4+ppMWhsrNT1BP5EcFfg
6/bVjDZcijk7KtlO+Xu9GymAFmRhcZwL8qG1SOq0Op39iPFurx/nnnHskqLx8M1y
eZqCipyn838TxuUPL1Ozs0MLV5JNIxp85Me8ttephGd3o3CSUdcp2tMiPmNmwZy2
EWQfPC+xRO0XyWyN3dZoEB7yayCZtLq/D2mGcwB2ALZ1ajo5bfShDrUXaZVztLLr
zOvL4xtDDzb7gWlZJhBOZ1BOPBoMkF+7DLaYpl6aKm/wdsLSboPlpnRvsNZVwK9j
VwqiUTsUZ30mPo4uVSCXiOPQfRzV+uw3Vz91Xq0xrFYsqk9DFltzXygzRBbFq786
24e+3uiCWT91r5Fn7r/GAIL1IIrfs6xRetAAQClqa0wvMDBluL0JmVo2aay8Rjdf
NvFSQo8c/yjWpG5gVe5rv+PRvIngcJSfVOjLzBzUpTaA2K8iWvyKKP0mobly2YaC
fTjZcl2/7EyX0uOj3OK4jWNClQSTF9S1Dyxi8VqBJZgHtA1uTE41wBKqW3dT7qqJ
c9Y3xY6Tjd4sq3OM8IGOgfTPjEtRzme674qtonzIP1m6wP8SyPU3fjJR26S77WtP
WBcuwar7VYEL/2DHDR3DrZPKCRcM8Q4BB/OoVx1IAOKifwz5eySe8ghEWR0a+B5r
f9IBBoVABWM/hqzF7Q7Jy4L3TRF1zd5JRutum2VqTeKxGxQ3typO0ETFLUrzPdQ7
Pp8ubi/jM2s8lYNw/FQJyqWPlGDo75yZaeEsoZBINJaondqJWJGsXQbU7NrB9hBX
uDNpoviCkcM/DWaPvBb6PK2V2ww2BpXu2eEXcAds7SfqLqIPZkBpnlS9bvtQdO00
bXq1vcMrNAc2VMI7brtNtDwKtis9AU+9YfPxh706zC4VofLi73pZU3Ny258r92AQ
XNdry9nbyX0tGaN7Grpi1+7Q+LdpLAYBblfChIfeKTPopsuwmHq0TqQ438+QBwQm
5y2epGmX812SxrlWLpDJIGgQTb4BY2rjG+ketcpJUFOFhniQXqvFPR2PCXB9qP4D
tPo09uYd0Dx7fUe/JzWxEVwxt/5KBx81W5I9lF9CCL9W/4IHyx9w/uo947DdVPpb
wjYfdVodN+N0SGdUIh06x5kGIy0eNhaU7FOQw41jg/ImouytosRGnOihbYsT/yoc
dRbXK0OgyCpUJtyYB3iY7F5iII1QHmWzeg0/KDOnTyvE56NOB9yUtpDOCbbP7I0A
gnGo7kgWPT7DF/aEPOyisxCKlxWrr0AYUtOiofCbfULkJa+k93iml8BJqboIja7H
bgbGKKgJF+BGRwzlSMY4hL4oEzKy+GRpcvDNrsXj+z8S+j5QhfhEcSW3w5VTWMzO
4PvznROKoYTzDkJuajDsybYyl5Z8LWF9BJA9D4zPYZZ8OipY2K1La430pKTh2EEp
TEh8PG/59vKqMq2zXBsuFmBH2mmUFYop536fFmS8FxCJFVIub1CHW+FL1YmhgkdJ
GGIPlJuiDp8dcfW/J4K74Rr82eIxk/heHwbinjs2i5FdGotw6n2peEdcpdnFRsjs
a4jML6ivA3rwPeXl7TtQ5SyBTVda+lMmsqQsZb92/6bvmWW81bonxTSjAFuKG322
uYLsV+plQkCEjYSlB1pghrXXZCIGwZzCR1QGOnFis9BP+Qrpo6Tv5iT67r9oLkZ3
fV27iEjTbNFX5eBJ7R0P48/mmip7fk/v9lTy0iWYITLLPfQnuv+lpqD3qA1LWk4G
6PVKbx5/rsXD+D/UuMC0B5/N6zBXLN1oesS4APj0IeRj2wXaCC5ZVEgHHZiUvCC2
XozVR/Js9/pKn85dBMxflK1AD2USA7sPE7ZequEIqhhc8u5Zwq3bWnr66ZCyeUfq
V0CUf5WScEJvUXsyvQBbjnhWuvdomkkx5sWiMEnrD00bz0YuVIbVkBIhCA7e2/F4
PuKcQg2UJGTGEKrPt+u1Pznyi4TZk4evhW+KPcizx3yuR1OYuVTeBM+kbOC5FiVp
j8bHROktW8KrrtC1vG3VQfn+rCt082cZkC4qtGJV6W09d+ChpTQOQAUjk8Zviy/O
8RfAiWxKX6Pr9ewq2bLBi+xqQdapFkHCyX2C5C6RgSD3419pnmBst0sjCds6/dEG
hLT4I82kSm+SOkLADXVV7NDxza01ihLu431Bs5uLg1aLs7UhiSadQlAVP6jrTH0C
ZAsWxgb9L8Thi3v9catmaEHKhezTsXtC4ASHjhkJqPktwkOomEtjtiWecgyS0jMN
PT5oUGMem3JsKXdAsA3c7fmGGZL0BAuXdWRD77Wlll7Qo6nSFkXgA6RrxRjBFGPT
HGtdloJl8tdW4Akax7NPCs0Prluy1BBTFOqNLhprdFzK6e8soztavQKaA3ih0w/t
VG3tuuNid5EXmSEuTiFCjMahUOsoDpiOB2KMlvQNdipE8lAGk7CVkH1o8rQ2tNGp
n5KY4DberB7+xJLEoMTjBn530OCAfFWh+U1sjM5sQJipTQVn20lUK1RfgGqEdOp0
nen1SMCWPqEBrE0iEkn+VrKginEaDeBcIOVLTGr/HyjQ4k0tP7GfNeGO3czIKMm/
qwjqlxs7cbeUpBjXSSP011ayQGHVirVphRt7cu2UXrbrsb4Bp3VkI/3LE8OkyqON
TjJyIZZ4jyuzaaBfANjyWYH3n+FfuOnxm1y+mxqzL8fxv9X6NzOkboAiyNfcDDSY
nda3MZrxm5FxBfvUl4AA70dw4kYjNW+C/Cov3QeW8xnPTBfFHb1Bm5aV15Oamy+b
JrZbO4tjlrNCHLk1TyYf1wY0mk4cK6lXCALzy9PZfbMp4f3rEeE5Lj3xNR/m/6uf
MKonlEc9YH/JWSnRx2ZTHs+wJ4T+L+ABh8VZtlrpkXx74dMBWlW+fwIM2IwS/q11
5irjvGNqEre18k3bG/lwIZMPU4G7JtguOzKgP006vAymgURrfiy3XrFZGLzh3OgR
XuyQq//Wtz3kZBjEXXwPIhgEMi2OJifknd3KTubcA/zOiZynP/Lp/SiBluHxXHar
r1zp6vRYc41Xiyv/RJEYK0Pgi6e19GN0TiNnDmDKUL/iyoL/yseRJ159fETo/yyl
rubVBLp6YlkJARF416fqP4seBqoP6Y0HqNNnvpr7FncdGgIsibYM+ki4DPSevDQ6
xDBPgViBo1JcxIgDXE5YRLjvIyufwaP7kZ35BsrqfQHajM9Nkdztz21VXrwzcn0q
3bW62xG4anpsHjsDndviPxPsXleO/YCLhwGVE4upIr4onSwjc11x6/7pIP/ieRhu
oMAyojzxlzY+0bn5HfpL4qgHEDG7UpgfO6nA0Smgu65FCxEyj15k2Hd8ZLVC+Ih7
8QL/dkAdYXG34uPdR5kwboQ9vP1qhKk0lJ0oLiKFaSPAwFu2joNL4/MzPDMhRZic
HdeCR/KzgeuR9e3ina6D2aei9RRNxGuSUepg16h5EyiSAAJ7rx0XmGPYm37WxTdA
M+q8eVV5OF0Fh4bObKLuDDRVo8vI1dx85wa8QHVy9bE+bQxNzZbydB3RRUbODKCx
sGa2vAr4wT6Wjr4+qW1guD2+GOlFHBQi63fl1hUmm+Rcu2RPTIuE2lZ8Ye0uu8Vu
G9fTAWM8bqueaghqVT1F5HEOzrsNDzgceskPdtGtvbNekIzdwG8Z0eBjiRV0mIQc
jVbypktIBz41+DZNwgvEIqUV7qa2JgDuBF/FEzr9sPC1/B73eySOhEn0P+ZbyPTp
Ev8fMYDZo3jmMLoO0yK0B48YYRW1WQS6ClSnOfXFGs7rQnKM7+0KXzu1M9K+E5tZ
cY/q5ZWCxTvydUYQ34004yECGNBMb+VdWaxyZxpeHA3AmR7VlcEP8Pz8sIKdUTN7
ZTNtuTElYDG1ImPQsJJSXsLR1TGxqVyBjc+wacSZp8Uy6puCyyVZHACu2oxNV1nq
aGUM+A1m9SJAOgj3IoY/NnAjfUAqVTC0kfpIvKfGQz0qNhQBguqHoVu6tZKwGXHW
Utin8BLwD2ksbVGxcXXdvWQp62KCT4kcMK7kwowmZFRyr/Oi3pS7e2hg4tTOrtiM
UhKHAnEV/QMe/AzBMWqPRdZBRxcjSlCPJaE5uZTZTUDhAJVHae7rj4ikMRowPbXe
D91VKDQQUcUT3cnk2EzBNwdrOg2HKnMG+uFRPFoFOrt85+W1Ikj+9aCe68Okf7f7
Q5kV+ojxV5HbBScf+rD5qXx13yFW7lQKhpW3rFqyiVcqFzoDpwk9yiSozTCXKAk4
AyVLpIC0HvjjXKHsbTdq0DXnyT7+empwtX/QFmBkyXje+JmJEKircavqumYxY+BY
oN4g4jIDsI2U58iGuAeBC5IGAv1moTMOdmfsAnNvdkjp9QvehLd4tClhlUM1DPd7
oXsRthcxj1fwpC77PaEM5rlOfVFln0qaGxQ6O2Tmo4qKtA10IL6E8Jv6qrcG6+R3
iXo+IO4vb8Oky0lya8Q1z1hGRBF2ZfxGekEb86FJhospn1XcM4MmWFTLJDBcB8ng
y7Rtfdc9ode16k/jusmSXu84i3+WpsK7kIKhwtxb5FMh6ciW2FrvRriT1f1FeVF2
Tw2uBxizX9WCXa6iOYmmU++lKX5scv2V4a6i9N0pXG/Kqm2WQTK47WYsvX5qTJxA
V1C2Se8uYq4RcgcCkrHLQacM5vfw8cAeJuZjkPCizkAjgIIa5+ytu44DdtnsZmsk
D8gRB75dmenFugg3CxjkX3xisNIBCi+LNvu403itOVTII+5XzWmrTXIzkXA5Lrog
uClHG8z1DaiBjRvJqCJOWmqsK/I8DL5/uUjkm8U0lb0J5zaCSjzlR8SDjGYzCO7s
MylpMneoKpjwv85crzBiP1Y0pERsM34IY9zh5njWubYeJKmjb4STgUbTIw0zwMqq
ihrTJuWF/6JPAPJPUph7iQYu1U50ZdCiXt+oGayczPTmiwhDDmGDFNyNK94I8O4w
IUHBWC409ds62fVy4EjlQWa8WOGZwhUjVphvlvDHr7EnSgHXcdTRZVB6/g2qjTol
pqHyyWRCgqdLtRjV6kj7SWCRtrFhP9/5drpErKAAnLItRL4+bjKxceU6FzMJW66g
Tf7noOVkAxsppwBPprOSMa1QvxTgAqwuWyhHUd3AsjD5Ei56SKckM8Y6JsGOXZf5
JNtrxTyi/cw/SoFgki489RXiNP9/FNqj8ESL+Lb7275NCDmIbcJMPxY3r/VSaeQK
9w1POPZDZDdZ4FdaotkQ6Xft4pmQBeHnzKhIGGazi2lv49WlPypwClEURI+9ztRG
y+0aeZYWLynl4qtbH7hErXo7ncHan+rLdQq1OlR3xQKkBXucC2Nf5gZN5IWfaklF
oHqksyhQprAMYpafYx4I5QUUs21VrNFFLENH8fwXtZuZFRdx+otxT9jCgoBF/i8a
YsR0kHFs9NIcPuIQKuvYV62UH7TErxGZ+D/8aoe/GjAmlVsKxfr9kATKnkORVKrz
5zMfcecyCRgzB/+dbGUdAXxb7KSkC89NTPeyv2QtM0i/P8wauLbj8z7v+P18IcxF
wRJZacxNKovs/z6lFJY1IeZl6QNc4o9ENi8qx/LYCDRS/jR808IRsuveEcBbF2Ag
DPFuTzyFh8QOdG0vxA2TxmcltPb9eXXN3mNCZg3TbPu2nGrN43d4vpyEmvx0hQZR
4L6avCN+Qp/I/DnPbBgljrE6QjLvDn558mocSQ8GlVNcl5G/h7ib5sHAD2bQbhy2
qs7R+e5ow9eFMeEFASoigCqR2ctYXZ+kL1qr1UrxZK8kYJtglnnXNF/cIEPagHNi
brygyqeUDsXj/mBK1Jg1E2HCTFshiCm4ND5JGn5FI1JaY7SuixGM2k1orn69zyMv
SIR+ucsiq9+wQakTCf5ORQQXG6aXrujbxJteHKfJ6gXk7fg/BWKJ/D6Mxnnb4iis
9JwITi/Wzxlg+qVcxDlhMYHIdHO4USjUVVWJ/utVV4YbGMopiCNJc3gPUkpuvTij
vg0sGK0J+WbwSXT6slB3VxJ5xvzopxzrdepmOW2HJpsjnRMgoVDQVSXOxWaEn8XR
5e1V8B6NVNIGkjjfebz+7V0JMLNZl82gt96kaTBVj1tvK9bDDkcWb6/wQGPuk/v6
yV96p1xPSYg8PrUqw/RMgHwGARhkARoRSPaMwUk1CPWG2lfzshmPCM+pOS1r3NBM
f4ZRzLuL0+Wtt9PjB1kxT0NOSnSmRqh7C4kfyTx8Fg4r0PWabL4H89fVynT/1Bs+
+g84tDu7Dt6M+hCaQdsBM4kcSXQAY0tTs1tinKAX8S5gCTl+Rtp42UHE4qyBiKUD
vFd9XeBrXhmhZoyUUYOnguzgQzpU+Ii35jsIU9y0b+1+c4FNoGq1AhM3/RlGizP4
ir3HIS9M8ZN7H7T+1F6FL+V49SF87k4EbuMQ4MYfBk9MrgJeBPSvDbVt1Y7G/ez6
knLkTwHgOsmdeL5aqH2QeoK2Q+x39u2cRl0AoWf4PscJAKp42OlXOhJEM9dMrf5P
Ir6WO4cnB6jl4vjiI5FSbo1b0UaNCQEpc7RUtnTe8H6+rS2dtQxDjl2tEOYt0l1G
ClUcdJf7M8He1L++sS0QYFshA0I67I+DZTqMajEQ/re9NS+ObQ+UpFcsgS7PRrDw
C/ta4zdSX+goBO4+zkNew70wqCMvn4J/X0rvSNDXW/1OOAb5Cn0nfjJQZaWhk2oP
DML2agEGjnu6/paWXhgXA3y4QPLC7A7NFdQjDdR2geIPwmrFCut8Vp67Zvm/fSlS
tde0iDqlb8r25vQFMJHFASbvIvOPrjtTtRiqb/8VSeIQV5/M7oOEPwVM7Lvnv2rO
9kWVBxsLlZl1NN0DYr4oJMAE019s3IndgH9F84gB0BrGwZjgf+liJL9JB1K0UyrP
h4FJpgmVkj8IHeqvpw8uRkp6jozjf2cyEM38ov3kbM6kbkoQ2XyD+vnhZVrP8/Iu
SWW4z4hv70OuopRi3oOrswhWon1DulG24F7O95VCz8/nlkT05cVUivmjni89fv2p
J3JVnHNcPBvecfaqavXAmNh0JU0wAMNIRC0j878ihlxjbRHYR7lJMNCOn/hbKNu1
BOFFvbnxLcT8TqxNWFqCnR1npo6CK3t5GW53nLpZCQYGWZ6RW12DZdaHU4AWc38B
R+b87g2r0+vz1oEXmidqV8FzqYordjM08dG0DJsycyis1B3UuaHTIa6hn786N1ab
wzhYNXkCt6NFvIaQ0yIPR4YHPKpG8DRHtk2DED9EA3pdsHtC6SWHrqhsLnZaf0P6
Vpb/wAYi5MPWrS/Y6+heYVkXGxPrd3QFPlX+pVdKbaFcXvBQjLQYMZCuw7h8hcJP
UzlVHVYs52JNsfhENagx6VwNS+s8dx79CTxWo769BZKqqSGBwX09EZzm76yxjUBF
eLIdhdz2Qp+43Prv1QkYQQHmYaZkYaD1p5HrvXzqJ1AMCSh/x5EuCanR7r22JWXe
NajZWtat5d2BRNeJlIH+RX9nvs2q7RRMYWEdYpo3/SH6dtqNafblwOr1wJEApjqm
XowvbXaf20WPxDZEBwFuOpxukGLeuQTcuon3sBxibgnG3wsb2IJJ/qrqleJEY857
B0WVbihv+ulWx972Pzq703kgHAuiauDEFM/Id0Fk5f1CpVSc4tkXNqZZBZsWExsp
vrS+O6FXWSKmhwm8AAK+cz87PHe5GtFkKBDRrODGbqx2V0NOfUt8NYfqgVklWSk5
sIktZeSGFL1/15xuWcZtAdgHqVZTq8m2J14lWwS4AsukOpBYYLsszPk9evdurJ0Y
r3sZq531V8ZzOvEF9Giv65li95qeg4ijb1rJFCnbppaMhqNtdu6pnHZPe6Ba7qCo
ls0IGN+PNiDYNaE5SSI7pUJDujCwnzGP2P6288naB7aOh1AyVXJKBpLW+1Xkv96r
MV0JJO20+wxDjfSjfripi7MH5Hg0qSCcnF2uUr1B6BKth8rMYcKQnAz0em3F2MOd
6T9F9nxhGR7vXzzeDDXqsrbDLoTz1g2LWItV40q/ZOp09c3mPUM2+9AY39d+RdwJ
kgHKjCm97IePrOu9CTTqpdr6BzXxmDErXQa0dB+fUrB2cAQn/raCBwpqZdfYjouF
RY1YGFcA2f+2WTgv9HkdLc9qgQ87Jsuw//8NP4aCzEYizR/E8eysrK3KlNKdEs/b
tnj7nthxAhT1JWuV8iZdePzXS1fuMP82G34ZCDO0wQbbfIKZHgqtNZValYRNXHtB
VYPhhd2mKSekYLPLPJiwCGyoPZPA4DUxr16Tc4Yp6uL0eDCEay6nF7LR0xwywWIW
Mw3v8fKBX9YMgvTd2hcSYbfY3flX4+BbkLa5NN91cgtiWrVm0C+GIky7D1DMA/ds
fJfKc1JQFm72Ov6L3171FeE0eX1tQPZXTTH2/qGVFLESfxfSJppy9U4BlLAhg42M
O6InCuXRcSFWZPHwggu/YsIPd6bvwcvJ+O4/6ApGZaI4qSS4Nf/JVw55HqYy7/L7
jcT3DqEjCDrr/rrKm1imE/OosyVmrConO9lWwnhWljyIQFiKbRzS2zHKvBWb2/K0
qJxmKR77wCcE/NNhAqqlnBBHkiBkEgzKTActLT1oeMF++YiTMWBKzHW6UHkveHVS
fBAhb4x9qbkWY3b9a1N01psU2gX3kQJStwzHq00gG2MDHPZwUUKIcy3KkKAsL3PR
BwHYgOvKhvjhHkDr9KMTqQqhAPwfBor7JP8xtXuXd/H3hDnTE1XF5T/sxi2iI9J7
xSeGcmtVHRrF6xUXZ8dwDzYHQL+BobHzfO0m1qLZpOR3aJqO/BNWLFFLC1JczQWX
nwjqQfMgNWk4v0WNiaAjQj863w3r8V0QMbL0lvbexwng1Ij3MM/lKn3Xw0jImSUo
5bCYIA/GLVOMexNLpvX8uwskTv2Y6/U3DToxBUHmB8a7LjwGUOUGbag+vGTjbnC0
YHOCJPcY4rYn9nQloSDNoK8j0IjOvtcYktoBKrdtFr0t/yzSJMmeC7VyX71TMKiU
Qtx1Q/eNvsHzIw9rnGVUkKE3TL4/p4U8n5argTBUwaEqZXzlMqRRHKAyDhHfhLqB
/813ex5+98GengGO9eOt3PbMISuaSd7DP+Uv6YA1OHrepi8r9zqkhjis3ywj+i+f
9RUCLcemQjwSjg7NVsuIQ730j9ii0PxBsAr2ukS7gP0QvDEZF3Vdexa401z3johr
hnXJgv5P/mqB5Yr2s/0xmOnKpHAgB3u497V6Dm2XY/3Qp6P3z8QDhMSlQuVPP1QN
e/d3oUauaC2kqJkObMEhCCv8zD64gni/3QpVLYUPT27vlN8HhjEmev7hqW/jcjW7
fxIObUEU1PMW2uqqx+jODTHaQWsT8a4a098YeWQNKjEj2LiI4tMyUAhsC8tT+QT+
ubGHU3szYVG2Y5+uQT2Ck+Bd8B5gYynSK3YD8NoOXzw5iAT5WBBjXPlz+GP8zTXO
EV1AuhM7q2rLSg/Q3XQwU9Z/pbVPkRZ2LUX0HGYSp0p9OV4O1jjw8o4ZEuHx6kAQ
YFsYe8HHX7bKVIhiHPJai0VN7WXBO7gEhtbn6pHJZVtNTzweRs/SXYZx+YqV13Zm
A273s37fl+AelNil5qmdt0/0OGiATsavs/rJDHNEiMouH1jFO+tboe2BvHdS/xcE
/6A1tPQ3TNMgyj1TC6wdAjA84dQwgmhgib9fbBS6lOy/mr186B1PrQgXNe1nsWgV
A5Q7avXbSzleM9wasW8nL2yN3f0IKOVBdrMNsTKejRqsZsntsaDH3CrUff90TLg2
xuMdGWeeSIx+ASNpMVA2vQyljUuiTbJoaJEXmrzsLaWQM7Nuf9PbCT5/F4DB6TK2
2h7r9wMm4g43wvCrYxYXtomBpcJ6/K3iN221LyHeKrqGLMi/bW/6hszYESPdx/Jn
vnIaqz90/lrYpmeLX2RZjebI+Mq9/gdroypiqHvyiO+Ym3V3qSmWt8F/xGHAMkMB
857q6qkAPqNVIvmXjVD/QgjI2bzDB57QDsk9H+sXUb1NILSCovEqJSQCV+Gyu0uS
cSnc6BNqr4+gDJ6NRsxq1byT9SJdimVDaMJsH8iO1mBcBvENb4qBRm+KQEsE62GM
8YBo09Mld+8jhdJ8N43KWu+LVJyUZXWrA5L8IILGKXxqvXz6DI8R6gPERqfWlSKx
J1rr/Ze8S7GBoKGAlr03hYw7OtsMxK0dpR2vlL0t2bAgYZiOMzrwRMZOJlc9QIIf
eitEMu0eMeyxBvQTFejEZbPOYzfR4LGPGQZRUOIFT+LDjPUy++4ESzoU6rRWPs+V
aH8x/6essu62O0BnCgjWWe5PDCYIiitA1nGXYxi6ZQq1QAjbVcXFEoQRNu1+VgSh
X5aKOj/MosUOBMBApK/TGeS3BDEdslOeeTv/upiRC+FhYCxZcENv0gJnvNFAW3Ue
SFrU4pQRCqTmLMwMW3eqbHT10HJptWl39VDrGdztP8m6CKs27kUtLF71q5X+65Pv
+ZLlGIx3eZeVDu6rmwWxDbP3Ssw4XwgV7W9ktJWm0hanRYIV507sEzy7zfdJ9m9l
SAN6HpMAj7+Fxb5RsDUh7ciYBE5giWS4WVahRLDAtv3pyfRXg1bc+gJ3oar4q0al
gsV+nZneE1hLKeGf4yjBzMJda+gcjm/HdSt4w2N1J5r7RluqCn4Zgaw7C1fyIpJJ
1Fj7N4Ah5qrWcBNiClRd3166u4PGhN1gxSpCiDywQYpuvJTYhtmiJNuE+FArgLgU
rr4NwgARUdTUFFRWN65bn6SeGTC5Q44yqA/otGDMVDiDP7JHUB3YBlwfWJkjtulh
fSsiXXwc8BxHKuGSZAw7WUIG9fJruDGqT/s9bVKAGRSz5UqLnkK+Ak+8WEKwOGWM
nZUU0ckqiAxReJ6e6uncZ5hCRKRHXKqe9R2kdVqgVonqrbhP7ItjWR9Jf8UzjThh
hg4S+5yluTLuJMyChNxq5AVjIs6GxPpGKXActVGGH2JoMGcfr6um8OPE4+uD9dBk
qXuxAGKd2VxzNUfjiv3kpbR6eTuERYCOIS3KcFUANjkChCmS1I27UtacaJ0Gy0qe
QGTmkQNnDm+jAr7V2HgzWhBI5ButpAdFePTgGavALbfYIzv7pddd5ML245i6lZvL
EUE87+nvAKOjKbLl28qIOQ8d/JTNILthAffp2qRAAMkD9W6aaI/BsoUQWFln1xBz
NUjFTPap0nFwM3861pSTiWNRw9Kcke5wr3S/DgB35SB6/OxBEADiWOYt1aCIGpta
uak65hypuBkvkxtwEPKKQEzIx6wF70X7c0wbBORGK9a5MolbhUVLjoOLRK80aTSF
9at49KPRirHwUz+Gc/Ppci4C1hHKv37i3SoAVzAaAgbdAIHpdU81veUzQ3XJkH9L
nV97WY2YYQJe8HiBNnTBrlzhfoBM1hfuK/3ErOF9hVUalLqHvYWPnLEgAlMMEDyW
FwDGkR4s+QRN0BnKaUDJs7n1h9yWhwd0ukSW7pyzJHAiQKu7pmPM/jxkw0GayjfE
feM6RiwEwyvTdGFMadppbHszXllX0ZgxzQg9IrZc4rhXfrrV7ja6s7YBDs34sJlN
jBr2pywuUYb3yvwAHX3Vt8tD0Syv4R5tkz30J5E0bzaeikD0yFDOpjV72R9YKEAk
TxY/bBdcTODQ5eyMZMVx7o59J/0/834CEzGMaaX6JdzBUohkU9k2orkWshQAyzid
hB1Wnu7QlWBVKS9O8nytpclvdLgE20oKK+Ztyj9t2EJF+TV87snkk8c6YrmmzBsl
xEiSqwA+hrsglWwJfsob8LBfAzbKlylpQNOE/UTG34g7kVmtm3cdKLHf7VWmypSt
TK9eXnqhZAlr+t1IEYeavQoZ1KgK3ROxnNXSbh3k8xrbzJGCw9NUvMJ0dumiTbwj
nDEb8tgXEIaFffBCW8cfCDaxM6jUdMEj79v6UiCwH/zuoaUbcxwc+cswxNQ0ndm+
QyZ99iSVSp/10XBlZWkwhywzxMh6/nrGphE5Q5nact7furqWSR8x61o0dJPqiGJG
SPZudZY1sg7J3KVTCwFgN/9VxpJGUuunlP64MUY4GA0dIrasLgyo03nWVox+Edrv
BexOgAC96hBdNNkqkR3ozcla5sSywup7KZhxFWIMNRZgSNDBPBNbzIeee5YonvNY
bA/QKZGj1Qr+Tt/wQAezUj6/F9YQYJO37pDvaiWoNzRhJodz2JuLX7Bfn0PcA6RI
5B06D79L1Jk7hrNtqILXZrbsP4xRhRugHRip1/Np3Tv0YWWf4UgqFjUd257mTqvu
NCY/iTjrj8HjEEZ0OuOT+txjLYGTAxdOiOGl7eNlPRmWaq5Zgy25dRiQoyYYFx9H
lpUqnRBVo62u3jRCXBa8KRPIMMP4X+UEwLHo2nbC5wopCAq+Numdy4KKo1ZG2lOP
7wwR7eTbubovG0N+iABn/og4UAF/zI/mLQql6lCdsT4yRNX4LwSuJ59X4CM0zRmd
lcBGdYilAa6UNFiThRu3rX5tFu9ynS3DrBBd/PnWIjcJnA0jCkq8m5gMpznuczVR
w1qYbP+wYuTq98ppwf8e9jzCI97y5PYO2txWceiUHACwEm5SZet1WvYn+zQ04NwX
SOk2/9RkU6T1RddEOVr3t7wCeT7GNNEwdN14TCwyVDsmRGl1TPBgX3fwKvwHDRYy
0uui6UcO2EbXojeoKCPve5ElGVAOSCxqBOnvI0vtbJOTnBUPKXeXVpW1Qht9IEwm
qsBUirZoUF1ToseVviUmHnBhVbYKqsnwo3hmTFQk037yZr0jOd9OdgJLf9ISPClJ
LpCaC7YgLqsroV/jI+hHaLY6PIZzknsXP9TX3It/cmvDPjzJjMJ84sedjfPsjwVE
f5a9P5jfE1ml0REVZ6b7KEJEvLyHNqolNPE4C6br3ciljS5L60n2e1YERFYEZKmb
gPK8tqFyB6jjbdhbX5f2lR5AekzYO+ECQo/LUaHwgi0s98MjtRHIZ8p8EWnQDX2e
IJ0Hn6+e+7H7etHNRKtTlhhBr3XL6xt9CUhsjHY6QJO42FyGWUOBu5O87Yi/A8Ix
uH3/v/rDEwxMY+aun05EupchWhur0tNDKXEfVVo1ENPvfmlIt064lJxaVHPLoekz
t+PtAGzhUlY7bn6oMDj4za4/AjE5d77kl5B6oX+iGSFXb791NpMDqVfMA5/j+Wko
YE3LqZQ4H7sBfle9FVC1CPQ4akKONCjouJ5Nq1Ez/JYkOguzxb99BkfWdClKf0kf
HH1YFB2AwltXm1B1EqTGzNRwKlb3LPjlHtgGTrJSj6Ck3EZEdVU966g4BpYjL7pz
ngSXn3J3N/EA1hvDONM5jCSNGgIU18if+Wc8FyqHtz3cz9djInJuis4QJtqtfJHr
7IaMg739X/KiPhD1j5WHhDcDvJ3Hj5zQZPKJlsGASoC1AfU798/3IBNygaa+8hLL
PEM8Hwi2//JsEHXtmKqXBu2tVUmPDfC9xmltfxiGVPBY9dyC+LrPXVb2TShNplJX
m0/mWD9pr2JOLzUw82OpIlwp78DPq7ry7aaKPJbBs+1p/D98Ag1QqFHBsx8VejDe
9684uAjXgdg8LSSZrlKv1t91f+5zhCvqmWVn6tXI/h8i8UoIS6cGc0hHFhWabe5q
46+rmTuZuryRqbqcBerpa67jpigaw5C8Ccr8BX5VH3750PZuDpAA/A5BUC29ZDrB
D8X+davbMIkDhVk+1nKvmDJgYJ9cJwf8WOZ68zJL7aXdB/d3ATFkXVeAHKG7hlWv
72SAIOPfbyNILGEwSig1HFiOnZkJXyPO4k6X2TxW5LmBb4pNZ3qWcyxSrcm0XcTB
YkcSF7p8GBPTMUr/rOWTyg2GDZgivNzdGhqDRdn/ZEUutjfey2+yUKLvJsD9mDDO
kTAq1NlV0xr2UJWbNpFalBPLIL6Ohc6EIqUUJLIR60vSqQuz7I+uLQ8Z8tXvbpln
R8jVb7luQteXM5mT6zDdjWSy4TVI8M6/2DXMMvfHa9VlyAq8aYIEWvylrLFWZfkw
+agrkmvQM9oD5sV2Ef8yCDaotzpTPTyi7pLTDdc+Deis3VTJWg2jLxnt4/F8X9p1
EHvOzZFKZz8AkQnyw08m18osMGS0Yb7m68Fc6GfAIZkPNkw9TFJjl+0LDoCgxLbY
q05U2Hvjx5bRcjSMvME5CM0G8xQnQwOMciwigH0R1gypLYddaMANVvUSe0tncpO/
sS+rO6aZoFzaHxWIK6IcJIgWEUXTwF1jdjlk1l31r48zw7Ic4Q1qLhueMFgUHowr
VMtKlE9FVmoMewzVNwsoZPH/KHQHmoXtnfd9cTWHAhg29V8AvQ7RmT6N40CFWFg9
mMzHqgMWs0fhMxsv+0wgH/YdJ42tvl0hEa2QbXHWZ03Tn+LulajViiMaQm2YTNRp
9/qN1yMICm6jwN4TOJCsZFq2VuhaNI7cCbKGOL9wJPfpWD4VzfqrWYeKmSY9oRu4
M465LI06yuXV/fTNEwJU9SN1UG7XIPmcKa6lrPe6vR18lEF5PwOicNpYUZ2B+J83
36iaZBy0CR68BEzEnImOmNM8KFhR9vPKuJpDw/xqdr47f7HgL+ghd5qzmbO6OU6m
Kuo7SW1rr+NtqBJrSY+lARSy0xS8AGZvaBiNCQvd9bIB2P+YYjkEu8OKRgAe8RpA
5a7e7ST/6EcAEga/DG31WFpaa/80mfg47DWTYNyp3x4bkXxVxISRnULNJuZRt86T
Ky5EtsSjclvXGgtrcau/YVYtKEUWI+qKQHTkJsBnyXu71N9SDTenIw6iuCBnEico
IPsLGpLnduDIRzSmYjsVxFPKhxTI0woNJmeQ2hfH5Xx4xXnKSIOqevT8WbDlJV2/
Cg3Kp0/Jv04SaW1vm+PXRH+YcBsCKr/+vNDTvIMZt5sXWz81+xq4v98EjutLrGfe
B9wcNVUhY09vZAsD9E7kE3HB5q2hx4TTRtlhdama3IAuwKwjLYUUxKpTec4EjUwb
LjOP3tIMnW5nCcfXE3TC6nNA6DBq+E1O10MogvynO2dmkDZh5iGp/7o8DFdNfbmi
9d3Rxyk3f8zbGwc6zdNxONSk3MZgh+il48dqJ3GMnbglI/Dy+vTZ4dU3tJOpHP+p
Ia2c3yPtKRM+XCsZDS7Pv1rxL+iAF6btRclQBuTlnJoWo04OXgnBvJaDvNXvs9cE
iPSlYmDBUTb3jvjNAWvXnjjxIwUeBk0350TMaUvPYmOceJsftI+wyHnaAZ7cCQge
cz91rR5qsNf7uIpLkhOHzlxiJf9QITwwupXsvaWsuaVpECVJj/Odya6TS5QWjeFq
Udknw7KtLyksT64Q7xjQVpTkIQro5o/7XmNgGAXz8A33PmOUx9Xz/H2rLicw6MwO
sT/uMRlpnGNhUQKueNUHLKgpOjtCDvt6Euh9xXPPenkVYEECwfN1nqIfRU0aLct3
fvHxfMXbc4oIlBQ9cYsOsPsOgCWwbGa2EiPv26zeLGkcX+xsLRWQqPMj7aY0E4qD
lT1kO8CtdoFkWxMNFXr2kGIAiLztUuxkojbcU5w6uR1RZgjKfeOig4MwNT/kWrGM
H+zLVZgohcoxRMrdtLAcd/3xAelQURNBgYnwtLFmdFPS3YU8OlNDRsaCDkcTXjVk
mUUeAit3oO1QOq7/BWHQl+f5d2jw7//q6Ywub13jVwIFiXboxlXlFayaJrMNcaw4
K6OkHr/NzILHJOlTiW3s7ShFz/Iu9fQngwAdNhZOPrC/0+jAJwidxbd9pYGMgsib
B3CiFJVbV6G6pAEVkZquCRoUcXHiigrSMziJgTRjbznlFqwswsTvRC5f/1kCYZbm
PzPhkXyLcx+xRpO2ReCMH75xokT7zfIjGgnj25165cNzGkXTmslwTQ5acpB8fu8L
mKWteGDMlXtn2xMELKOdiwM8koZIiBU8XytdjgZa2/uY1T2vIOKPw1m8xRsfXkIm
QHC4OWVz0Lix8fVAGPamAiE4//Q5TEAD5Ex0JQ2F74OkWowFGAZYVNwSZvlNat+V
uIopuue6+B3SobG3koNglge2B+Isj5F16Q308s2mwnBcTPv0x6CGBdq9vrzTUwB5
e45nbRixfch02P6469nqwyOVTzlEowuccc/lzuGkrGDbf2Tp5Lfz52FoyxmiUuG4
KP45RipcPaTF2KfAyzjklHYPzoZVxcyEG1WbXIAZhFbmqxIfw8INxbQQygfiVt8v
m4QMpoj6puT2YFJ4QvwAyPGUMcmNg8bjL2NkiPAjV2d2avXVZw9adn3FSHVIv7T3
vcwlu1c1u2ptqMiwYyUPOi8OSSgsECuf4eON/qMu4bX7ndSIhM5LAvQnkncdb34Q
vzLdU+4a4DILnvWVXiXk+VNymUEPqWjv1YwSv3GuzXdRhkIfFrH+W+cDq28pExtA
OoPW1DNfX4pIUz42pe8/93v2dC2M1wa4NWYh0jcjPF1iZcXHlyjG26Qw2IMV0x77
I280AJui4a0BNXsuyuXRFyt1CzZidAhR9qrAzd14ucnBIJD7zlMrZd5R75BzYnhS
EuMEJCuxgU42SBRgJoUOt4acI9VieRLFmngPs0WgKnAMNzZe/KCU9o9r9FkRuGfx
8IhuDrv7YWmPUVgGooQgOoKbLclzL6oYeJu7b3aVR0i0msKJP+btF9deApQbsl5l
4iqQpd1fpDErT92b8F9pP9jiiyl2eMrFTO8kjX3scMPr0PfS/sh72qMmqq0inwcx
6Mq5Gb77mhTUgi69AGnmMJJgm6grsXhFkerIGmN0HBlu7kAc9Rx57bkiYDqi7Krk
skGUrTH5d0xqg3kNJDZE0MgLUCbVcbwjMeqsaMu1XXGPBUjObtLG57So0fgUF3Hb
jQ5sp1BgAeorr1VJVvOqfgPZs/n8sSTaZ8tm190psjsaRdTzWLQ6vzDbbfP0QG3n
fsXWzJ8yYtA5UlJ2b7AoAp93Kf14GR9aYIWwtxPwJuMmYFrtaOGpXOP5o4TKF/P8
jOoNtEw4or0ix064qtpmEjx8zERo/7C5i1b691VTwcpxuHccNqvoAxdALLyGsaw3
b0Zto67lUqYj5KvQaC756GGNim5wCAAHzm9N6c/jEnqdwhHos8YERkq2pdbsfvlY
v/pu++RXpTKyq4unuclMRa87cKaioKM9cKlOqZpZmxj+dxIEfvHJ4vlF7xcE93S+
Ja2yhxtyxQ5dgbxHmbA/m0rdfZ1J+z7fp5EeNjFqcy2hdhCFjV/Oqfm/Bm8utKi5
3QLjIBd0uHtiPM0hDpy4mB+ICyQYH/vgVE1XTTyKpwHzFZKfG5HICkUGMq72+2bO
9TKWqdZKTDXTABD2ehh4i2LqPL3D+nZ8jqMozQhbRhVQNjca4lltrYOJ5MR6tFwE
OEkRPuhbzo1pdduvlO9WcKw8TwoZo8wZXjf2YCmUMv9ilHXhnbMQqAfAqU31IwJB
DvAp09nMYzBR0uxZTCx1Yzc5IdyMZNnb0r3Ln1ktRxsI5g/5SKmVMGKf3JJcUpbK
1Gw+ceg+W6xas9CrrQwYkK8M+6ZS9n8+TB45dM9SCmnPXuhRzyCxfHapkfNNCxsO
CcfI0Jd8hTpv6pSj0QAw7sUoxBkeyY+z2jdF4kRoite73s9Ai1Zu/MX4Zu4yNdpY
tG8hScjValQVzfW28glhkPAtOyZL6OSsWphSRTkssjBhs3sRtIFrTp6HCpkJUbtW
YfwVakGT1mxJIWQJ1bplqtI+ZO+3ClSQpU4hd4cDPPUmczjPEY0Lw9xo2KFW/LoH
p2LnV4wixkv8WYldM7VGOLT/FTvkdm2K/JC73Q757cvlC8SGTqgY07PUvNewsXcX
iK7ScDI0FEEO/CBHzpCVD9t8odD7bXMIv7UXI8+hrqCO3VHkPkQ7YDHWeCxCWCHL
6S5qyRVQMCEXWMGPAMQ4DePQmlar2imdmcgT0wI0iUFA3ctmrU3rZxsuyfSbd0wO
SyPP6LW97SgZmz2GYta5FLYeMs4hxfqCfcUuCs4m2yefwUD/5AVtU5SgqMlvWlS1
NK4/zeFE/qLH/2tjHTe3Q+CnG4jYYJZgTUVoavsNVV5k2lzQsPg5qmIfRJwYuzs8
wIpZ0AMQO9ASlnFLT76OwRS1bk7QzEPKsHd3TgjvcHytsMQCD3HrqLughMPvyxMk
jnHVOq+OrklbVBWoqH113JcGIogQqOS5v9b2QiUSWtkKdo5Sm0h0vj0+JQzytPO7
ikjGkUgnz4vdRvePHF+J3h95T1KGFkwdsAUwDpFyauFSS0+82EMPtu7kQ+a99jPm
iuSIuUx5CtTdNPbrZ42+k3sOjvmVBUobfTcnO96Roc6RtaHHVm7YJhFwMeWCV4m0
NmbI5elg6NBF9t0JvJa6qrLLMZj12o/rB7V9Fq9rb/CCOFT6/O/QLMPCX8PhjAis
vHj3JNvKg2hUND0eu+M1et0GS+962rw75+Vr/Bm8250gZWBFdUB6ErY30Newf73V
540/aDCanfyIsqexYICdB0u+Y9lGqqtbedncu1U2fg2hIidH1BT5gyZIlR0b92Yy
YAnWLmxBNCn336wWw+O+ntpn/zwtF29l5Z8JQxDd2JEq8nB42I2vgkssje+jdItr
FGW+CWeEBkxt/U78SLgsUxYjnUkPmKWCSRJvF40Ds5JydLkoCormu4U2ylPmqBsz
/E4Q2hDs+V47k2hvci1xIyaMgrnXT3b91mtJQvamNQ82THXdIbLXdbyhPOyWrjEC
OHRyjvdk4KAqsoqEmC/7gaj4GGnPZXppGS/XkIRmaYuUnNUE72hcfZ3nNlXVjLvN
n9KtrTKl2RLeQ/YaNrJBVV1uO+egz5LiYIJhpn7EaOMnEwkr/OHhGLVsdHWVHbAJ
kQF18gUl098nD6d/wJH6tllpvbp1x3SAjEYg3rTXBZAMLRt0pL8csP4dpPTNmILL
QCIgWunVzZ4IEqecMPQRvftzQrdiF3lMSepRWPnMFrj+rAzfy+rmon5CWVrOX4OC
cjyTw/GjAtFBlliRqohUSSLA62Na403B8qB9c6kvl9gcg1/oZCtr4b2CVSXIpiV6
tHezTGdZ7BioN9Ykxd47qTAo6BUXT35vm/xZR8Z69oBNYEikmoS9BpqQ7cSE1RqA
9x+I2PP1w012zN4RHxMgaaHkpKeeD/okzSsuIl4HdCNRvqxNsr7C3RFtN761OHKt
+snA+EGAZP0MafGH7iVqyjqByJgJDSN7w+GdLEahVWNEYjTzC9+/aCKszxM/CNv8
DP+gkdsy3zBRBsDcKRnuqRzxeORlCF/GvrnqaSUpSJ6Z680vN4xSyEMsJXOiswB1
0rsmJa+a/Y9yN1Z5Ual/MEo1XGoJ8B2AXrhDjroOcDW5aWUnDXEHRHGEi8CDlkqj
OOzeWL6LhyGRftE4Q5zhEkbzT6l+ZWd4ct97mxqs1S/sv+2hbhLqNDOoK/rdMsUS
R6Q5bwmBZkiEeJ7MXeiKiuttDo1RarvnW0KZs4F9kDg8vzZzbS8lroQROHNLHqyX
W6JkiOlBbfKilYXgoNwpgxBj9mwwuV0nsoYEvOK44G9+SYZfBGYo8YKsY65oa4Ly
oghclFKltNjkDL0cxfhIrt1IzH5BZQXP1px9CdURxQDjLV1c6B5v2m8v91xzRpmk
2N/SZshiDT3qIFlBgdi9+DANlPVE29PZ80ldHc//oST5WMLdj1NicbnJkEo9hyBZ
P7a7fTkWMj/1rfbNmPSw0y4+S/SKayXOkmjZZZbM0G5rA8SoTuzkDp5GRRSgVYpX
4biQlnCdy/qlGWNVKnMwar2V82CFej3oX8/OnYBNu8g3/C6+bb58BoALht5RySCI
rEYl2K7JnLYRR3p04OEqcaztXfoJHOKscYUG/qF5gBD2InXKHYKpeBs0EuaDG33r
SMMaYXwnRxAgVvpcAwW7W8Pa8krp8gfBQByF2YOusDLDz5scThZSgJrllWm7aKPK
miJAKieZeWsVd85xLdcnoXZA0JBh40m37csJbMlDiPjSmQC3mcu1MyfROCuFZ88M
kqGfvXVW2fiaV85mxLvOBmX8/BIqVlO/io6L7ZcMP1mKLMK/ll1iN6UqTjghXFyo
2z/f166jICNLRso8gdaCcbl3yOI3jZMRBoZgOuSSGCfFTaYd5N8Wis25+mMKGj9K
kkSVtP/LLh+E0qcH/F+L3e7+BSFfA3l/BVcnK+Qo6DjC18fymTXjKJidMks7IJfz
uuUCCe35OOXaxWlnC8u0YdbpsJF1lZ0ADX0xKBW+fa4qIoXWDCEoPTQW7WB/EgIf
EbEFGvol0TWWvW57bJuWXVmtIEkLvorM6+hcE7yXraNk7tXtQ29B8U8GMW4xJGWF
OsyaYKnVme13OmLW4IQEyYyeF9qczbeLX0JtiYO4kVEy8d4P4n9PAja2S6/g/ID4
437zsuS2W0FOknZQ7fKRfo02v/trx4Y50FyZe9zCnLOu46QFTr//MhDNVaNZYKBo
D+cQ4SpGvH4I2n6TJOxDpzssqc4olitPzVnA9V6rYmrbiOyB4r8+CvgzXFkQdvnT
dZa8UHVxV02CEQco5ovLYn9mRAadeu5k0NKNJPLWJMqNwjBpQ/U8ySWz4CCxIOeb
F3vX4gYp/cOhfMW5gXscwIB79pEkeqRXEatOj7krOPxmKjn3Uy5gCXUvmskHBgTC
Hv9knXilyg8Z+zINFZZJMep5T6v9iXwId7iGihMTIj7wOn41M1UXLpMClkJ1ZeGk
5/6EkOqOQT8dmibGWo2bGJzg/7HX9nT2kD5GPE9xA7B1VqIEpltiL9/rApHhh6qI
+6SM8Pte/zHb/2x1dUrNzMCqM/cqzuatEHPwlws4qbXiggnd4HUCA5NkIIksvHSC
KL1lHy2LhLWG3868riPYn8OiAiPK1MkPZgu/ADhFD4wn/tKYzpuxnIsk+SXjShNl
R6pju3zJbwzRHFYoHsfZ25MeyCSbCVF5SBq0hT0IYnu9mhTcHZWqYzEnc5Kn6FQH
6BIpK95SnCorWlxlYmLYOQqLjVrn6ir2RxEK5ndg+BiQZ+ExHQVIYFCK6GnZyAge
CLnvUj7nRO3+sVkhHqa2UOeLLb+uGH617A6qU48TrSdWIzhj9/8n+2HI5IcJIXRk
FikbM+uKXBe4Z3DdXYhvbi3s3WEURAAq0zxhbgc3GPqES6c8C7YHF79ad2CwlMs7
Z/LHCyhovoyYPLmYdkbIPUmWFNn/02JWgSeC9BIW9+HYZhO4FsBgybnY05mifzzs
F54Ahz4+8SvnytgTvpKX5rZnbi0eC+DdiG8lUqF1PVB9ZJMaE1ZT3SqEgHIP6bYK
MVHfqfFfxAIW0L6lPntddhOwdmC7by8bV+oohMhh6rH99INvx+0HzcckGQzpUPE9
zWSjbeJ5DBOhrx9MYZ6ZaSr1k7kvsdfcyQnaL7BEVAOFjX73X2DyunZarfkLzAGp
Og6KNgBsQWiBF/HE3z66Uq+AWn1A6Jiorq/bFkPWFCdTyh5LuHovEsAetl8nO6gf
5GgOkpJyhtzw3qVCmsTFOe1YVGGGD/DUZUe+xD8CYVh7fzCLjsD68E35d6JvUdfB
W9tsqkHguXwJ7WtAbjWuPgLtTTmLttO7N0lsNCi7R4UbfXlLxcyGa5MBg63QLRT2
8+mYBxTge53iLSZmRTd579+3apP0zKqGu6wDEsyWRzRB+9FkfgvVP2XF4pR/oHNU
0XTyFlV5XD0xzuINYDBnKcw9SYGnPWkWe+Mhwv3BbNpbHaNzm/ySEHjKDvk2zqfo
2BDBpUpSc9s8DtOuyGxZ6e9ezDqMQ2oHw+dT313t+l7It7EvCa7BqTi4wrD022+o
R3n32jQYN3OgznrhilANElezjX2u6p23fNDwBrqLrBO++fCsLPgwb0vS5cGmVPwE
ff+w2WykbHF6uGwhy3BZ3H0j4nf7g1hSxAFNMZO70Vo+oYW5/lZ3ZCitNVKUeW9t
4qD8QyZjrTkKlTuhgNmz6okkbUa79cOk/mkei6+Rg108ZEiAABD7aPwdsXCk1owo
SXZ9ZEq5sb7113RFLo5UvCMKZ8HEA5ZINCRdGspf4djzdhfixDvWzpbzAbQ71v2d
OHviMo3c8gBeYQlJV6TdC2HZVCzam3UDoRYYR6Ta0ar1llaLQWz9HOmE1ipLiRc7
YeXBpimP3KKXDONltGlig8NMRncTVbz5hMLIRvHaqyBShD6qF8Zp/A2ggllZN2sB
bB1nB1QBEdAexxdSDgPhHoXQEeoUfZElxJ8g0Vbu7EN+LEMmYHbSh1+ByMg8IsC7
7b88D3k1la8RKoycROE8yK/59CSnYqX8tOjhvz0W1QDlG7ALS//RYWgcUFSSmX3M
GZN3TjTXjhCcbwYB5gS+zWEhBE+g/gXxPhRGmvFyS0vlCWcsRSgM990nTnPmrA+5
Z5LMubCI1jwLVguc2akvxH4SCD5B64nbwGmCOkSUTkKX+F4Tgvi6Riu6B+1C8qJx
7T8U/mIC8O6FTZwA0KskGK9cTL5a3sEb7KY+tjzoqcgRp1mcXsOKHuJcXArsSH7u
eWVMfRVoUCNbZkDqj4Zd3LwgqFZm70u5PKkF35DoXdbW4geX7fjrcrEY6lBbgTRl
3r+LYArcs4oq9r0TASdHqk5ez1IQHn3fHin1vU679BPBdHOpUX+3UsRHCYZ83Uzs
RvN4chHV+iDXaPEWFTV6aRGjFakyo4fMXptsvbV5QAoDuXjS0S1o06ujNusCd+IU
8WV4YSwJdfoCn1gfFQaanBo7iIulQdTBuAUgxx+WK/Df0X/Oz39EGw6ccGwEitYK
9HSf42QxkQPNHei8OuiWzE2ZdA+ixXh+fctIwEO2wmd83g1M/JFq6SSDeGn77urX
+wmJdTERxuIX5EYUVgf7eEuSv35WHB8gsQ7jyP705Uc56YGDq+gGq9KrcHczl4mm
pjIEqKPds8JrURU6xXROtI0Uu5UNmjWLTI0FRLlFVEAbDBEAb+GF9tsuFoJbVHLN
tPa64R/QH1Iel7AM1sO9icqK9xYqVWzsOmqV6cvKnJwCYNq4rJsJm8nwqBf9JqfU
NFJ6OjaU9OFJxLivqPzJkg5cVN8VwwM9ifU3UZKVNsnchSPU9h7/5/Yj3c1WIj8R
3YU9Hu2Wj9s0egXwPkWNlmRBIYypTLe1lIXMhAAodptf2vCYPsOmqyjtttdJc0e1
zbe884PuPJm+RhJTxy0AxBkyOHxpcIPAbsKGpQCH2pLun/ry+IpeO+oY9fLwXqZ/
vsDfmMjNl4rzgaJH8Fxz8M86DOSIoE17pOyJv2h10V0XanLjrMBDdTF76TnN20P2
VlbYSQlfor4UsWBlFyfQpo4XJ9hP8LmVFG6UiE4Rzf4IFIcqbFZK3Ey0d0o5vxXj
YRmeJS2YNb/ZvgxhXtabMOaP/s7Ri/u0H2X3yIOGwQgtK9qiS8EaW49FG9kUkx28
seL2WWkjMuBpgr7xD571rW8mO79RSSCDCWmrew7ZQAapqu63P815xEIDspS29YtP
zu8NE91UW9RClYAxCFLJ0DD2WAbho+7ZnPD0eruG2AoCaYQk7NahWGka2cF2JUfo
R3A1XIHyFUF9FZ6GmnMKmMvuI4UjtxZHTDF8nQtTIPzdxi6Uo0sRiPqBD2QlkhFb
Yke2YwXyjQzG+nHkfAKVrIGlYpHASPgPuouoXbmoQ+6qK9pRPHxSfgglmmr/fWma
+sjwaWaw1WCo4R+aRTOmUOJdF6dp55yXKiyX3J2mRW0vdRenAa67bFjpWRI0OfhV
15634NpM4ht2HpPfgZL38MFDO4dprD/eTGubGP9O88HXOIEcQmp6a5oIn5YXI2bX
acNUC3SYw293VLxrV7a0uPMZr2JfOcmgVJTbOa20Puc1x4fJUPpkTsxUD5urPxTb
3AOczUkD0fnoFmB46onZvWTCCPoxrBW+eBc2GjsZxhCdXLLOUd879Kt1zY/3Z2vG
jl/SeFR3roBqqCO4sci+t5Tt6DZ2D0VKBDR5LfthERycJDcg6DkYkVklthAvnunz
L4hcVi/mKYvv4eCJ5wmJjUxalSgKsgylWs62IIN+0zmSOphnmtLFu7E2a1Kw8un3
x6G3ZzU15Xoc7kitqGVmIt82d+cweAr6RUCf6eMrBOgMySlC5U+jFyAcBD4Ong6I
qhUg/Ip2aEtCFkX9Vc43LTlZkUgWVS71c6RqNMMiufxV2mw85TIS/MFHQbMamhRg
+BRP3GKzBd4OkiFwAeyFs96jZv9OmY8KqboB34GRHEFyXDEQ7tqjyH7uxUaxxYc3
sQT2aLk+PSu22BswncdzkzvQo2wFEUYwRhVoe5M5TSwfToJQ0Qse+xRYeuVXy8NI
oFH7HP9mx9UnTq33UYbeN/q4iQ48I0hqHQzW070K/f5TFmmRnq/tyXYSXOEXTxm9
5xIsJigqbafGxGgmTg/E4bIreEiamq8lVz0ybif+EV4rjZFKAP3rvYyy1iEfjoqk
dZmHV7DGqfrIlpJ4mtF+nMR+1ixDLPMM7hsyv9BlERHZArao95bIXteos7TUUs89
6s4bFkNm18LY+AV/92YyL8wmY6awYMnoX7CFh4U9xY2YdvSTwXJGbr+asaIlGINw
NSHHtlYtTVJ7a7mEPmMNVc+xRranOt0xWi+CyDmnp2YMgUmreF9NO+K4/1hJ7P1l
3I1QJc2LlBqm7flsjcrKP+s81AvED3HWfL+IxwXpweO0LPHzKwKWUE7CipkKgw0R
b8TexJxVZTW9dtcXTZuR6S0sRw3lrJRzOJQZ0zytLGEDbn56WtK0he57B+BucXya
5DKVXb43zFcQJXSR0J/qVs1rrFQdiMZtzX93DwifACffFXhhGJog248WVTYQ/EzZ
doGnP/AyVLV8ao0puKOLm/wrGJzENasDBYSuuCLNxSGRI9T9JNy+UBpqb2vHqs55
X3Nn1lEaMBzxr6FVyekGnbogt9sflSOgdIRIrXyd+Yu3Vz6b4Cfk+J4fILcC7d5A
Rg6FpT4np0PwuVuiCQIEV8OdKit3kRkvWt9XyQoAzmrWg5pn8JWcWJdh9pKX5vXg
uRwGu1nVkNcw5aGHz+MxoHkyFAq92D9bccnCQ81Upt3jSC8aJL0msrswu4jBK5YW
Cvhrq7v4GBh8phlMhHGydpqNFE0bVG8dKz20GxjZC5ipTNexhTc4aLG+8mhZc2Op
Lta5thokigFYyPN6BkyA99J6w+npmLU74ql/bANaNAjdFvOmFkiZR/e/kuGLd+Ip
+6mznydyhUU8PGIK2B1L4Eug03O+jqLrYEtne6MFM9QdppQdPoxDmBWpq7Y3MRUd
XoxTnGFbMXsmB7RiwthigwKJsvTbkMc5AC3EsLVa5Hul82+6LX3Xc3ux98aVWak9
Xqm9dgUlFthdpeHJexXZnnMFQYvzgOmTg3AlgVGj26oHUp9IiCKJGmTQ8W1fekDt
Nvc+ypbURgoIu/q9wgAAGQMUn+GX4W/yOKkk91I+Q1hCs9BD024S3/L5rU2ejG5h
Xa9Tom6VuMblJp+cTRFir9bc+dg61nQUvxaP7V1jXh1ktoFzEQuBs7M3Lg9VCd4k
4V1YscVx6dWzSBIelI1VueZgyAcLjlUWSp3T3D7EhsSuHSTeo/z78sOkFTH+mPAv
vVOOCsdXXcpVFhj2ZyNYkbM8HQB3ovG/GThYB4a5EyUWufxXctJQcTg1s7CLdSyt
2C2Yr55mrf7qWTrGlWHVgapbMXPfy+qgfp6E45Nmi6dORsElXm1R96erghKZzxF+
zpjyJrH7LJWMMS20vsBGNnpDx3uUrdMImaJjElJv04RWAzDsed/wMcWJ5JigAbU6
wjywK+XCSawZseW3fhCmJSbyli0Rr7OYcpZ6vlpGrLHTwlCMJ4Ol0HdUaOfDsXK8
vsN6T7NngmgPcCkwTKh4j5+LYjUTWroC1rwtp9EY0F8yfrrmLVNKbSWLPm0q9Jl1
Uc4b+z8GE756w0HMDpUrVGSXNVK4Fxmkq5PN2IAVEM8QDQTWAWl4IYmyqvCyHTIi
f1sj+Td4kv/3F6/ooUnY5uvIkpWuBGCNKWW9NPmFEfalEscOigq/ARw5LU/D3dwo
w3pgCro5u39RN6m/ExdzXu+jEthrimnE6IimTwJ+g4IsKSqkajNeMoRA2qzuD9SL
ZSBiq64y+qKMgB82IIh36nZ9/j5gWwG2HMCtmP58+JAo0DGzhpULPz+8NGdUr3qK
lxdhUi1M8T/jUNELVIXyLvxf3nVbXAnQAwIXMWLsVTZgAwZI+Ks6yW8iKLHfPOdF
zA+kGLUUNAO/5wVxY7qF8AmYLgOgOzTBFOp3UV/XP2oGi0QoM8OuiiT7RrNidSnp
zDkZlsLOzCJIjaYfZSRl2hxgsMv+BimVk+aSDDqif3nUk+ZSFmAUgY1fMT8HRcly
dV/x5sfO54qvaYzQ7/nX3FIHUKzvI+rOEzgJmRWg35uz1qUUJHgShbEffurnC85j
MBwer8gYOTX/JVu391fby9HlNGxrs/F5HGWFy3Z20qCxZ//OdCHqapeT7No3IiJ+
cIPR5aci6vnbrzxR5Ym6+qXS+g6i/3jYdPZMA4Mzjzyg+rPaepAp6jJ4YwgGadQN
UpISRK54Cx8IwkbzpQ7PQx0yMiVJpe3le7RbMGWrARJCNknLLdjP6hmIaEG8QRM5
xQF7GX0kgKHgB1CFRoAsFKBuAHVWofWUIeSfJFYgj1WSfwxarPCM2WGuV5c/meIe
coEdB6qpaRBG4oOEfVFhtRLBpHv2I+ulpDWyNuM11k4ROKDiOoGkmIGeKaKAw83G
4+97j7/+/3eFC1mL/uz8qnSaxfQDT608mEYN1VmPP9Ef4WpQFBaSTguLwCL76QcK
odXUpADEMkDe25A6WSscgy+Bqx523weLi5A1CLBNDXOpvLaEC1FOKsvXcOhWc4fg
sLwJGh6Y678IVN7Zzl//zc+HrQfubxEicr4gw3jk7bCNXEFxbYonQX3pwTVbduXn
rz7EGnQ+ZKFOa6B8/INl3xRFlUtIuzDmdLVHUQvwh3mkx7U8Emnr6pt9LAU0s2lP
6wSgcNSW8dTcE0L9RnpSNFPv+3YKFKkAtpOmgVegvos+1mHt3pNglLqcWnwU4IO0
xaXw4t0X0l03KMPoRRA1JOG9jeZrcaBtFfouC8Ylhu6ZOmaPiieO5B8iG+XW9qvR
T2BHPhgNLW5AHzvAVhIDQdwDVXQ6nz1fs7pTxMl/b0uYLWV6ASoUJb0HaFcXkrZk
f9lfqk4yOKCSLL7h67x8iNYBDwQaIN3IwpBTq+COYjDR6HGlDLzJPZDXIYhen5U9
36Cp+vBedjC2fABWIkuQ4B6tt3d4yv3RUrEZMUEm/H+zCMDBNjJJC/mapsoLywv9
MGS4kBFL7Ykmv4fcC04Dqz35nXCUAXYgZONc3LhvkMgp1efF85CAZJScL/Redj0F
WTf6DQKmqGL7sGvrOeh3s7uCjj6E1S1lExG5Je4RhZeviN0j7gMiPsiJvAu8rQJu
kCPKcDlCMdhXxyagJz18kXnXBZ+DrSgzRjm57tkuqzGslJS24ZpeOj0nBDxK4We0
y6kiXAfFUWi2BZRN9CikBvbHfVqkEzatKfKMJB98T+bgC5M4263MkNyJ8GZUuhG2
kq45Rr0b919LbVma9Wr9PRjMtPreP0GRPW1nXhh9Urv8YCymVEmb7phjPpAxqvC/
4kv/fLuW09nDAYy5/RkEwD2Yi8Wfr+mRql0Oe6MxTXhRO0xFtUdZz3IYqoZ6C80y
IBDquIt9ZTW/r7CIM4HqV8t1+AIsJVERIzWho1rrKWI2YtsOxr5/izecizcn7vx8
xxw9wl8Gcp23GmkYM+ETmwuTEgH83ppI3oppJfimxECssP9vPZMXm14YBEp1nAuq
gXS0S2DMDUV6Df0vi6DfgUQhLw0PHs6Wo5RAIynWyTUVCQyKXW8R6KB0SIZtUSBr
/h1FOzpfdCc41MGCecntrpx4dEbu1/VaRY1r3ZbK6K9dDR70htCqxhbtn24d1vc9
if/wDORARzqCpn+ZTHbUPkqAmXXyJKU/WPoB8BedQQzP7DcgmhuaPi2hCJSi9xkV
29lYhANaNco6lHRh01y96bOGb2o6fKha9Lb/Q9/ZsFGzwkQGK275vJkwiT9noztc
3biScSLiAUZHWKWRyDJg/Rh3cr2/fWdbBNiHOiNpZH3HXIJeWBRZW7ZxzGcJu7+E
5FSzqp2w+isEK2NVzXvTy9jqu55U/wKX3Wfgcn1P7O5i//IT1yyaC4lK7tbcu3S0
TzEtS4MkxWcHbyxcXGnsjqv6iOWqJKnyWMQAUEpA1jRGPyXn/YISBZMXusRBCdlC
8Ilkc1i/c4Ap9GmJfSr/bz6t9aEP2i5PhSHL7uTxfedDRw5LfTuxzTgysjtTalrj
w7urf91rGYvkfnep3Wmah5t7On3KtuOh8RPob9IsiPHgAgQSp3dOHOjOr0bAzNKY
oV4vRPBjC3szX864tuU4K5S52LXA1hFGs+kYw6wGxYxSZHrDXGEj6TCGw+sa8kSY
LVtdsWE6fPkz0aNfIGKP23UF5CSDqnC9c9eDBhzb4iNVLB8J/2qLUplyHOM4x8iQ
PClhX8vFqNYLQG9bUKh0bzXt+FgP2JoMOuwdc3uZvrBz8OPhgQXnWvdD4Mn9DxJp
RXH9MkZ/LAiAwLEwuS7HUdrYYCqcoWCzPE7OwWbLO/vA4xjMgkp3Yh2xXYcWUnuL
UK40e1+OD52zV7bkUg+VUOAj0j3bv8rpImjnSEoJsE+Pd7IE+p7guFq9lgBPfxQm
3cYx4/rf4CRl2CVu8mhmKLiD2Tu9Z22hVPpORK/bBv0PGDfHbegEpWqM7F2gUL7t
UtvHLnSPmERSCdCcLJ8SIci07AGsYaVJJjq8m1goHr7d4B3fMOenDBgkAhgNpilh
T7LsOrBOijE0Yrrc6igvqhXMsapdybs8bGgmso+MDe9QoqJFgDzvyZFIp1GiwB3w
Diz5xhxvyoIQeK53Q1zguTuMHiIuIktsAr1ErkLG7gf0kYs8ItTjvp4jAmK0d9OA
UEh5xO+Yrsp98eoIZ6/jFYMxP5vbGqRl923rnZWZfMxTp3YCjGc3yB5Vtog51TGY
G7Sqeg1eqsBGsXJEQGYrFRTthhhjSJTWL+zfy/pY9p2Vebyj6GnJhtlEmGOlwgEc
mbdsywdBayzu5fs121cPMsVSXuuc4iOBGyCTjz14PZJL5Aj5LTdel4NKHYPujH8K
zVV3+GDeVKFndToL0lCSM4GSy6b3qUylyOx4hHT+oHGoPY4/4o/Kf5vb4L8AsxYJ
yPxuUr0ser3vSgLZ1OgiGm3QuZ2cZixqjMow7dc8H0AAxIK6RgXXlS8YvysL4jHA
E4vursCnDCZbJ1ETDPImu1szf6bQo61j9vNlz28uBUUnb8O1CDRsk+GP9UKJc9r3
aq4F2h0rgbTPdPdaSRf3v5+wfHwC2puKCIzDhL4JiHY812Xps3WnYgATRi9aZfHp
gqCWJVN1WVan1ztcsZpeCX78dRsRUL2+Jq1PHnHvuJm+4x/Vp9fNOC57MOB52TOa
Zd/dNk88NZB8KUIMGjxKpHILiUKlt5isj1t2znaOTNJo13Ttpbf4kfn6mgbDYkjv
U9Flg2D6f2g7/IaV13zSBeap6PJfg6yF+jkP7/iRKo3Vx0ii64WtQ0Gnl8gEscer
pm/XUfiAlKbQKN0gDJB2RsWuqtFsR3mVpYw4QYXzmdhTliCtpPryVeFtrsRD3+J1
3JabBIncQvUisc5dXPMbXPgUA0H8YTmoa21oJmAljZkf/a8s4lVqHXDVT1l/LyK1
sgePxdhqoD+oe8xv9ZSxFNL2D9j60fF5rpqJHzF/2nr7FFYS0EechZdJLd7dXgVw
u8b4F+qbGGPkKbSsi1mLO0b8mzs+YRGRGGnF13oEe/Gckdt+6wwIC8wiIw+DL07c
vNI42zGxQxjDxhyJXhtm1V2BgVmPn3FXhbt2uWvUOotka2xFpwRMa2JujAYVX/G7
hg6zdHVnhqc/R4oGITNUxMyMnkFir5Ef53VUOzHcnWOSYPwZf7tw6dVi/6Kkb9W3
g8Lvyn8iOcDVU4cf9rE+u7WEVNNRzOn7CwClMRwcBJPSHfgloWRLItMsyhLFygJv
n3d3CgIoOX7f8CcciXmx0dfnLZebyRl9dBra19HIgoCWsqSwJgizwkAZYQQ6GqNw
lz2gM2fWiTjftzMrexT2x4ZviOCDnHkzYMCHVsxIRVn85njZqa42of+AbPIwm2ga
Y2DX2uS68eRBl9KAueNUi+VWcslGZx/WJQqifWDA935jX5V4hXY0BRMFfRY3cONj
p30oVHFj5rmaY7crJejw2lwEsCWYrmldWrG0lrtNnpscJX06bZDKuSAyxuV4jnVd
hXFtx2PfXp6Ij/2rtwReSz6oHXMsHgvHcGN8X2w8pOwao83mvlM2uZ9CkHJoDu4y
pJEyfo+TWLdVlT0UuV4+J0HHQxP8rhctPpon509CbqiTVnBtk9dJJPhDmbZgPk9H
J96vF1PFIl5yzWLIgEqfGKyFTgVYQAMEjfWFsmLmHkTVWxQ0G3/poVXLFpb+vZTn
Iq3vlb8upoMr0xeMfkSDEVVsfdmchGT/rwI4tWD9slp8zlO4wn2qseNFzGsYu11B
fo0t7Z0ZWYWdzExH+aDJP2T6TYDY9A3DP2WTYGocdr2//k4noEh1ayG8pWLm++ry
ulO3MBPfIVleSgvct1iR/TAI6siVniz8UyKtqAgCWq0dV3B4S1UjaXjn5HDgHuY4
q+KGBetn04EyXxL6sW7qTwuu3CtfI4uy+cJlKWIS8tFtkX7BYjP2bR/8qCONehUK
19iqHmKd5jG55nbYoYSdyi82f+iigs0NLTxaO4lhmwBMpe5P/t1Nx2EN/O4NSmo5
OViLYeDUsEbqcgX8EdYC9ALvZ1onQqKnhsxxRNOM2yh0E4x8jDeqPeHB8szUDMJ/
gVjJRT1uGug4b+fIH8wZcJfzD+LdkAWaTAmJwAYad12+vkuSKpUJOUtQ+xDmoWqw
2Y0GL/3SEhYE+ogvNa1x4aciwVjFe0q/kO3R5yQfgTCGHFgIA29rQhT9QuMisYs7
Wqx7wmUtjuEzN0OMQNGaodLMYEp9rueXYcpd9t/G+s2PcsRaFBu69/DRc2jgvfuM
KD29G9wChqHl25WgbsmemCaGYwwt2/fB7f0QSJXc6iKlQzF4YSgQgjaMh+j0sV97
c1n0AhuKhpD9wq9ttRraX2TnNikYrnZTkPwS4LpJJgGRxz8HZZdwdi3Ze2HZVJ+s
rF4AewHMcGBHNrztBM0kurTT1S/J7H+22BIU4txfDBfRfX8S0496NjA7h6m20UjV
YiM7OZg0MliSA3jv6SE9rrXRe7W9wsawuxjYlYQ9Oepw7MsfdWu1ViHS2vztH67+
BM0uyC12ijBQIpNNzrc6ERTpgRsa3GplvkwmySaaKuJuVK55jLW+6a+766y9dAS4
cQYXK2zDNVtZhVvALcs6u+MYh2xQO+X4H8ULGrpBqRALxUyshh8lHkDmeRPtDVu5
Bz4JJQUFrMV7Yjd/16vmf2IbqhEbkP2Wx2OhROczaqFzEzNAV10CMzAU3MUn9sav
tLWwSsUNt357O31NNkOV4JlGxcG2Ysqpbs6NmhCtILoghWAC/035/fztucii+9l3
iNH3BDBEN1cKWkncVtZJFYw0PiKGPdmkAmZHQK7EVakFV4roQ3SA3O+H5W45hE7Z
p+TA5EvKnmPwbYiSTX+omi3qK9ATl7278T2RkGmIh5lODObo/0kwK8WSN3Q+U7/J
PeizRPSfN0+2TAiUarUrIln6FNRnxqZnBCkTnQlTKoFi7dXxRES30pUoO6STDYew
z3hHYLwf0vAEKElJFJ8Ehqc5/JV15Ol1OjfFbpTPR0ER1UQJEs2xiOdqt1qYdk+O
k9G58TYAjm/9EW8eHNJe7UVZ2Lq5SI2DJvAF9LWj3H3Z7Z3nhnU4K+Xm471uQUku
Mqbu4wdXyiDV/yJvzVeoBlOjrcNK0GGcXtOgWzDRPtiqplHmoNmAhb3wjNp8v1KC
IyEtTZt2vHzHx2c1EZ/XqoxvJfFKP1+1DltRlWjTuYhTINY94rTNjKSoxyG/e+uR
u+jhK2Lz8qsYw97BS35SBFvu9CKRnevHLCXTkceyYPIE8O02O3YODntUbbzjf76V
C+nAr+LxkgTNWcQfLMjAAxYqkK8Na6FVENdsYgTVbyUhKlMaaV8M8r79dd+zSWnV
4nIcw22z0F1VyKS1+oOKsgyYVwjRc5PZN+RJ+yvWBtCn2jVzNlAy5u8gIwu+AW0s
glejFyDJz0U4MKcCJw7BDio0xz+1q4TbGZTByoHytCZoSB6PB8o63zTVZwjiWuXj
zFLrgfeXkdJ5qrHeNs8MPXdWaLLkgvKy5aEzMCUoEB1y7sBqEHPEJxzwZngHbEiM
3Dg8o5uwkgBJsZ5EZuH0qt7Xi1D29NP8eMuF9P31TUfHigf9t7ZG7cmEMHnTI7JF
/g8/gEi8KK8cHr9bGmg0DZte1bL4jfB+iop+uIreEqs1Ho0/2gAN3na1k3aIetNh
LBWJvGVY8eDftBuoNnAEX82C/gMQR86NG6J/j+G9ZkHlpmb9no/y6ZARxiJJDBBb
r1klJkmJUdB8bv1isAJGFXNFrjO8cXE+dmHvM1G1CZGtJ++MvcUaIPIPIZTZeGn2
6Jsh2WWT1tqWOFrnhLKjsPxL3wAWhhzV/owYZUbP/8WjWxtYndM2/+2LE8+brrUO
D5hwwijXK9J9WcL+acsu9xdjnJp1ZQtlhFrfvFwbq4QdSwitTsjlU/e4V9b6lKVv
rXRKybbUMx16Wr4gluT33rShGAOtVZbWkedO/eCqeDpXvegqDBBhqsuWFh/us6w+
ngEQCHuAlJJOn8zwQ5TAKRo+5dcl8jOM8kkoM8PQz3icPcjUKkD5h+kTH0fSizNQ
sdr1HUlnDgJV4ZNfRVRYxrKczPHXyy34j3eRCGMUAQVc0WLqIn5T9PzJhNQBJ7LZ
L+Yfey/jKoeJ4EsqDabSTMsMi8BYY8AEGuIrKS8kNkkrjnfaVTCP/yf6wKEdCBz/
iabO/R2WTMw6TnEg1COKh4Ki3/xXfaGnYjl56Ywia6K/153A7rebPOHOdDSmDvRh
mI7a6BpPN4V0rRYEQcy8EKPZBJANS2DaTzkVqLvWxJ+8YYQJOsTiTarmSncMhZSi
eD6OdmJq7tCHZHe6DBBWEqtcDd4P0Xb1/nXsSJ50GpOZFIw8NBNKb6E/IEV9Yzzm
+xSZgagobkZ0Bjnwm2H1wIH3k3ZoS0zr8ORfWXHKL55F22ZYApk6AR/ue7I51YG3
2T2ux3zJ36xKrRG6Np2hkseh1axTdgQGX7YO2WsQ1iHi9LY4W0Al1sWSCaki6kRH
VrmFdYjDt8EyCLdzl/jHVCJnlqwR1y2xG+qgS3lXBUPToM0I2CZvJ6TDgcYF1qMH
rEM/BW05b5VVCdbyMjYm2/F/27lXcfSinwZMzZQIfydGO3xO/JpUehJAUnR/W6Sq
t4x+54vl9lk0/NKcMZ9weQZhyMXBisWIMs8gUyc5pl9r/KFijh6u7Iq+B0AZQU0U
myld/RFJSM2xOCb9DXRR/SjBJZoOpMFkgkAg9sV+Z/qBNgMTEZDqIzVZrnWzBWeS
EpYGh1Sdz2vn1yA9vMFq0lSLIaORT93xtDiZByoCncFZxazfePqz0d+imXxWUO44
YaQ2bLdOmy3uBEgdxqR/ATLgTnICjqLs59UyPa2+KU6i4j3f8cd9P+IxQzROtQFx
L2yL1QcXl/abEiYtf9mczig8WoHYMAQkJmGxLQoA1vytIo8inb0hGkEJZNm0oiVf
6U5IY8engjBmpbyI48z5vj3j4x/yA93kZKIeKl1p06Qe6BUTmAk5wsBstaw7XCZt
4GviXcC0Vzyii56PtfGPKc0veYNGMZXWbv+IsUdLbWrcKLU+oykNAx8AizhIZB5B
cep4pqV4qqFVrQDiMvFdSmYhlk6WYIgPRcWdXdM/vQ4NEVFbICrm9B8dKiPIPMOH
9Eht3RyqW4OL+Y/+hmhMG6N979KfsLeGn+DEGPt5wySOqn8DSzzH8c1P5kJsju+f
kZoglV6NcUfXETUEi2Q6KnhW1MYNbin3j94cDD0E6y5yjmyFNQT4mA0hnydcuIFs
ao1z3mIV5AoCyYng0HDnha81r2QkET5LjF72UAW4FooJp6HjUb5kypwhNJ03gwds
Ci20dtc9VKGxyQc7zKYpuACxuW/ov7Lj5VXCqfSoWA1UDQxbo5ZQ6oXS2Mzb46Dj
NaoAcAcuA/mNN/dNsjd9mmT2Iz5z2bkXvFUv7MYNtBREesMV8aA/JO4eqTzMwA5J
+wltShZWk2i2tOIDmnXV8Hs58MZX3hBEj0tav9FX24M6XefvOv7q2uN9thjvHTG5
iy8iBi9vkhsm/x7FsRTd5Lip31fMt00Wkj1/XWgUG4aK0F9DjPPKA8o9LqHGlykx
PIbJhwQHUY7w1mLjpCU3yIop5nOPr4/WepMoUAFL/RSEFhzqce0JCJgXNt/31FAJ
4BQoOdnHzQ/bLEaDhwhLI+/JAFqTPcA4pX6klWieYnMEAEZraPdoD1lMnuQRn4to
Q6z0OnL74+Q/Y3P8a14xHcgQ86xnI8ZU1hQB56EF0rElAk7VN5ncFdgRID3V3iT4
tpM0fAIAAz2QE6iL0pJ+jPOWWom2nO/6SeOyDBLgTzbmr7456HtsQj9nwz/h/mK7
EQvsbSktFS7yGK2vGKX/PnMogt7wMfGnmZZWIm1oVkGOr/Elbc3ubZjZlag2vV02
d9QJsv9J3kO/Rk5srtidyhnDAt2taEYNqU6MNdBjYyMJizxx/RwmY1wRC1Q2PYIY
uQeDRoFuNxMqeWY/9eaG8amr1uQAeXx5jGmmaZSNuWRWeUbRDyWiJ0L5ZDi4HyPe
yECeQVjzAmhsdVybEeC4Q7wT0jchsB2Bm20PT1z6E0ggJKBUdWol/vtF37ZrPcgQ
0rh6q8p1zhn+ZuKFXGZn+WIjEyyPOhANVzimMM4Wf27xjZfF9cFmJp9/gVw+FjLR
MJy/Qdw4mOi60xBc5lTK7GlErwE3CqKISin8XhVy/Gs4mcx1ie5Vhab8x22aweur
H5ZvYHh7axmO+Zwj3/SuS3lm3nymekFlhDPrcC3Ez2bQUzTOMozSvflFgj4pAnTQ
6gx4/UfNC7VzBmV5XjKyU5KtKVwN79aaMnaYD4a2nf/t+5KvrO4+mCMhU3D09RaU
S3zVt+3mS6JEtkzjzqJFd/S7PvYos04Ez7cxYMMhKTlcqAMt3GKi3wsL0ZmJ2kb4
jsOi2/KjDhGm5BimOokk2tyb3qToBWz3q6MnuIGHzUEytaqctqRHq/Vgr4GMUU43
PLOG0ov8b4oWU7N6XAucOIPFJeqaR8guBimkBqY73yvEVqer+qMpMX2YfweOmAjj
wLdoyleQVvMiIp98FxZoJPIA5DEBpiky31zqGZwJ08qaLIa2FO0dUtEaRynHff2Z
Ua+996OHNDI46Ocfc8vAS8OSiFq2kRhFp0sNGrEbOioPbrN86tYnYBopnR04Ujzt
tHKKEavqW5lahkVeJBmLWXukj8ZkLD7dRilJMADRZTRqO7Kfv96XUR6ovHxhxTLV
lZk68sRJxQawOr0VEmMZPcKNTycmZtMJk3Yvta/w4wLxUkuvAEcn4p+l+hrQAEi/
B5v34p2VXizuua2P/LvrXwvOQ1XJ+qeBkl3orN9sZieH5gVP6n2wYFap5R5y1NHa
C2cibeghJaQlxUgvp+UcL2JtMWpPVGWLAyXPDyqInygxON+3jzmx0vlUNbPUFSQk
OQ3sflQeugPsE/1tKxAbiyFYctRja6rdB/O4q/NqYW1V1b4un5Nl+Ys+B3YYNX8T
xfHsXolWW7KrrZxb/r/Bi6ORcpiprSosF8JoqtElmx2qQkPV6aLtWIzxjKC2eSH3
E5zlGvfEo9qZyv0V09l+bmz8GdMXVp6wxzDV4w3LcVENaaGorSdRoGMNmABvDumw
8ecUnTk/iI5rDgyjYkqYXPNyp79l84Xq0QnrLiWEXudVa3u4aw/7Sl8e1IhQUdZ8
pHXxxrRUIzDWrHujUP+9ZPok6fvb3WiXSKWtSDq/HiqBQQ9eoBUnlFEtWzOigVcL
3G6YL6Gm43jUDtyLyl9hKN3qGxpJnbmoorQ4P5+bhzF8HeBvGcfy3pMbwbDFOugL
R+8nSl018m76b75WhBy/V1bkJV1XUVD8UEFoE8efPBhRdMI68o/ARsQ1Eix+gfAb
25WHVwvMuVna3uNYl5lWneQx3nUIK/WvlvtyezznKoJNABGMKS0OoLgKfu6lviBM
b+vlo9AvBUrtb/bW9otGplknweT8pB36lIphFhgBreTtDutYNwlgs10uCppAzsPm
40j0n6KUWLy10nn/J16cLN2Glc/5ct61MM0dp5dkA31Bhy9LY97hjO74is7UENLt
YXyoGDZ5EPFmpr8CG7tM/xPk3FMLJGOJDUQblXfzPQ8nn4Bb/frPIo2Rsq3l8kel
JxmykZ3shjTj2cNNGZYML8hkPf3pXLEYahBsT2UA7UEmV62I6+0vYUAAd9qwBWKU
4xU3FLqiI3KRSSkR3H8wqINGDL12JgO7ID1J0opQEtTT0r3ox4RteJsy2JO+6Lyh
WKJ0nRvpgbzg0iWlxXgG7BxVoZNE9swS7gTGPgL+Hb6aglbuUjf1knJWmD2CnKSm
f9Y5zafmVcjf/epGblLeGF3V/QCix5o/ILpxa12rmIZf8gbAeWDk4RF/sklcSFoL
5eJ5hVfa64gz6LmsLG/xbL1Mncj8KRpMoYbTU5erXLEgBMbXKw/LuZHTLYmtRk4i
DO1RH+jtwthEFgxPPFrHMYizhhU7KscGf2VK5NUjHUUp7evAekJ2BWShvUqAWBoM
EdskNiiwOLogMBwDiKx3bz74MbS8swxwflIVslzgJWErZWNNgmL72kdRzWFq9xBI
dI1JZMOtWFTeP+4LnpOOkG4mnIx/pVCrazWYMC3PSlxTX4ZKvMTMFG8JS4sJq68+
RI2XMJrz1j8a6gBaPfqKNSJbmevepZfLNHdwRM3J21EcZS2WrHrGpQwcxUU7+4Yg
/sLO3yAucsUjXmBefgAg/Ko++QEYmU8sv/GWQPlPmMQ46pOUCqxCsTjK1SRdQvI5
zV/gLElzsTxL/FedGeLbNO8zQSyiFodoIggQyqXrxndTKrynxIpmw0pCNoMZmZHi
sQuBmWiaduQMyMZiq3eUjDzzYv2RfgAuK/WYeIoU0gALiUXc9YlauZ7RrbrdrQEs
v441VcXPybsW5H1VFg2K1DNuTDj8Zm6E1tCaFp81lXF5sdbGKDPo1OrPeHWnK3dn
HdNVjxa9BE+NMDAxktmUUZgoIrvYVLtru+wNUiHkS06jhUtbNrYQnBoKKHCVhLhe
ZHVbCq2MQXqV4ae/psdHO0wZl+vULhTcUzSpJ8c0wKTVhJ6q7YgE6/EvIBJOamoW
S3WbWBsZW+oeJTaZFpT80FzfU8EQSytYgLi7EufBTqBMdW2md2JypGpSdgAgCeNJ
W+3kkR+gW6SjdYtPlBLCmWmIKxfxAdVcwnqkjfD3gbVGpByCo/kXCl1Bd8Ympn3K
ClslbMxHxgfjxDwnC2LB3lAs6mL+2gHL4pnER7qWHGU9q+cLYir66xemuL+q1lfy
gUfNRqonz0kRq8qZqBYxUxC/E831QQABTGYOxUXqGOdik62b3gVWlSYyVOPhpJ/p
CkRtU6hlWYJlqRcTEcCbsyBnu8pZi76z0clm9Hy0zq97CqYFvYQFMKdYP83xSA94
v5wpF2Cs1aJQYg8auMiEITbs6mZJ3LlNGMHDH5X16EFla39O/9GZf6XWluIUZGh5
sWn1K1ExK7t4atiy4gP8fnO4y+W6SXJggu2DSyo5Hg9fXFHU0dIUO+W9xG+3+NP/
JzGo3ponQ6AZIs1Qp6EF3Q/wlxvUveJjMYWuWkCsZsLr5it3Zi9CrmaQgcKSuMm0
DvT3z0qOUJr6v11iG+d7ORusji5uBUDk1+uovQ/THC9LL24ucifY+w0Nib1h+9Wb
NZqAhpEiXnlRYnYFRxUzAbk3vp7g+NOA0OFljDKQQMXzxwJysn/Jf0rUorqNTkqa
L5HYNQrV/xVLIAgduUnrpGzIJx7W8X5F4nitr2N3YyXptkIte1N7DapQ64+kmaZV
9rUogXG5D0FP9RlQNiyjLVgLxIDnWYsPY3mxNdYrD0gy0l1DwMafGzu7xu8p7nTU
n7PC53OZmGDLpRXo9UlCfD3K1wsU+AuR5C7FPObeotZdvsTXytu9XE4FYKZ8i+N0
8scSTEo3bKapd0n+kEc+enrtT1h8MBOyPrL28hl8Y9XKp4gld0as/Blsi2Qveo93
Fl/6q3z5BvtvVYo1qeCAyrc4d4src8EjGtohNmVA3on8thkzN/dOLsWzYXekORzg
pZkBG6wD8qXWynXNU4zoQ2WRQbQxjb81THJaKGij/G0soKqd7FDPJFdrp+5NerYY
wZYkDeMjUyILiaIQZ3S8xGCTw6HgqdvYAmeDJU7WSD6o9F/YzLtpVSNx9jaYuhXV
fKO/MPecrX/TlaFFCJExB7QDfJBWdC5clfA+6GwDHc4YGyTWs9l+8xAxLlVFUAmH
HnEtsy+fsVPP4u5/Bw5mTqQv60CTXN05ElIt7f6tQQadVG7OvbMVrqXaQe5f1BAh
cUTVV315+v16j06ATaZaem6d3M7mR+heL55uB2WYdCmvXn7IHCtDCUam/+UJIUJo
fn+yIfGqpOWpEz6FzO4CHhYmRr+uCSO3VDa+QoedJr5KU9rbamIhXqE/nR0uGIra
+Tz1KfRgxR+p2Ps6Wvlxeepa5znWVu+ruKG6mZAN75NT3W0v4aD5EA6izmbH2vrt
cgBtEntlzQVj6hEwIps9C61LW2q6KReO3t5a/fmnW3TyNwZDvf/63g7cc+WUeuap
+1CLR9XjUPLc2o3KDCWNrfib9PTBtIIOuPVkI8HVx032Qo78b8AGus4jdnxKruil
oMLlW0/eCL5dOemHRVWOl6uHnJ9wITWn/L+ODH7HuT7W6YGNrZjIe5z1piinwjO5
1ISLSZ6+Ao4cBaVz1d6Qnkd4iuUoOSB1FQ6YCAVW9b/Dx1V4FdibOr25Sq2Uv3L7
sjKq3lqsNngiCrHtbvS5QgYSxOZK9qq5KGnnAoCwqdc5HYvCs9KfRj/LYGlffovY
v5+Jr2rJZ45/9oF/qDSY+G8xYsiDZIcpagLJreenj4m2sfO6MGifhJifnib6hAHi
4MqX1jYyPOeNhP79N1xN6wyf4O3Cb7LL+6IhQWpJfY8qaSkj/sgCxXBJmaT88nTM
fieSuL3pmCGlJiobrYXQyQicB1SRhjrZCXJGwNrqQ03LQq11HM/n5+8ZQln6laG7
iwfTvnuag99yS1x5wwktQD2TtbKQU+kyQnYlGuvdQI6GkXalDFKbB8XGK7icJM9V
7L9Gl+mv8twPZHlWmNCq+NX5dLT64YdFyh8jzbYp3ui1kYopNF0yo4E5+aBMMPqU
DvfQInpWm2SGYZUo9GIQhb9qJzTRq/HZVb2DR+p+zHeHQuszuWRPJ+QXJt3BwkDJ
VbzmQbskHyTNA7o6Pan7nmMRROcq9XHsfiS/CQiKPiKfRSfHg6pInjfl4wsQ1x2Z
WNtR4pz8emVZ9m0HGUAJhxsNBRaFppBO5GmBuarVlXmSsNDQSluQvDkCahvMsM5a
UNxRJuokI99PseYzFBkRXbYJXg3EVS6OV0zquQoMvxZqXYKx1BrZSkTQ7b4WwtOd
rD2Yf5vKdVS5ex9jyH+B6gd514zT3hZOrujAZJzpt2GvnXgHTn3AhMUsTzCLfG/H
JUDYGt0hDCiCjUDP6/W7u6Fu9V75x9y406yUm+ZpneY7l7yDxwpLpwMPQCJZbb2/
m8/6zH/plX83D4tiV9rqvcpzIe8aDJXuF2jHvIMACZ/YzcD4DK87+WLVKAahLMZc
WQ9n2ddXIUoPHfPJSgD3vqMGnGxH4jT6pxBHJvSvrovP9ZQv9lwlIDsQv6frvNSD
6u+h1kTFW2/HPPRTcrOo1e/wnM3gXrQwvRa0ljrjhWSwa1Ka5ZzenOiAxZFXkJeL
3j7jFdZu/RTN8Xr3RhLU5Y4KeTmH0k9kpuvb5yTkgBKczBsY3kSw1QYkRRTPqZp4
7EDtFFVXUpxWL/Xcwt6ncToOOe2vfH+7hz5oSVleVDC+oS4aG7T17a7C24Aizz1c
CCau0WH/venRkDY40d3CDiu/HEQWMJ3wMktndHXz9wERQyWe6nUjNoLsete+7PtO
QvoPoCp3pywFsiuRMtk3/0m0Mw0GMcWaJv5dg1YLFiuHr3zOD+vypINvDtatom16
caeLfdcgJQ3EDI/9qH1hzz89ixXwMTZaPDveM+tFS9fl1wveWbWjLLZASom0T7op
S4qL6SuswPl4AYHqSkcqZU/hBTHhs3g5SAhxzMBRil2XKJPAg0zres3DWtwOdPNZ
lb7vSZLbtr7jju1BS3X0i9fpOwJWH3K3gj2xhIm7sr1A5A2XWmDlVm2R0G5LRGBL
dVkDsCutLNeROk3gKsf84Xm46OoUKPvRxn2+Dl06NXZM99zRAM533G/VmVA2ZIqa
K4K5syIuC0P/33ZKpVini32Ak5JQuWIV5EoGTIXnu1uZZOL4hM7sCes06NhA3G/C
5b7HQGHaYUJ7KSssqYqcQc54Ud5Id4ogC403hnVvEyqxQUw80JcLrpYRGGE7I5Ea
c19u2RyaoT0xzDRW1xedGPceGXjcp0vmpqoUhXvEyF5kGFDm5mHoh09ztZfLnhDH
LU01VUN80FuBn+Agv1V2AdRuN5zwxvWSBMcbDt3OOOsceBRTAwE90hiABKpRcmS+
RyKEOBTGqAnST9ANOhrvQoG9ZHKGjTx+xsnC9TXcDr3p7PtyK5kRJBuH+ExruBiv
+kZlXFIujC9LxUX8WWHwBo2fddrwft6EoRAJdzCHZ2uEt4DkoxYwlQ67J2R+t/k2
b7LdIP/lMTTH2GOqyBmpZQGleXMUwQDyGQpsL9dJhd1mHZxmDm2luzSgW0DJvIaY
Ws3cphFWcPyuMZwAaSM9U3e9aakrnYd8n1vNGsa2Nbd/0qpeg4Yd5uHgfVTYwL9q
6Zm3ZCNb60sL4hvpCRB5UhQ8m1MB9X6CPgnQXgjzMtcjgAWCV/EclRuHyCnOfNz/
wIrOgHujT/axc/rXuyRZeGY37jhj6Gm6MyrRTYq+6ElnQPXtfWRrc8vuRu5iIvQA
W2OaKAC5HlcHa6LWmvrOY9k5C0FwXGB6QEwxETMdrvorjQQ/vVKcHm1xOY1Yn2KF
2TIa7DH07RXxalEMqfNluVauUx001pDooxuwtGxHea0WrXApLN3VwDgeje4e/b6W
TEiSQBJ2XQiY+bzU2ilVvfZBo+XgrmFmaoUsk8c4wHrrJqL73BYtZDaXZafsXPdB
Qq/3T00fa1KJDa0orTPs109kv4lva3bkiLJHd5yNpKKPcgRmWvxxNWdWc194urn1
OfuJ5/WrxVRflMhiWXwfmMrJ+EYVuQ7Mr170I83gg91ddWWpR+L8pYiSiXJERR8/
qb4PKb5tQ6vbjJfuwXnLbk8EWWVMHbjCTfhOF8UNrs8wt10aQ7AMD1VmLfmAQlWk
1ZYGAHsZqkZ3bQYFZUwSZp2Kh20ncfjkFKfv4UScfBNKQxX3D4Zj0tGGk7CM+61W
mmsaugrxhPC88nM2b5Ppn0UHUd4ySRLa41ZgZQLozZadAgcSq1bg9PPXyp7DZIhd
aUmhJbK2QGkAVQakH2LLru+1LOJHCx3TEQNUTfhLQmGLcXo8KwDU7Pl372TWrxCY
BTOSvnU4Xw9FkHP/RipTXNow2OAvYGq10hgMFl99HGh+h/QTSXZ6X9FYDYwF4qIk
iz0TaGzbhT9/lqJa+rGfoU1U5f8F0KQ7H+8MCtsBf0bW93g8uDyrOZbZxf/R2DSh
b2ApN3dg+7kL20rMrmEvUjTpnnQmm8Ji2EZ3eMJLp78fp6bUXe4+Yvj8cMvhPPt3
kHIuQ9AtgPkaK4tgs4LCKwXq7ZGx0yXWAhXRZyi3ZY8DZhijhpoCvcusehwfvMNS
jeb1fNn0E9KQ8q4arTcoojSRG/rC/NeeTHMZr95ou/9Ll6kduFeJP+sk/ueD6HrA
4moZU+F14D7USrJ4GhihVKSKdKgcg++iGHvgyZffway89joDTkGvNFEJ4yH+RV0F
8ExMxWEXLY6POI5bpx7yT/bqyNCm2ybRy9KFMCa//OzjMDu377u3pYZW0rvXpjEB
TinD1rPYfzyoWVuiq14PvAKs76sZ7cUPQg04Cagmcc/qTwIQtiOe+hTmVTkumHas
izCXnNJQoDDJZo+h6A+B1xF5vTpuhUecRC0eSFHCeDaqV9RZqfEY+Kjon7GRNWTh
BKd/mtX9rJ5hTyw8cBa84MEgiwfBo/pVSCOPTdMeYDBGo0ZNYk0zwfNjKRX3de9G
smJT6LlC3FaYaSzzw9afkVhyFv/TIn6Dj3keF/UzCIXGdGNJkprLAu6cqCKv3pNT
xWWZodsUdD/fQeiTHmw8aCcysu6Ppw/mCw9vW2+jQr7uo0j7DSPv/p50SRQIJnjp
t5vDFo6VOhD35bbJDwPXls4ydSYnTC+bANw/wL9hphZ/y2D1jGAutnQYGOuAo5fd
3hqRD/Rb2jlpd0zFzFHd2LDIbJqUBI3QOx9+FgNyl76XPhit1cw+5LD1zG4LC6BN
FkYQPP3wr/0Jum0WKBVkk3blLirNqPj9fkOV+XMT+h04e3/JD1ydqF24lk4unQUi
3t25Qbm59FWr6EIk0L2SovQNelk+YFM9FQ9XvJIRm3wbpiEDvxLuIB7Z4vbPLxO5
1hPFjtFJGELBIItVz+1wAJM1U8xmPlo92pwrRTfkndln4QsD5rN2d+p9tTr+y5zU
nY8XqPCPDZpIY6wW/CbwyIk5Po7Aozc6zCAnemVq57ssxLYV9U39C74X3n0bGmxB
F4QKE1Ch/SoXtimOrGbDhbaybh//ZtMWOhqPAhnO7n65BVvE2hd3EDBsZ1Arjw0f
TIXftkcctW5IGQ/nPISKUy2aGhrrR43uOmodosr2TtB+iVlLslqTqQfdD6sTL7j0
L8/FGyr7GUaaIscVvTw1+V6aUZFE9g8K5FAWY0TozGNDaZSVmZE4KnoXXLJgEQQL
PAkoeloAFKnXek5Yw7qEHf3DD75neYmE09JaG4F/KVrEQ7hD3inSTtM8eaP+NLOB
1sacNWZWeQdrzthRfX9M4BqLs1bDnr54pUe/cD5XZai4ER/NIlkSX4dpLdx7d1gR
AdJYJ9CHle0vjvAzuW2eirYbjxD7qtZwZlmIF3HdOqjIUbwbAVRji8dkxY8RE9r0
hBW6SULfrivoDY0RgspbtouGoqktTIwFD2/hDCxW8cp074DAM76mErqm1UVnA7rO
CRESTgpTJWJbl0+ya9fWTBN33wOocKpmzCQvkcpC59VQLLX0p+k100l2OfTPQsPB
TJQpMOZKI3z7+rAAid0qmkxINT4qmgIXjJuGTvG1n58MSBMRPY4SFE0LAEGAhIDT
jGfir1euit0JF0nPlfFXROotDduyuXVYOjbAnv5YJn4A1XI37MkZ0vvEYvoZe0/N
1kMW4xSMarmeZHfIcmfa6j56K92MiUkOwYXqdgArvkMDxRjQVhkqVLkoxTFCrW7o
qIoR1qH9FI8qOVielDs5WQSYAp9O2o3mZ4LG9gDGR28C61uOnLdG+Zp6PTVTGSTl
Lq/9p6ZJIVFgPfchCwUX1OpYpIIsWDCjytXSZ1qaW09YjD56rqNIkP1v5FBGnihp
oRifQvJaunKXT1tcuJ0LRmuiAFpSt62ngBX377Haz3v2EoKpzOCssTGDimlgGu0d
Bg2Gi47GBFEwvDpcyA4WzBVfNunJaKzw+TrdBIA3SUQFcxQ4LbmAqw3BuSbb8iL0
CJZvkXr/U7JaNE2cP2HZMpTQb+yBDWxmADg9HKsQE2VI7jxx1MEDJAoGB3AirZnH
VQUCawnTaY+egE0GPpQetiDsG6SuNqS+o3U2LU/av8bmEmXEZ/jXuY7HIN9DurT4
U3E93NyTAL895EvEbYrdwxlMYVFK8sq3mPvw6wPMKuR0G56Nr9Ch1i3kPRbslXtu
X7EjySne5fYMAKl7V4+mFrSxphqVzYrzYyZiPAqif/sxNvFgjChkPvq8hF2O50Lg
Rdzu0C0FequkvkV33KVGm2LiqcfHDGeblzOUiz3WaNW9bTQaC8N26oNTrIvDJpDj
GxQFA/Ip7wcm2B293LcRClBVUm6iqJgeeEhiGn+4joMT6v/Gt6/oehR3LoBMsS35
Mk0B8ZD4Y/3Ub2Y8ER3QV3Fbc6456j3WpqLw7fN2PO/mrc3MALQ+LKo1ocm8D2OT
IAsSfA/TiATi6e9njN9V9k5nTeEfQIl5/ITciMgWkeYC5LZtuV9x1I/+oySScpeD
Uyr9znis2cunqQhSHoex+iTPw/8fOkF2lH17R6032k2EyOZMWI3xvL5mjlEM2QTt
WQ9VHRVXfevyjWgKpipx9rG3i4ADfeEkJ/AQtPrmuyLwnhUDq/hHJkJA1vvyVFDn
I8Ed9LxjBYGi4X7FiO2p2USguaqucyAId63VGJ74xDBKhnBVdQk1yo0KnOnEBG16
YEDQwi3TYPtD8QdpmwMEZpdbM1My6ec9LUpnYdAtB7WrlLKslx2upbs2/+fE4AF6
WNAuMLbScID2aQmnJl1XYW/T+AvFf2BDfepqy7/GRqKiF3qj0Mbiik9K53wrwOUt
K2aKIxLT+Qqub/6rxYoLotAjM30nqqzbZW2cuPaZoh5zwQgTvusnWTABWd0M/Pfj
OvtJlYn0QnEHV1Pq1IDbN/VBJzMtJiUd/UDUk5cQ0s631QRB1G8LrFN09che2GzW
b+Gdmf8ob8j5izMFQAcggYcaVl9BKhHToGVXJDUp5Mpo+Hfwe4RIK1018thA7BR2
X5AhRgU71NAFh8rxsI+irPhVHu3YvK+YFVoKO6uMoNDrQiJvYT6YH0P+xObdOD3Z
EFhjMOps0CNVjWnhV5H3VIQIORRhVeXBNSekcSFP14VmhAMDr/R5LIMutOPcysgu
lV91DFSfz5LUjEdrigPyz0oML+p4m/I3GFubcqTB9RzyrJu62jXBvKifLBqTzSln
nNdssd1sz7irqDxIn89ZvbGEYBLOOf72VWWb6J3J3KhR165JY4zwqA6cSQOTO8lK
ml2AY3oAuDV/PQXHaXVqmSOgdwLco8bvLxzlTmRbXvliMhdFdKLdYrDhhCf8xOX6
T9yp8Bx1QQttxNgHABaSjjKpQPEnYM6BZY8fQ/Es38uKuTveN4Y/gMysTTW+3+01
XcLDcDalAIJhzpxYVBm6xiCwCwmc48nSWovqcHjFAkvquugYhV5d5PoECYkIRa38
Eho4XYWi6/G/PImMFLQe1LjSpLLrBrbVAa75SrA/yBKwLDRR/FGymDmaS+S3D7v7
GNGKrDd7jAyIttYJCLWh1visqLd+E99gV3ftGZ6x0R23AGDuX8aQFgLlLgQfyBud
rYCknQAEVs1UKvPj4vLwCOik+MkvIkllnS1b3mxA5o34VWCNrinZtWg56jpT+yGB
BT4pYvKh843DwsbCnu9bkYuspWVoqYd1eyyqDuU9uPlhRCwNCLEE6Xi7Es2ZkCex
I7v97ooywwXyQ0N6kzbi4brrc8zsg76TC8nfn0mYoH7gQMU3aso7V5Rfyy8Ynxmp
UERq+ytIH2kFL9XpVJ+q5CELnLGkfPW+Jkh0l7lyRCMI59Za4TS4g6aFT2Ggdscc
yvCtT2c2Sc9xM4cdEIdglqXvz9SI6h+zwzXqc7t2QlcK2WU1XZmtNJTivnHfjG3I
02EOegvKkVPJb0fB2K78rrJ4OR4yf6ofSTNn8S5c7wI6BzM9v4GPdTF3yOWFn5tG
P2Asanz3FbazIJWyA7fhKyVgzeYjVM9qLKGbWEw7NxuOtLbDMipTvQsC5xSo81qs
oZewEOmtdG+J9uC23UYXX2OZgwj70k1QWVEKDASOkAghi+0Oi7cNE0taM0si29Mc
gRN+RzlPOQ7E+3JhcYUtpKxaxEJI9k8dMbeHWT7lGEvP+XEPxwYW/rG5h0mQ5aX/
HukhyW/BTJR5xtY2xKdH0aMVRiJb6N+wd2SZNjjS0ExsRUPKUesMOVuJnbmYDLpf
iVJFt/+i3gDw1dqSXCgVrQJsxHAR+3W5H4J+KfbemBSvFl138B+3/XXPqks03NfL
LW40ktx4gcFQ05p+/O60fOhNEYMOoRkGCmn2K1Krtse6lLh/ONeCq3s1W0EgLtIM
WICn3/TMGOEfGptHvqlbwOt6Ej4sKLHZVQOUTngmyr6THcQtQvPW6KnIZAyvkhNG
SBuDynYnNJwYJV6B//NJNDuTHNveAYQMC7ttDbis4OM6QQ3g+ERDfMMq94bpko1K
pFPRQqbBXAyUObx0Rv8deML2z9XNKgpgEdadYjdCILk0b/F9av1y48jhtcw2n613
r1faL/etCAr7NLoklhkB7Eptq/xZng3MU3K5TV86ERPiaw9tgeZ8SDWFKnKvFpuC
j1dkDXvI7Zf4wClS+AUT7QBZiOssDsLPE57+Lls7E9y8fHu8qdbzqlX72lcLc2+v
1AYr4kfQj/dAz0D4ybCInV2L3cLId+xrrWBfjG0pthkVvtGggCs1yXoPrLAJz7wf
TN4wUEQ7zZHTGUDVcjIW/4DBL00TF26WlDVQlSpCWr8by+aXo8J1iE42zqjgb2Tw
79k7NpCiGf4snqWCHrkRV9DVMEsY0GZJnfO4+zNNks3BkEiFu1GHbadXvy3daVnV
qjWhNjhNGWtv21flQoDcs1lYIPVuXAV09FGgXduXmxzyAbOlQ8iCmV095cyByARI
1BkfI5UtrmLKgb+Mg23YxOkJYdUEj8XDkmcu6Sv02+uQMaqws1qBmC8RqG4kLOli
CM7hWO5QLwMYF/JRgE6sX5WwCZxg2RZ6iaxlhHKX+VNwIjtjmX6YHzvQoWbS3Pjn
s2d/qzUi3t5laXczhwEo3+tTYcweotqzwnfVykVJe8jFsSDfNWglvjYUauRznJBD
a30Vm+uzH5vLHPvxCcw3hFgFDzpXNV61XSmFJ0zqrlSHzGbBqkO5Kw+jiMgzpq6A
3cJYBhO5yvTMBzGYZJ8bT2pTDb8+UUvBBWAe3XFamc6bOlq6IFvp5YaEuqF645Ag
TTSHsGYFXWislrpyvdWqlgS8asxYQptJSnnrUuav4a3k8sfSaYNvgKBTBh6viIqA
/Rg0ahAHtLUSCmd3x026SdZxtiTkVruViaCuIWNnUNb+1fMZj9mzTXOtDspsD26B
2kLpFoumjphKgmO+UoUwKBCyqTnCIcepz1H3NgYhChMHn4BBZuDL3r1yLW67U6xH
8uFJGMri79KG7nhfVsoQfveYsxEjajYngMmxTi5GukwvfeBhXO5W+rba65nvQvEk
8Z0wfajSi0aGlqdhXRNmBlVLktDJI21jOM+cDuu+Tllq65KDVJ6vCx9DKfsqJyLZ
9LXCZHjj7I2LkPtgMCFJjIsYilKZZUgurPl4zrSPktdgdolGfMQ6kc1ZszvXDQpq
ZklWOXWZhkNDzql+qocJRLIhz1jGI/talVhVdjcQ82uSbUp+PfbBOxBXJNYuoxfe
oXJEMtTuu+oK1HQClDAqK+Sm5vec/oCXMIrG9NuWoloG/pgNgxKXZRPyCz5Ybi7y
v4WcLu4DSsrclmSyZl0OsnPA6cbRDVe2eHFbye5Kq6xopZkEgj6SUD29udkIovYs
7D3OO4AfRgCqGke0QJPG4l+eOeWXS+ESqdXV8+F1LMBtzB3TuhjLOixT2A/IfZfR
6/M2SexkzG2xpO1yKExOnPkZI/kQhOLl1oIQJ3qfUtYhT0teUX2allcMTlq+hu2E
yTzwMrkl6U30mr4nRdVRsZxZqJOU8RCoUU5dGosYzJ8CLWkymhj/XjKeBzdBYHA+
Ps1yVfAXbCA32aZYijhMrltqnl+t0j/S9mxnsTCeEuOsV7cZDGIHU3QTRRlExAS2
gb5ggDaiTIVA5y+s054pBYKSrMI8RoNd7iM6CzZT7qQPP7CVAOa0YMWCjSdiMdnY
gTY1FaUbEyeM9c8iB7SdD3dvrh9zaQAhi64gumFj/0i14DCIF2mkqy7uI9WHLQKH
U4kO4m1aHSRmtBpGh1w2O1pKPgd3qML7pwVhlyQk1vXcYWgz67VDCXktf4U5P5df
NOP/FBxTUpcaYimG4sLG6wq1TZg9KgDn2oJn/uc20c3TjuNVKWMaA4rhlv5EceXx
ZCHt3sg0dVxhC+qoNxnThgfv78AKrnwFbg06ifG5irlaB3cSQkYon+/tzxuE14lj
804BfQapp+MeraPfeTOe5UGT4+3fxA3Hj+ro5ZxZWccszIbl09ehsgLrKE/hDf3d
8ZllaNanDpuXryJCU1VDaIM+ThDh2QrRNCuEL11r0umpEXiUMiqvqXKBRmYxzvAA
urmaJZqyHQVCF5PJufLUqpl2zVKZ67nHTUHv3Y/LqRue5Qw3l+pvA1CcIw/GmxDu
GXUyjcyeHskPPZoUgZMYr3bM4QROcfOk4m5epwotOxxpebb9AsqggE39B5/A3Gqy
9XgpiLarwMUe8pLQnT+2bnoXbHDfIG0iaeg1Dv46xxh/p40CjI4l/Ud4iC0nBU0T
BOdA524rCjUljcw7LRAUU5OYSbJEtas0OQK1Deii300bFzjBH5qEs+Uc6ulTa7wx
10OIcLGxq++qATjRJwxnPjV+UDS8ULFA/lKSPJB2XszKM8AADVRsVnQ2eNapId3s
GRis88gUBtVgZgRxxmLXa96u1Na/n0fLZFo76cB0h6fyQhr4uajIYal/DOdp+lPg
0iRG2Rr24/leK3itl18WWZNeSVHQmEPiNCTXTb6Cg+8G1XijAABzhNP1VsgTUpJp
tiJ99V1CD+Evp8+dkbOh81CeGrOM+QA4RJbDaYHv44PDEo6OOlXU0gy5Vq/NsXLN
bY8L1q0P0TbnLvjGACVCuLpgbcUDaj5NovDEJ5aC4T1TcFhk557vWVK0v06vkSV9
8LG7yqRFFcORCvAoBhRg1xDophwkBFpC35f0hs6M+vhDZ+QUw9No/kSnIJ2s4PKt
8w19RGpB/6sAzRjs9ZhnnKeFxgUf1H7+kAXY7Kpj5J/4GZFzPwo4fxesY3tP3gjJ
FstU5evKPyB+3pFpf9JCycyaK4NM96T8M+Iyis9rC6dR7HXyQNBnfLimQPCb7FkR
Ts4R+5mpOCmAKrAG/DrdUmTs0vEyZX1zmHVgaZ1xGCSuogJHqOeNTff25XHbPsP3
omSi9x27YTAcI2OMVD9jqMGJfOtCQwPplJ4hSGC+69qshkDn0fxWOnkVZR7v8452
jJNMmNy2DJh8l3ZMcU4SPnwksmjp8d0G8QNWPVWIRfCHSN0F7AQR+lgTRlfHZkR5
k4qClZmHM8ukB8TWAgsaWv5DmPo16dE7W6MZC43dIAPBYtvSynyREV8X1HltMqid
Nd6ju2s2OKB3B3isW4RCmkEfYAL8Y5BQ18WJhUDyARtDlw8DBCdwFzL4AcQ5786W
o6ZWv2Uv6pdlIqU6r1dz9V2V3bnuiZOnH9VUN3uPOFsW4zrmXPa6YLI5Imq7IGgf
bWm6HvpBjLfBnQ6X7cL3dhvHqM+PPVJ219vgFzgSQzkd2yHrP+EZMrY5gA4oaoSy
9OghA3FmTQe0aTa5FUTIIO+U9ZzzBhOXt0ovAw/fPLgGJSJkdTxES/eAPAuQq/3s
JS3XOPzh/j1jlBWZszVu1oeKYgoUtQMlDWqK0x7In5kNJXr5lG5zHk9rWkFRjdzh
lGkDo7M7KsqeuiOC/ePd4GbyccYWBU1C3f7afLg7ysEcbgjuykpR06DilLZov4mx
DEcTo3BLbvMoam8wZFsR/Tj/1GogFiWdU0vxgZ7ji90sHTGAA/l+qXIJpeAxtbh0
KJYJ9V/TSx+FgWA3VS+C7qFOLn3xEh5vlKrMwA6A/Npcqi+jThXaWLOGVjGFPTGb
GNW1H3wq0QU/Kj/syfufuFhYzRuJ9A2OApNso6Gnrwvsc+TX9pxKlbVjaM7hEYsy
FDm07SwsvkXOfofyNS5vi/O6cub4rYRK/A0dHG3xHg0XU0mHGPTfSdUN6VeYNDaw
6iZ4/I0+7zGdoCz4KLmclduQjl5/oiyUFQ76E+TrJgQ7sloW3ZRDkDD7ajs3YrN7
GuIh4Q7i7PfwgrI74pbH8FA6JTUELs+ePVtkQm+ikYnUNG3lVAg9D3AN1tHZXobd
9/jhJ0lakq7Q2UBMEFthFyirG4esfsJdKJSY6ZBynGcGTUrLX8ntani/Ymi+3B+T
8kCh9CM8hLFL2+/+R7I7yVU9J3eby3QenPAoewjjBaE9vlcoZkSPNTBKbCiUvlxm
6uyI017IPaK9PAPb0WGYMhOYnykkEmnei/Fo0ZzmN7Gc2TFvR/DZmBdgTaUZuY+n
hGBTj/4Gp4YuGpr5rgdjkDe+fcEP+ey1EMQhu4qcWfP49z9GDsWj3oILJ3COcnky
CMEZbrrf4VMcbAzpBB9esYWS0UjXGjEb5ElQc7MMBmk4z6wp6gtQgoezWX5+Dyap
u6//+5vtB4xLIWy9TxlUz8vz5xbIMv2dHjJscYVtVaea9/VimVZ/5w1UX/5s4IUl
zU+8HTiJIcjl0J3Bzmf+WG4yG4SuIJgpfkC57iY/Ea/Twh/E08MEjlBwxBR4633S
pB/Yx+N1YKvsXZUbS8e8xIaZX2PLiSm/+AqjeLbjQfC75/uf8p9YrBEP75eUyFyQ
QcskgCKg06sKo3FtrDxmcUi3fllJWLN8NpusMsTu/yWP70M3MR88U9ylBIoye6aP
HsRU8a0ymChmdLcqe5BjEGqGe9Fi/h2KRoi4tcUASYk+EOYwNex5vXtHqaBk+ghG
qgRxVaKzINsC0PUe/zmJEeyj6rp2SKmWjYeovsiwVEFmZq7Ej4SGyzYQj2XHvX/m
JMNR/MXjqyFuMTVYq3J0hqUYJVOeoYLCkWbNiCG6P/bxiuyMFNluteSYKnSmepDg
pTmkBTBoul6SJ396MgNfNwvI6Mfl94cjOF9YcQdWr23teh/nEidDqgPn0pnhId6C
DOmtpfSDmR0welcKwnO+zChl7S57FWGSyaACRITBfHtC8RRm73svutx+z6yvKRKs
8LY72XSjFe6IwL9MMBdaSeaJHSxVtdWeUFK2sbld4Nda8180Qr4bPapZUHBAwj/c
PxZGKtm79Ke0cUvAJtIscRRvq4ginkmIBh3MCtOtYRdKqCrZ+qbVKGyVdcdisovu
2rPWZoRYlQAmQBpCTqgKzs0AtSevrKDFLA0yRtEqM/EwJLbjEOudYySYQm1hW7D3
aWDaqFpoc/SSS35jDWURZvZFI8pAjCaEpDnQoZs6DIKpN3dD6RojE5gVZR2BQd40
JjD9dfQsuDmzGR/p+rkSrzSb8FvWjcAziR9ljTrFMAwX39Uagjn9kHHlpvEISove
wqUTkvnZMjRdrRaGiZHDMdyA6gbIkx3SeplTO+qV6k+TBuauJmmuwq4TdnlaWOVK
HUWf9eoQuc1Zq0moHQYe1CSncbKAl/evx06y1zDmCisHC8I0dGHYoOdfxqCWE6K6
CTEmVWzHj/TPxheljGV1ZwX/5GRdeDTfSxE/SQs/deDF/HseIZmnf3dyfsVO0Wax
3XX9Jl1ALjFITDxI8IDmxVuE2N4scv6bjCGJmrKziCaDIipX9Y2JEVNuKPDuty/P
SapIq/eOQ7uUWsV+AD5JOIOqMREn0OVd13g1Tl7w9pOy2GoGn/J89Bx9Y+MPo3vn
kso98EI1xa/oLnRuadFyNPaehMGEah5ekxO7vMM8Sp6cWWKiB5ZY3DI0HKwyA0Cr
rB57iHdaxAA/paNRGOu040hm3PS9ij4JFtvoSsYs0SIAYiSD+PYSUhgipwcchVP1
h1AY4EJWLYVmzDht0Ee/CYpEqRVJrujlF27K8XIWt9dJxzMpK9WhTss/4qNHgOev
kaFehCe+eUl6S7/K1AB4aF3ENhz4nrdcjMAZ3t1oPvP687yDrJu7vQhgaYzUQM+P
oby4CytpQC1UxUmdRBB/svKJIKvjZ8MlESPnV5JVo2h4KSBtKNr3kv11oVVpQgFU
ir/+59hDAhttddxetPfPiZ91PmVVlhcoPoYIgbpGaSaUu0dkRrgMPV6TAf2cfxEg
3HRQ7pVJgP+hWfGoJMsMvjgku4vmvzPFFTbzwAWPTfVDItiRatT9v60N/eI2wGD4
6RRI2fD+pnWB5zetJuwKVU14RO7NQycSCNYIB6zmOL5d/geNu3OPtEYvu0ahME5w
VjNBOHxVyhL5hCBKmxC57Ww1JvysLI2sQ1pHGL0GlYhd9IAudSR0QKwh9BQE+Zhn
C5UKsbRixcKcTgyxShEnwQLMELhgnPfdr6SBVZ/BsfNv6F1Q1s+N/0wnEtHhiVnf
4IbhEQ3eogKy396v3GKZxwKUOe/UCkfBfOR9VVE/w19DUynZ50pj/B1AK52OZXgv
WxVmMEJI2Szusoa4ck4e3jMeGhB4RDXVyEGL49UE1EwxIvrQ2OnbWolx9JpJH1EI
XrhvQyVQeU8Lu0vmRIG5+Y355sbSMfRzFqwCWeO1UM+RmKUFZOUDRR1eo2sWPt+q
wcCjG7fUYZ6cQrNTFRhag6KqXUOUYkUgYcMHpzu4rt47ytuanN5RFcVJFztjn+wZ
NmxNky6Nc7WICEbunTWbFKcm4v0xhj7tmo3d2bXtPXte70HgGKLXYJrUGziO63Ky
J0zsNtyWT5mHlxrEZ357R1E06w99dJkgabob/Olmgp4cK6XEdWLepIylX7MI/FBs
1h0F36qHzLbhEEyOVzFsbRUtyZY3/SX3cpR2zRti6Pxt5DaGshf2IEvpfsOEEedU
i8AtrebAyQkEE8CtQWm7k0Xcp2KYxZfP1LOkIA2NyiZz0pTG08LqINnVBNRQWyK3
Iv3GoATjVdXZ36qql8CZkdqpZdU/KuhzjWPTC3YVW6EMAzDVOFbJ/5YbmqVIZpYn
QKWQYtdeT1BLdSs9K4opHKlpUxJveORyAbCxoJe1xH4+sgaoZigh/lG+GF1v7kwQ
+jD0PIfCFLq6+oU9Uyykn6DUMXM6lMOyBvfP4cSH6JaL5j1DshQiOMquPsJ6AXwM
YgrinakMIPf8EvW2NikLF8mZs6kj5D/Ck3nyFkyOz8ueevIfKbxSjjVzfZoImQrI
4d1Fy4Br+Z1c7588o59LdEgkvKGAl5R8P7swpodjbSE7xoTyvd9tMtNKng7fP5Zg
iofRrcCDczIf1wc31H9AZJ3OJb6+e/zMcHUPN55Z2/TrGa7IIuuZXukWvnP6Hqe2
NhOmksS9ehMoawraORhHcibUO9Q11X5TPv21/BotqH1iL7cNe19Yutn+X1aUxJ4d
wbvSzGLH1wnvW21xdBGFNAbzGmxWJPvug0JzvE5N5TYftjod9QoY/gJVFcm6II7P
Geea6F8NW/QAq359nzA7eB71fxl4RsV5nJ30Ll/5KOoQan99PYf4sixv/HYKIu2k
CWfEOq9XHREgD6hOj8RmnT2ykBxzvEOlmfCkFj6PsHnLhv/pKVYxQyQz+22Fa6eA
qdy9oLNevEQQdlpf32nd2ORImNuJ3MA8l24hV4/InYalSx3rJKZTJcUmGrFCfbjH
LRGH6LM7QOvzzEGRu0tJpnkfxJ4nhhLeq1Lz2/ObPh2uGT9XAou8rYkyuUjUF/Oh
wchn0V0rqgysbhCFJ2eWnvD/B3LxnbG67vHYRUHMP3pzdnXWXM38T7ds2Y1haznD
iThYSPoEkzglLdx0GU1CZLWwwhsDaQu8sKJ4XcGkjI7Td+bDds1m1fvdZ/VOOcTB
DAdgVYhwDuLftGLn7OG0LKXCklVSQkyZciVxmsJTtcSbcOlCYlodPS6zNyNjrrNr
QyRhpNm4OlqFIlk1i0DHIGpZgBfDUldt9wIK8qRSZyR8f9v/8ir4bptNQHr3HeQv
+RjRDHjqICyGKMnI2YZcE0y/g/EO/7fyLf4mSkQQsa09kg8YNRdwRvqt/VKV4365
Fpzeg+TZ3CCQ7qnqNCH/3w7/sWG+hKasc0TXGipxwhg0t4qAhbUs1H5MwaS50+/w
b1r8HrbdPHmfpQnP7Lkg5WFyIkaS+SOOH+Erszme9OIOeG8XKJx0fssvg5qmEpWG
bHMGwpWBj1Z+9tF3fIoLP4OXJVKD9URJG+f1QNmBgKqpqk8yeRVFqFqtR5q9wrYf
WfNB53+Y93myxaeJSITBoGIjyNTgViHynxygRCx4gEUXx59meG5rJNKkSm0WXW2v
PjNqhsbXS8zDPfCbpNRkYoI9TX8Icg217GooFGfEzz6HSYHHaGktaY/o2xtW+nfN
g/yM9R+U9xyxTc0bZLJX3PBzpWJ2qzXXLo/sda/MsfzhokNd6b2KXsyxOoiqZhb2
I9XnHCiFLChj/cQLrelLvuloELmcrdRXJas8+uQAotl9OFf6uwbYb2sQkv5C+yb/
ZRat225XpvKcaDwgydccCnaK+GrPhE3zIBM0FbwhIg0nnTLsMK+M4bzMMgLs2e93
J6CvkIrs0is+YNM4RuKsNmDreyL+dk4pEihG1QSZRr6jSUaDYOZQ2zEefJt0NXtC
6f6axatp8my8QtnCSv5UWPxsclb53woDAeXONUYy20egD2DrwCI0A+3KWDn8wFqH
YBnUrxGVL/jLcHoO26XrxgQAEZiZI16tvDd6UyJvTNPM4CcH9rCCFuVkDvkZQuLf
7Wg2TYejjytkHpHS9THbu1UZyQ1uFQk/GVa6yB9BxUYgzhlpDhxlNzExLsKY0DkG
DoPnhEO6YyXFA7laLX+WE4EdFaLaHEre/EIzM17nDJz9mMRrRxkV2nf+07RM3QzN
qhq2q1Lq0WN3bqfrtMMjNGlSko8qTRG/ion6Rz06eYXa+liWUCzwdrafsdV4QImW
mAgvCfuiENuuxSWhNpQQvr3OR1rD0+gX8YAKlSSWvMlErL8i+C8pOxhcDPLiQjbB
4O+DMwGD7PWGdshdn90pctkz9rWdkDQ/Et/EWie/EoEaPtKXYfDH322dfqirhHNR
MaM9wYOMMuofIwlBwwE3QyKpcp6akX4CW3gD/qTUvA9peZeKXA5yynX0hudw2q8F
OO/b21TFJEdVA6VsNL55Ev6gBsUbbaOePDbAXrL5DQwJtpP1yDPBPByzBRZytWY9
NBapYEJO9CKW8Gf0StICRkC41L+7CaZ/UUA3leAq/whBQWapjzvflFXbEq8O9N9A
MkUXgayFyLbvL24JXd4dA5KxyHlPfJ3aK4H5rNzNXLfFq/bL5vpbpJy4+Sy63fNm
x3Psi3uEU/ufNNhjFCQtgxW0DNEexEJrtZI3HS6mTNnZmvJlKi9Sd82rH606uTEC
RyXrTfziQDkcWvlTt29RrMoCusHnAmzO/CPYGaBsNPzj1KF31uyCHG+EuMs3FfEx
yq4QSubONUDqoba0zm5rCwX4fh0sn5g2wHsEUmtCDfkJjQ84COhFqoxMmIH71stn
S/FJtwP54TuBcxdSCAqTe1irIyVYtZye3ZvDx2j7jLTTajCoT89Tom+Xmrj1k1Dp
13bacUzBo9CVpzpXEsHLLidDB7rvgL3S4rTBQEiM0tFvYsu3jGNEx6qZORgWgcNb
0Wcl4usw9d2feRWqPue9tFo4NUEj32Xhmwo/k3mc0u7oixG9UXICE0z8xElQWRDG
TAiJAwF5aP++KImV8aBb1uldLlkRSuo0GIDAg9u1CXxJ6A4DqVjbUvIrmvR56EIW
zM5VH8ivyOHHcmmmwDcl1xfYqlvY9ssE52+9CkXyLKJFLaiWhkbZ5VY14h/cnr7A
WLzfoEEKcL+mdkki+4+l1NnagDbeXzChUgNeQ8FxDHGlXt+ibVJo4DHv+owUPzaH
r89EWFDLYsANQdIwoRhdRwceMF4sib8dEwmF6cpDbhsBhn698K8y+7F95PTdDTI1
5OlrkXfe6lj5RYENnUrRLlMLITMte6XQEzKgvfbicY5JHVHbOFqIm5/ewMu3OdPf
YcQkUY/CQhEwZc9HGSETfQWnahv36m5mPpFVsf2R0CGpbx/aDOgUVh57ROtWifEs
QSHWxJ9QOpGzF6oEiv+GPWwKtfh24pO8XhqfzAOJ03bcQmzUzFco5TpDkfvoT5gY
xtwKgvMZLvA1hJANmrM2rgOmVrNT7dX3BEDIIk0/Ee9Mg4CcAErsSJKhL3F4rlbn
B+lDKQaJUTcTiIW1fM72zUedJfOwVytiC+11d5aQzeZl/9Y6cEAN5nlx2eow4Aej
PJJ1nmOSnGT4bPbs0nkkM8/ZQuU+c8rTuqDCHqN5uaNn35ErU+T1qTx5ZYVx/zDp
YVkIyBMyRrjV2ouYDueP53hF96ujnSxxKkQJ7PMO3tCqEOs8JCTRk5/OzBVE9bm6
RK/ifT+ggYxDniq322l3X2NaxTbTxz0OvKYzIh3JuH33VRCUcSx5MMthsZncyJT/
dZW72Rp5ChE0qdssF1rLFFgvUuG2HPVWgvQcyQaEnUwYTgE5eANfPBhAs0nuRmqu
WEYGlhzEZ1kk5DpnnWv/W3DNfxFBZfRMbXSYYDoylaCnncZoe2bQUG8giEPWVMXI
1J//xOxL1MCJvuauYenF6qzIbXpKpniXlGPwk4Pok+U5X1hB/u1SlwpEl5e7qi7W
N2BtiXDTZF7nj5vonJvDopfER7GpCaE96d/be+TJ8Bi2eKjHvQWE12Ac2q6PNGno
WAfXPClJPLIHtPX7RGp79eZGCZkaVBK5laWly+wADUnl5ky0wpS12AclwGgtto++
biFRM6B92wJmLiw1Xn5TkS8PJQKKQGl8qc3jPXWb1YFgiZhJoE83lpmcEVrtNIS4
v0KnnE5JjNZPPZAluyO+w15rX9jRQXvc00CD9r0nB2pJb5vUGGvb/J0BBGFJcTdB
HBm5qCvLqoaGN75N9BVSpGUBEoYLb5TV7TSGxW8ihK4PIwqlc+ocOyCTYwJTnF7q
u+maOtqNgQp5pD4Iep+p6KEk/e2/KjRBDK710QhZarhQcB9cmVsY4wzgAOyF4aB1
7zJsyhuRm7DosvG2alVc8CfZNEJRELyxmMwm120ULyUuHejrfB73KAyve27rSY8G
yBd9BefH1bgN0pa+o1zFDJSyI2iNayOT+hoKOSmAHl1n0Aws5VNSrDf+ZpLqPmU2
ltG6/613WuwZusQ9QZ9MQyc/Ns5p0b6nEh10uSfVI2jeG8Xy2l6JLXnt9xcDUm1D
qYk+6YGY6s63iLLaPmmvGUBtobluBCAl1ZwVGInkDq7uzJ95wSQwPl5PXQLIjqVE
+Y4lEY4AmPZI2CEa3H8Kc2ZtHudXXacv4HX0nOJca/OzdeiBWjq2IXGZSo79UqPJ
GjAjHv7YWM5WkA6rs9O8tegI744UORygCv/3I1CuDrSTpBlw2nJ5CqPf7+Z9Lznn
Iin4lQAhy7XU2x/mxLJERtANBGDz05Swe3q20zfY3oVdciWz2231fBklrTwsvX2u
9et2ik2DJk203+TKnyj5NGlBxDWLXiD5KaVUWpvhCBTNQKpkaqD6wYTIgxE1vJgF
yaSdAa4X9BL41DQ6+bLKlFW16cEvNd5uCuqHlycs3P+iTSX16SkX6PVEY+GDkGCH
6Gq3tM1LpNWaZYRYbsGm6gElLsQ5F2JGN+kBF9uhsr6oisTGYz8we1qoWPiN1BqG
k3IlgBGF6ab7InvN9HGM87vrGXzzM39A6u1IZIhf7NVXAt4leNl30gbp1Rcib5s8
AiuNyGCNJO8w0wbLRkSRLGvYoGemAlq6ZPQy9lz7g5Ql5bAawpHObWYFSV7INxv+
f2jyhEc3NXJWKTPXPzfbvSOHhlD2D0kjTb41WKcc3BxQLtf1sZtSokpJQRcO2nWZ
YxmOBafGPi9WI6RBwwmB0+YD8GIWDa5U+K0mGn0gaLyvPqsHsTgiRrhYnTpjJVZY
tNm6I2rhZg9Yp+949jEsFATS2lc5eU7gqL68UIk4GRR8/ye6mcKrGzMMv1dyxYRY
PKThpAQxudTLVFwYfTMP1NVY+8fbP5ETDbE0CtNGpdZ2stXQ0WY8u9qeG49V1D7G
YIDV/KraLPlf7IyEfMX53kXhlAE8oPQgfDC6a7qU3JlXoU3T4WbNcLin3BH5Q0H8
aqeo1MgM8412Dc9ifwLevQyb2Z3vsBnGKrCLUaCXpl+lETqNCZ4Cxw+sx/QCm5lQ
LlL/xFpk3euNbxM87UsvcRGZc6U/ZtktnPRRAkVY+A2cJzuv2l3CP0O3eZ8+vz2y
Q92XgN2Xk1Vu6ismITVxn7apDy18Y7mEIEk6qkvCiF4+TewawFtKhev06fMgxJt+
SYfMwCeHpo/HN/rbh8W2jrhGUCzfIpVl4U8GqQjNovL5LgpvEBiOzeQA1J4iHbZZ
i0hFtEuMW+to6gb77qoMOrMSkkERVq/rlGyc9XKwNyZslZRG40IDyoQhXHID/kK/
G70tX2B4azXkX+Tkrylo0i/lRwKFF6VmUw4srVYG02Hl6SNJJXpfBxPemmaq69mc
3NyNQUl+eXdUfYiHVRJYgFF3mpdQelysjFYWWJh10wl5vu1Jyg+T+ZfNqbcub59o
I/mIcfomgTE55B1qeBkMk25Zuw2PWfgDZZmResv0X7Ooxtn5ijWbH/vdbseXUN0F
ow7M1+DzvarENmc8Pg7OoGTF3Pkvumyw3oNfRu8pJQB32EI/WKZg0/DuIH7WRl5G
R+Gy64DIhAiEeuW9nOpeHEFA8fM1mVkVhhwAewcznrB/9sF+5z+uo7/zxEUPgi45
T1WJK1UuRCJAHfzXh29+aNEpeNRZM5JhfWqCuDBfewKpCCHDKRLg4yvqqVe+/DvV
+wOjOkl7e78m60i04857oCnczvqt0rSJBEPihH0RNCOpGMc6ghIB1dooCzCLDOvj
i7/rENt3VkHAgjdDlPP424U8IHESQ8cZFrcapM5CTFAZpAmCrGOr0DiI0hwoB9VI
1C3iXVO/o1qQPNs+Zy+0PO4DJYKl3Pyu1yhgH7+JOJuLgDLkX2G0FaYYLgrcQ+4Z
wodQxkn60R2jSUbPtFe3AVHWCGig3trfwViMH12DKD///DzEpbKL38PF9TDoldUO
MIQyevTbSzIdVm8HocUb4RzRE89auXqc5LfHJgSm+1Q3Ic84J7iQFcGVvh1ghfUR
NO1E4ySD0/Txs2Eldn0vXuLrtFR9yjPyrRzKrP+1oi/9YruXOVpw3O9ckJovaPES
EXWBSagrp5gEO3WcV7KH4CC414Jj3qZI1nrYThuDwtbL+951/u4j/yxuMvNx7PUQ
MdOXCLf4NZP+IIOOLeBE0K4Pxn5glXACGrnaRPhoIxZhOQlLkmFxOvcDvYZqQ86a
ZcwZk6tr5U/not/bEGcbscswYk/nG16Ntzwq22EQMZD64mHKb03PLzAW5pDD0Yhr
OGbP2bz9TcxIQfm21kG7P2ghVk/+pLIYVzYYWogelanFesFDXTItOd0xIff598/p
E5z36hMo3V2RSMUUld2IqOKcr68HzmQNP8EcjvIWOG4bw+EziNEczUXo/89btiFo
805H63hao3ems43CH8z711k5UJ0bW7zEOhzgsTu1toml8J/EZaFwY2OAP+CQc0f6
nQgV8DGUDvCoaCD7D0JBfXFXoqGWSLvRnC1wj7C9z+XW1rPGVzrUdYzlEdanKK5H
yd+XJoNoaUwy1WzJdInvdC6QZRRdpx23zsEQwGWJZ2YMMaolardcOTwUjiOn4d/D
/08zWe6H2xOjdQ9hvcTcRTV2iiOWKPtyh9v1+d0LpoGjoaDF6YZKssCsfbl7bzCX
kfombOz1hxgdOj1wOzsOP/7n5EarYkhbJa0303WKpktwz5bXH4Fd4rCs4+nWvjWR
gmp3uXxshGj029yfghotX1Eyg86CLQEpXbRuT2LY6ibHWQipBntdC4NShdNzku4K
DiLKrfS5hd/xGLRdIHEZLh6nWQZ0OgCjYUetP9qkHxE/NFcbzpV/B1TKXw9Avh6a
4iLWOj96jSfFhK7wVetFanG0rN++2ulHmtX/ageMzk/SxbuLdgvg2qqpkI28BCQb
mnxyCOwcYwHCfIyVoqmxXWe0loCtEsDokl2TfXc5z4mIHatIFzhdY3m2T231NVw2
7olr+VBFAf+MvN9dUMOhvnhq4Wf/oKz+qxKzmSYV5FmC+V/XOq8RCG6ICfJEXPXV
QV4818ez4zc+9whzqyK5yN4PMlWqh2DyaH6ZkOtEl2Dt0lsrK52xruIHyJ3OhlJd
vuwLSQ+pLRiujNpGG/UDM6IdkqYeLN8M4C3c3VGZaKpMHBSMKkq73H8oY+02K8ZA
CNxTv0CtafxUc6pED0yU6Pv1AIqlroOTSZDSJgJk8jTFioZzZ+zZ4al+aF9vM5S3
aZyN4GKG9k/eMk3KZ2VL+iFmv2TxCXFSnKnCXJv7sL/cKDcKPEnX1zmO3a2ApQmR
FrEz3yyJs5nT9ek4WWCx7LYB4C9XBzBYqStJouql8GnihvJC1zBuyajvw6dy5CeY
pcdpYBiVAH01fAUrk18COF1kIowhOzXz+puAKcoTzDV8FZ62u5DPVTDmI9A4YxKj
Tib2QrzmZvoeMlCaVmCA4BwtTktxi8FPWWK+74DsXmhyouEC1EP96IXPePNpaf9H
kp00koKBXfwqBTdlNlTZNVj/2GUmgz3tDkEqAYCeYdmE+AXeML788wJIeQuZ31ou
VmXe8K4ImSe2dn5kBiWyB10jCwMidIgAziQ7qdI4Rouq7H7H6smuN+0EwFee6rTO
lwiKvCAdb9kS8VHir6iJMa8Q3n9NbHLhI53j4EXMh4t/LrOXzparFg9nR3g8Flan
0bgRNv+wRLtH0LOgUTfaqT7moWmW0hNCJCUY9ut5TfrKvsP9qtb5lodr/72q1HM6
elS8PCBMdPKTJo/Dcl0LG74VKlDmtYRaG/aBTet2aYcvE5yVATPpm7IkARGKEPNP
o+MBccQEsaI9kKcrWrJ429cuclUCsq+3kKTMkHQMicbB/kbwENIZfms+SKvpgPt6
Bx3p7lqrfFxlEqY+ghKXw9+eNdDF6EqU4+8sorccqkuSSbubUN4LEWKN1FKfB0H/
fMHSwiwdqzDwhGNFESvCDjobgLZ1GMemcp0AKImBWffDTnOlgDVJCJtbHkQK4+oe
X3FXVXtz9eURPItxczNF1RD70t5x8fLLjgLy9aG3B1XABwnETni09tr75aHvbYz/
b3mkhdKvdZR4zD4u1agZnTeItqxpZkcA7cubuFTKeH3s4m/fDEsShAq/wO1UhMCo
wkNmZuYNU8I4GcBu7JeBGxY757EkBDFKfqJNSSqM9J454WwwO73YEBKRjLoIbYec
+nTtTs2vpPxbAmVYAiFsuAUGhdA4Iq5sJY6UVy/3F1h9xhdEm/rXI88oIMbt/qYH
RxWqouIL7lOhraU26xZArk2gHNzxk88OllH7q4IOE+uw/a9ZtNAcfkp5ohKS+rTn
K3BjaeyYFCWNs/vGCNIGVV6jUhueOZ58GDOfAdPFFoFkUNTq5dbTjwKBBnRkX9XQ
Nvf1P8wHLqdki7QJC9Mrwi0DKGjYy/Y6GvVkn4tkP1i+XbT62QIBmqMSpYmPqo0i
atUcNvvSjycTUkR/QlLTWiPAPiAiVMH/IHdCYdR/ezhp1ChypV68N5s7JxgNPqQI
gi6QY/UkRt0sAbLYnAbCr5HA1UN3wxfrvj8Of9Yi62avWRU4dkogNvESIKdCSDIK
iA08ngAwzRw95i+XUhQkCTVf7z4Z1lGN+Ok9kWf1oBB3Xi1Wgw/rAqahl3H4/7r3
s6XMVsZHFC/DxdPeibstDlLRjGrYisFxw0/xsX1ux9XTuLUi4EO7DhFZ3ZRqmNSc
pzW0T4wxMclJzLhZYKqutEhyIrQGoK+C2d1DX+Pv60JNW1xEas/t4Z3WDLEZouKZ
Rdv7oko0QUVcdtxvBdjJCwdt/+Xu/Jc5vG8QvhS4hV/SAQ2mlHJMv6iK4tlSiVqf
Hbml7oMFr90UM+SHNwn5UC9gGF9aC4rpcqYbxsrwOGjzHUoxymQqPl/EN9P/D7+R
bjvNKg97GrMsM7AmZWRN6EYNv/10IxECExVYR6yutatyf35n7NzL9BubA6723exs
xudng1xb5AX/iWN3uk+fqcywNwgBeg3zKEuKrqsyeSIw+9sN4LfU8ELFrGG7f58M
YSIHJDNHFW66+iNVxD+SrmOrmpagJx3gGykqQEEVUYJByhvDpVVY6MJ8A4xYQA2b
64s5AHdrOOAjlGw7v7tMnvZXI6oUtGaSXzN5RJY+dYHcVKO73BMJMvxwcujwVLZx
8duBRyb6yNXPuccBiYunnARix2gFHO06hwVgjq6KLditpm9OrVPbzLMhA1LJjmKG
8SNNDPTCIBv6+eigPHqPDCcXPIcjAJT/FI/VpHUizBv5B/KOJ7Sf7ZkKDC7rVSiE
Q8jwoZ+IJweSL/4yihMwBv+Gl8EkgaqLr7jTeye/0wYuxnV9XgCcS/Xs5SAfb8h3
sndtYZhT+dhHXqvPZDVbhzRRG6PWzCGfmNSNrzhOR3IeIyFzEk96yZnBCOI2z0XE
IPirF4z+4xQ8It1F/b3hS2ypvwl0CAsmFczgeippQ268lMFdoFsCrZeb+XMO4x7Q
uNsMQ8CdkXtRLhTSNUVEfpWeUxPKO3eBAUWfT6vdouwdAO0MgnXvsXEBXCZTWXlu
zjfg50szNePx3zY/zjYZoRRXRbsSOLdAqcYjvg7W8aIk5KIfFxBDeczDqRYGhNhG
pNcgVsbLCvEDqWcRUcKEXioLMlmqAxbiEBfzIbLgobNyWMqFn2rfVQEeBeoupY8f
pqvr7SSTNrCPLyXr841Pfr8kLw/vbte1Xt3VdVH0F/+S34a8eQ39q0qHTwn0MzAw
Jd3ai0oGrGkI4pg4SYcCoCzivvXcBgOnc7jLkKRLmLMy8PucRNFQUAcaM9GT/Cdx
OhNSflzGXLrZB+1ZQKD3BlWUHD+1h+u2xbPahYsyNZSPWm5c/czouU7+2a000Zls
ckfhdBG7CwdS2BFgTimI91/CGfS3IhzB/gTFkNDTY1wCcb8ioAqEBwHkxbaWsQGX
H3KNvEl88jMuNjHJAwkaYtTHPKeeUBKjrk9uq1HdlvvjuEeeiNKMpN/FW+TOtxJE
qJUM+dLay6Nb5nnRNYTB14WG80DjBgdAlT07ICAc6KYy8lLAOTLdGiUFH2L3HMkT
BA73RpXwW6KIRmaHx4z0QU1KV2BBokPy+SYFOK/flosUy9AufCrctXXpVUXbs6S5
ssQ3aZyP0SnMTKa1ymFyB0IgxF0Qee5DnT7/b0NhVEwNZzq4tOLvGKvlmvYeH7OA
nYFj4uF8n2AyS/1RvEqkZ60Uy8lnvpSofS0vIs7+f2J9MRnS6HSEy5pm5OjkUdgQ
5mRjSzAPr+AyJH9Jv6kr7dHxyiJKMegL2I1RTuqLKgI6qg2OjLLWUX5Am7y0gE8w
xQmNTbKc2r69T/XEXRjDI9vGUajEvnXUXTBNc4Ly3QTDo+PFNLQKeqZdp1yRAn2h
lWxRlrST0Cw3gnBaS0oda27EePVc6VmVdq+/9Q4dWbPj1jgYH18yRgyBkN2yr6Sd
JsGtnys5jy6aT4Wz72YCgcJxna/mzkGzPQH0PCl+wO1+V4aZb41xJhhWcgpA3Idv
pRnNa3gOrPnzdg8QIjkRagP3dbRFFr3iFVaa0jpEsMM0jxoA9MMwcqHM2uZbib8B
2zRBwNGL86BKWbufK2sG99p89lC6cxuLxOk+YHY5y+5wV4aMGRu8xm8GY2QPZVtO
U7tqi26KT03KKOzhRaq4WVvhTYmt73fPS8XX55JZF/QuvAiS4NfM6GDAhWDxIWHz
TxnYctqYUGT9lGDSkpS3XAadAo4lhTniqzHgfK+65oThzSruL8h2DPjRuPNSJ5i4
NtIOTm4c8nY7j/QcnTIwkvrP9FIF6DA5VcGOPY113ejhiHqPDrmIDHfEBr2TPyjo
OVtfpnyqs517GkC/VkvZcjU5Dd+fwD4dSOV7zQHtl1QxFOT5kTxlVBBExvsMW3B4
/QJx282tftmAWAcXhY2vv+5DpGjvwd5qZt7Z2CFdJAR7Jk00DUvjjSyYFcudW5jW
oaa9iy1blgsVFW0IcH9ze5v3bG0xTPK3yJxb65Su5kEYlKZswrkY6gcOFSDS3yhY
RYZt2SYt4Gh+ZaWKbMVw66gxn0VCyM3Au5d19EV60t/xHT9GfuqRW+gKhi+DYGyN
jWJk1uK7GLKIgD1cPaO4/GmMA2PbHCbHRRjcd1ga4quywQajDJH/OgZvre0rCwco
R02POIheE2p6SgEHCea96dkhnTV/LvfxxYj3JA+J5hOSpeCVC3ROCtHABl4p1xJg
CxdmIzXcqLktzvZ2BAn+tJOpCgfCqixnr/83ib63QFuIFbM+Br8zwcQrXZmTVHJ/
cdtWstfrK1OOT5qo3Z+QPIfco9k2ndC8RwMCWgjfuEyJZsXMa2ZTbKuTtXrZ3mJf
HkVeNz4ibXn73/QIO9HwyZWeKimCLt9eQEhJQ+qRxz8hb6ADzzjy6POcwY4UVga4
NLmyt/1ObFr0Mn9Ijjgo6YBg4/Fpubmu1odgCayLzgagt3qw9w8zdL6MFKixx/OA
LbM/UHKQVs16uzz0KjOYRlJNj5phxT2nTcoXpBkg4YBV6cr4Q58+AcKkyTGr+H9i
5kNwUBlq6dgC8PqufUNzEnrfH5O8ixle//zm+r26O2pigkIFJio70PQSow2BikgY
ZOWnHyyyEa4SnkzqcZ9Pbisqr3l5cYCP8G1gAsTTTEMRA4XI0IgJTu72gCU51Phz
jmwJK6AjoGCgnBCSS2u6gZlM1U6tzOIldZp3IUplYPtIeIxBm3WZMotZzKd2IlGq
W2aTqMCkUspg73eAF4tHjqsH5QHZojaukrxlbYbvkI0x76yu95NL1QKVVLo3Ll63
VK5Aj76mPZscL4g8b/IL9ryPWJ5A3yQJh8E9xI7F7Ma8aXawJGKlDcDKSRVzGkQm
Vbcg8tWBjez6eRyl81tjjV8vsWahfznYwIkHfZBGvJu3ynNRNV4yjkB/orXZohwR
zHVagRBhOZvDYuwlxKTLuCd3N6OgQ6tqAeeoQ9+PG8zkLL6lVDPB2MC8rrW0f02f
irzM68NNVtY8XP4dvpWIg74Ico7DzG64Qqpv5ShaHQFL8/wS3Vu+C+fZPwEEtNAG
Dl3PLwMOpwuB9ozF2flGJ38vfQGPBxq5DVLaQAT7sKkAakTHElQwHA/PryDN81x9
r1LazoHSQqJTjSWcdI3okhHa4ChegGU70LCqWMlolSKy++V7/rnIzulyDD+dfmTF
udlIF2BmprnB7uLcqy6LXFFebiWDdJ8eSVd8LWgDJiN5fVoHbjWsvwCJgsjoSuOa
OFdEUvZpW1vENTWYRq+a/PTjM7ZBywdvUL8G9IpvIK2t3g+MHVJmhrLZljSAsE75
lPJ/N06CSweHv7aANBQmR+ujAi60ZoDSRxHP6Hati2q1D34GtmUs12q/Bax3LMyp
Yc+T/Z6d0V35+D+p42dwMwhM1NcMCK8yQ3BMlUfjrqXSSvnj+/EjPa9UsqDZkOHg
NMFbcwXLwr/1gCSvucu4hBMS/v+7Thn40+Nb8ji3Fd/+429E1gOJlX78eiqIkRjA
0uF70FPbAtFS918xrwIZZ/0qylcF2ho8NYmXAHUZsJwGxphZHE9YeDooosbnNprN
mt0Qy04r4wGgDcTCra1Tux8fFdHsNmu/oJYaPk/O5TrCLHvEyI2Jk2Kk7EtoZXnb
nUpPYuiIHdEOk1snTP84FkQiSx1uIaeemwLgA/Uxw7N4yMs8EUYpeuZYMIPcFqxy
VPwuLOQHTHhJR2Kxg81dQRPZNUoM6Taq+/R33I6WOQAlD+4iCTYnlkv8G1MdIt9P
0qdszw7ZeC1D8tcqtjAKYTP2P1FsJv5D6841TUwPphVx6+pv/+g9aMW0J8JbnpjI
xXUpKLXccDqiVhkw04ewoWCi90pP5IooXRBgdP1sTj/NnZqR7E5xlR9fiLYweA3p
8WkBfgiA0g357TLKHYHixb3QQl/Vb5TxYBiXXldgps5dlLBGIdIn5zl+2qIUuEp2
/xEnA61RADwy1IwZWKcY3Ha3HvC+u52oGeOoFXCCkgW+ftkGYEoKtn7gFVz2Cj1D
3U/E4KTOMhYF72itD0ZjAERY7/RO5VFByvzrToYiedi219dBb9Rm1++41crsKx94
pYHHmVX2E2feNtUMSdXQIPD5ILH3+HIxwQwBfdYVrsK6u1ZbYdHEtNMNg0f+FhmI
h0Evse2Wpba51N1QZfFaL7lvVkKh8c98cCqu4dEM6HvFS7wX84WSfVLWxBNbipyO
SeuWiso0kLw0+K+bcvHNlHQelI4ZUBqZAWBEobqyyeOcLkiRQQ0Cgo0i5JRHf7y1
lE0Rsb6KBha/htn8ZMKuYxSsacycoyETg31iIedgRmLzOdMT9r4XVF532zDsXVYI
sf3d5jnIiHzCydFr1f0Lq3TSOuVsNv/LGa/KCRNGq583Iw5MyiE3G3U5r2yUFcmT
DPzp/RogidA8Z/Bl2iAp+BYcM0cdB/GuL0uHcJ/CFQqhyUGZVByUR4ADiGYAYgvs
YU851omxmMbJEUjExTbH3bAcWtoknbyH7/RRrxb8CCRR7/BFvIFeQGS9RwgpyG9g
o/OCJQhaozGO5Lipr+jX+1X5GezFlvIdXjnFARpE5i5K6rBPMn70L5/VID/Aj0xr
jcmkbsKC3TYkOJCxpKKMKmvXLxXxgA+teJRyP5Uk1OS3YjmUsYbfuhMYGgZlOWmf
tJNwwLFBOoVSvnuiPj0jbxlagfE7g9ZLTvnISbJMcMmu2OpsfWS1VyAp6jw0gtEd
dA9s1YGcCF4bf7VfRpKZrQlO0eajNaTRVIhQNszPenUfESSG/qwsZz0SmMV1gqk/
U5EVUTlpwZEmyeIQrS9RViUoHylvh3ROhDIJJFwrb6q/oQKj+Qzzzeq6gSdQadY7
RiKo+Qo0y4m2baVeoDB8F4CnMFGL+iyRIa+W/O7fGwBzWRPdeBRkV2eKsx7G/Av3
Co5FrnxnAgrKY+vIk1WqvjNTckQ3lT8/5FJ7b0hcJUBXtf7otHsx9y2ARAY2Ose/
PlnimZWJs3k8U4Z94cMfevN9OrBRBe9oQH1mrMVeR9mPnc0pC0+HhdSc9ydjzERF
G68qNPfpAwcQmLVUHNWR7IXltuCr9awpj+s/J+IleUCV+oHr8atn0i63l/hQ4JzR
1Cmg8UV8rLaPL8UrT2QWm5PGCZKgVAS55GQaHBDxswa0tn8yZZRYFSGDraiAADYG
R/gWq70IgHV+aOKqMQ+3mm45RFPBCub/cytGAhP+bqUdeFGaL64BOzB2m8UTlcGd
v2rWqgT8soH7Fnp4W4Zi1ldF5SNatqX0f1HW/5or0VnFIxmNqgLBjDg1odvU/UWZ
NhomS9NlEIBWXLyC3b2ArHIcbnAu9u62XpNWtPiTsb5b+VYvuUAZxKahxCxGxLFh
fDqnEBXW10pX6CbbqawnTdPaEOYfgLbLo0DRPuW+cN79g6/XjBrzN/KGpublQqNN
n1LWASYESsRT6QYvd/BDfgiG0NJBAQyb0o4/wjGlAXiHzsgKEZuFWTu7gKosXbUA
GPbYkYrPd9zHNTh7HOadqZ79dE/PtrHO4mQ6E9HQaky+IijGgfsQKPS+3PM/7Ywz
7eNzMPsAew6EaPydrfyLyINsPTbMWIY5SV4M5zbGVii1hcnlrvmsBrs5yXvCrUHf
m4DEaJP8CfSEUfUD11gqYXG+caKBoCdPqAZJdcyW7JvIXsYl3AHwl+rAJKfQ8C2q
C3FBntXErNKDIBHYnJ28lbm4INml1CiToPak2X+wZejIxafT82jg/xbNnxCRIMWv
FSmCuWBRK9F5plOQsBeTvvOLVqoQhvRSh3vSoNpZHLEOukZ4YNkOkG7V6X5cXhYK
wt2W7ZtuYfT3A1GescDBcdkhwM+igmwhH+h05rnf+V/F4IpPOn/WY9AyORG+ul6S
X0dssBDbRPJt84LZtFGq8S9RvT0xPXqsV5og/iZMFQ27h4wH0O9VMuNnykpK6uSl
LDqtTUUMGj6IcgoqiMaMeZNMYO7Sdn1oWyrMBDPAzvCi9DEMzyAoESmf9VgmyV5y
hWRcr0QxsVk3PXHH9fWg+B15aJFiHhiZ/wdDq00kPs8bQl/yyHJOgYMYpuv5rQT/
sAz/YFO1M22JPxpGcX7J5ByILXp5EHQymI6wc/FGky/t0BL6gCeyWZ1Gho+oOAXT
b5/u7gHz7C5dqSwTVkNLm4MnChyEqAkYSPzDi8BbrpZq2a6npsrth3T+mx7OBFNJ
HjZ+jUJvnW9CXhP7syNhkTwY84ZWPuAV9mfDhIYgtcWquEj3RBPv5XvE5969hSxK
ZdV9ZKJGXvIHT26GgHT+nvdz1K8YN3KjHlEtmUpGykTsGv5dF+rlFXlR1X2l6s3V
OQpe3gfkAmAnAvGswLVyzcCkt4eQusKm91ESGnpBoKTolV1lNQWKoijPu+7VUwEP
n6OThPQKg03b9JZwcSak1GwwdTSCoNlFENNipAQeq6Fg4FXL0BXtRA8b7ccm5LYr
nG0E5G8y20zSMA9CS8ZCS3rRGXGlek39iKpvb5ifM/J89o5lWkHs+EiRlsTFWdCo
KXSyr2mbrI9cLAI4Um/0KugqAfAsmD4HNNe+Od3a9ceYFKGAv1ZzjV3BXmFlcOzJ
ASBG+BgU0ttO3xndllluEieLNNoROxZtjMxkRv5Jivoht0OL+w5eypplzMT07ygg
UpCOfTtAOiqyhsKIOJesIidLRW0kC7hPsOXL4wZF1TyKxsbDZ6z+UPzWRZ2SUPlj
ISmF3x6iYiHbpPT20Lvn/ucYIbsE4NEMvN7byyTlfrsP3ytWozLRpTnZPssI27m7
eb9o5HQi5NOD2sOAZWcKQ8rApPAKf9BXipIr/3LvdlJEGvstQZAwUFs2+nRnes1d
6EbqwSNYXynPHTlPKky0WvPh45mVwXyy5G78b3aGEnHfCk0JQ2nOXjpX3/hSZO/X
lOADqkcmH+NeZd7y65FqHn1LNNp8jetoMUZr3G83ja6FrJ9j+kL7rJGgn6OA1hPt
1y4r+ulS6J3ZQnWkWlrTTz61r9oTnc9ScQmkvCt5wIbU/jwq9ipi6iN3g0aaQ1nl
mRDVGijBKhQrgyrEiJz/gg9gRHzuQT6+7YHYmeACYWW30+lh53xTfZB+yovAYO6o
HxXUIdiaVeg9nsHPi7nRUtXMtirgLQzevbGMfQTFaDn1+HnxlOvaKzgDOoZ168Y8
CJB7wpHYFk+Mpoagd+DHrnQzXpfaUXrL6KJHlxmZzzT8Pug8nilnNqNy7PduZjXj
eqVGdRrX2OQZkxyqxzbGohGq/OBNUrEepHgkBNN3DWa8Uu28WH8cbC+D5lAJILWV
7rUxA9uMoYfXcJTCwLKINMvKylQBmqi9zfeBo38QLn3vFdiPqjvkFpxJo9jDjinx
zu7FMCduxDhLBkd9/BDfMMCWUoL+b+rRF0Gxd5Z069LW23dsGvEpxMl4ZiXwgTn9
y629qLyy1+5E9VmQBUp/pNI3jjj1ptdLP2wQ+XGHg3an/7VP19gBMKuNBCajGxBq
0J03GhGrGzRHlO3BM//M/AxxABncmwQ/zm3y0Vfsrs5HxSiXR6IVaEybVJpv8w6V
g/nNrtIuigqdqe6bebTTVUyetn/Qe0whverUFbqhxt/M/kMRXxtt+JimGhAtVDcX
FMT8PRbUf10WHwbOsmDCU/QGfcTC063xfOcL3xdzvLAOsnDao7xOUh5dMnXWthqn
krBSW/EgGQwSktCGP0NdPWsiHo/zjAZ0+T5x65Mefxpa37xpvVZYufijNRqhB+oU
pOBdLrwVEBaZWaBtPypF1heUMZM+WFxBcYKvqP/g/Tr7k6UJdFfjYgQjH+JqdM7q
ZEbJSONLW5oeRtf3UK8XO80GY7KUKe2sBjKAmzJF3J+Zk/j3znhkodFPRt/Nazky
DTN0TT7v6UL60CjSJGz56M7WpvmmdzC1xG5jG9nSYgjuyUIQB7n/gZ+0ic5NvNtY
rHIPkIfNNUjjh6cdeP5lpeYVPq3xTp+v/k3O1UJm/L22cUnnjc2DMZIk+eyW9/22
mgugRN7/R2MolwVCpZzo2D3igkcFCm/yNCCIeMk/fjy+U1QlBxDmI7xMeFJtFOOY
CxMY+4MZ5p+AlL5gq+jNTLrOKL5hpZtCsWyXW3TuLQZPbYhP+u7Ss76wGtYlqniF
3k24bqP5BvH+QwjDpRDlCYXc5JONQCqXlriSAWfPODsFwY9Q0iM+vlM2U0FvBA1W
3Azz4neQEnwhsEB5FSlM1Tf8d9hcclORPQxkVw2xf/3aFTSWLcsxiZR3ZFyamlt9
wYJZSPK6mRso9b934ry8nTyiq932gAEGsVFsafWRQ7IylKTHeh/63TqI1K88GB7H
X2b0i4DvdlsBDvGGACoAwgDe4pAibszlnDDI1a2v5DpLW7KPCq4xCWZpD+SisI7a
pEJEpP43rB4wt3WO09xvPE5vsdzATZAqHhQ8ZfsIeGtKT4nrXceVtAQc/614yX5W
EwRsCShOKVyInSLrwA/i0XW8mTwXfXVTmAL4ncg15wYwv3Wq2ZwsJMutM930cfip
RqI3EQ0KcXLut8ny8lZWyA+n17M0IRNmAWMwwJSlvFm8dJDxUgzuUUMv9ljSzLLo
xZbAofvJJGi4GA+5pnlNMHRC2RgaN2WYQK51LvmncWhMkgAjjgW+1+29+uGKCinP
rUDvZU0WO7Hcj/9kuUu7dUVbt7UwFP1fhexwn4hfBaJjhNaTm60eZv2mmRH0LnCb
L7SoGNXeGgzYNvSLvtoE1bZbUXBlapbtT+Wntb8KCtFai0yC0sPWLk9V5mUcunOo
6kToiLXnn3FLGAfOBLULHYxvKHpZLqIcbwu+BcTJyiuO2AXqpzaDi43Xq8quHT4Z
xm//JVNdDpEH8UwjzIY6FShLtL7IzpReGT2X2EWPy/heA+E5HEkNWaTTXyS6Po9v
D9nk9v8GPhVrk6PsB0LVD/HIENDfeIxUBBKq+9bQiDswizCAk8pzsB2XM+1mfoFS
PbVNYPvv85ew6GE6khqWcTPGIic6W9/Cd5BRJWZdcGdNlYndDktoHV9kP11lz9Bt
t3oNyv5qf3inyzf1K/Wkfv4PWUVZgTqGImy5+1MRQkfccdoiHqfM1RPkOJ2zvuD6
jbeNmLc6cFq5nY5P1E0j14BjG6Gwn37gsIl8mgM6W9bbmAYhdU0ttcKRgEP1gX/n
pcnapaXEvFSL3qcsKM/Hq4RNu4Lpy1WlL8m7Bhc3f9Y0dqPPXOlkXwXZecMM1b1u
PFjV2zybwdwp7zDKuOmgtbYKuCkMCMXkM4MOSP3i0fqE/UmFTDptbRbYGOZS0Qkf
sDM2Mu8nfNxIvJNZAI29jvZS7bqZT0eG9V4XXDylga3J1SBWLHD3GV9pRmlsAiwL
O8UaBFdnnzTJcmHLgs3kuSog/X2effLVMWcKOk+qb4R142yXeGIfky4+JQN7YFWv
lW86JWZITfXEND8/DB2XgKHXgr2Jg7NrsG2bgq6E8nbfpcQASEeYRielWlvcgeMB
DJiug6Ek6PK0Irp+imR1cOKlb3RkBI+pq7mVLJrhkMSkmVNtyZvY3GaRHcdBth6s
mzGpCROMkXFDPUQPcwPheBxE554iwfJDjDgo9gOXJXrwro+zvVKMe4drs2jL2QLE
7GYm/Uy+++OMEoCwwUYQIK+8d9cjhjaLFc1skrWscj92bg7hHH1IyJ49gDzsLCch
gTu4a0yGo8mvTsDWaC0lfSRZRNL9PGLhh6SFzq9RIP3acswvFdAg2Sl8RjRWrBsh
la386asdzILY/QOcEj+1n+YnwBX4Ov7nufPG9qpj4AwHptzlxbfsUF6upXPDhePl
W+G4ZK2oVPwm2GiiSMOMFeQeyYyFGNDkZeJ3Htm0u92fRxB7/TU7FuBh7yarBk5s
xE7bsbVL7GWynzm2H4su4CZBiQwutv69NstyOCOrtCusI0G6Hvv+174r7yunlyCP
9SBXAXss/2TLHM8GHNTFrLRUvLL7dVFk6BtUJSLTWHFFGfhgGAiHCyP9bdNopwtQ
VBdxCRJhGON5G5cYvAYAjfMhsWAmw8Ovt8u0hQQ//5WFndpew73kFppT6TcQHR4y
oV85JXTUuiFPZV/n3Nz225enAsj7yPYqBrzAl/gIAymbjzRiTm/xEdkf2Y+VLSl2
zW4bKTMuinMoL+ZChogwhOEvsDXTBtuaQ44n+dAUI4o/KJWg+iKbFWFlZeN13Bfa
6SOppwHKM+dxAxxIh6g4QRpOycJWyGQpOVmpVDYTvVkS6FrtfplcPc1hWeP5wuYi
RAOLTSmNc8c7Qq0qHqX21NrDim8moKrn4PZ6YKqBNgXVnISx2dbPAXDW40pTYPmH
aMnNSfosgN9Dkw3nb7Gwh2KLfXKgYf2uS6w8nZjtqwSzqQhHZbl/iHwsZB13qL0W
MU8kzDUcG/mzH9COogj3K6MJ8zVHDGreeqfeCzxXN615aFz6iuf2NTHodK7ZTOtn
JljvkVDNfMBA7dnw0fUbJKs9Rcanoffgm+xqBAympE+PufIKMfKeCRObgoVltmgc
VFxc/TT4WCdgjhQ7TEjkXEm2WBvPCixFeYWgQgEDV0Rx1L7GswePgc+0EzCqM6Ui
cgzP/TYD0DhlMkD6/o3hoKJTgGqcS3cU62CUvH0HgxtT/5mlpzICkKJk7Ui3XOzU
GWiFh3bcfZd3Uf11rcRuSRQahg+KoetnXhhsdJZY9Tz+eZQAL19HVxN///zQz7jT
nXz245KotJ/ED7fGUvxSUrzSlf+b7j362q15h2fKmxyedv1QfEDPw8do/G79CUkg
C78wmOSN3aT7HYG+hwmZhwf5aka5fLYGuNIdyNECGJwoKEm3l3EJjsRlXGunQKbP
A1Z8bzEvakgRj2qF8Zjqej/LaL+d0fh46TRAtYJStEq2MokF27tI/c1x2mrAuS6l
dWc6gcpklubNTVA2N2x46/Qs9kxwhHZfn12wJgJhZsfqVrul3rAnqkKlelNUjUn7
OVcUFBUHRi3hr4+wlllusGsmlKkd+PGG185gVq2epNPrhlgs+a32V0OCp0GPnpFz
4Y2dlXRH/bw3uQRMCbdBRVl8m32IxhYzgDwuFrAW/oPu/6VkkXj6UCc3qZu+eoof
kYGZNPBYHWSWum1fRS+rwWuROdZRwYTR+egIBTzuMAaMnfokFb80T00YyY/nkEGS
J63gX+muKYJaDUhDbK3aZ8P40jfyouQsjJiw9xECKHgROK8lKHtfIrKagu4hPd8t
LRXEDPvUbiVaQhoQaV2pvwGN9wcQZz6AKkT1I14WH3JQgRRMpfDyB+oEghlOv7Ch
AgKHOFaDd/ahmWXZjH+DxEYj97DrY835dbjN+c2YjrFD5XezbfMdtIxow8b+SuUF
tfsOLCGc+2+dYV14D4Ju5UFsGFwEyf7mtx4lXVvcbXFD87uYR0iT+QxUkk6dOiOZ
AGTu6R8c20/FxoJa87jgtZtME2AAbVyWQV2ozxWyjnrCsUzfFIRUpuKM9yfKjveK
xZgLYOQDQq8dIAfXAhGX7MfkTmji505AeyjDyKXAoZEa1GBIC+XRzYKFx63ovjeN
Y9cGD8NNMYM9jAudxaRmZrtJyN2IIoVgQ8uYuCApiXlp3sbO/h8OKFyQqot+Y2pV
P2kGRdw5vZuSBhtRDIcJt09plFa4uTcRhlFxV1rnGPSlswPtdgZ4Wj5CRqxnk2Tt
doq13o6LK0gj0EIc1dPAISLkdRrrrsjs9TcwiDCTIOlTQfnzVwPVJG7XtV5OBxoG
nHA4Po+a0+rKSOy7bIiu73cpFambJ46oeDexjTkMx95kEuidS8bPX7Bs4vbFNIGW
x0BZdNUxTij3O5qPjNX1jEDUWSIwgJ2dInTXEv/jldKzTY6a34UIJgGePF1qszHF
9cgNUlLauhg9JMBGBp9+qYNWs4FHYjwwBY7MVKyrZLXP7/neQlqW5JJ+xzPZqtkS
JQBlplPrm4SXhmWLD7KqaT38Nchl5UoGlyW6xNlxyME51z1YHheA+zAXvBYyROxG
cA1Blv90GHm3cgHwKIwL8iKyCmR/VXFl8Sb9Bbadu0Cznzn8k/+EwCP3WbrZCPtt
bexBNaHgU20FQs1CK03c0gjJQ6eCeQZ/+4lA4tUVBGtfYqPLYhExxTZfwIeMi2Uh
AgMLfgAJIsrD99RGC3S4KOQi7Xs0rcJUQzInItSH+kLIxxBji2N11llETU/nSjjx
i/SrKQ5JvMSJfKoVYY6Ce/9FmRuS/KRyvouxjA4uTEGR1koCpcwhvAHGDmv5VTDM
dNkG+HGoFsldR/nWIlUdsnyHbQgUZrxtEhqvIXZYQ9C+f7j78m/1VXiK2EPHa7MY
FZh15jYgxbaclNz2ISTgPEWUg7p5UxnaywpLBBr4X7n/SvWMYlf2KsUzbcsFcsWC
pPxJcLuFO8NCNRHQVimgrVNZpb+LIyHW089vd5UL6q79V5luK0upOiSeuEBOG06M
pSL1Od9wqlSyzPGBLpKeMD8m1YFtNiEE+SQXEyWxZbWuEo7xoSvSSjysw8WQaVI0
Ff7LoxMeITZaI7sUsjnIj2HpSlvsThjM/x4aqukh/Flpp+MpM80QQ33UEu+hP2dt
E3uZJ4OJ6w0Kb5T0lohgp9gqiHcgyT+D/JaIms0BFVtEl5vo7peUZOz8+VtG8Cnl
iYZ63s+6ToXWWdVhQXR2QJlfHUXKuzfMQczSNoYdnvlP0mCrM6e/GigawiADMcO0
ohJdFhKeOfWd9hvLBUz51ZRUdzjj/a7BIPQjogm51c3MSKJSIHtwkaoLNeJktt7k
n6f0faOIJABOCJXYwqxQNBMu+8P3AI4Dgeqwmr4bJWDmTM386lqh8GnJ1f/F9NUb
W59rxF1EvzAmOMt+OnA9E9otQQ742BZEPuP8h8F/veaiKdXXXAC2eVxqJJrcztCY
ijaaEr4E5h6Nrq/kaoN9QmmTPtrVLQQB1FedDGQvvwmtTsW3/fF4rPWI6zVe2kmp
mllqct0powMO/pojcZDaVVRgXa29JXtGbxcYTKOXZe/ixhJMbGKMlAQrQwEXMboY
NX0syuRD/VsNvFVmP1O5vjXav1gIuIWbZszx3lyloyvlIPmqzqBiVZoEeJG5sU6U
y4WASCFwxJba6uCU7vDPLflxdj9vsjftm+18t6GAk8Cl+oddIE2TQQHlf6KUjzqX
lyQdafNeD/j+lVxioTmEKR3JXaBVRFH4g8WGhL0rLUEC0rW39lAtI1pNw+BZCfXq
4ZWQTHtGX6gXYQUcRuuD7LBSWa1tlg6p01pdK5PBtro94uqqLdt3DBbe2oODnGdr
HKFzvvEVt3sNnyANAkQI3ytUdQCwN2OKQGNs81ELVhFMBtdwzCq9l3nhUC1u0IHv
x2xFrCx3aDnxnsmb1rbZvIBVzKo+XblqayyrqWJWLryJecVp5/WsGgQRrILDF3Sx
4JeNfyt7iyYoZfK8ZcUBDdVAT29RkBbOnwl5U5+n4jpG+jzS/yrXRPAH9ZouY58x
ltr3G5e0U8ehE6SUZ1+exL1ZocKEfZ5AJSTd6bHSYMyf+ermZnnxSqXwBhuOB6xk
1y5QHl5X848lyYFvtO4kJJGJwXt2qUHmv29FkYe/rtI3/qr0AErLhJk3Oy25wbF1
38gEndbcWA9tcu7Pa/f/UcYOUmxEXXFlvoirjG+g/Ue5nPpe7J/fKVgqajV9MfQe
vUSOeT1Clk6WrhF8LBjIaqQwaHTVydoI2itahCAC1WnFyOu94zZ/ijahsl1tRcFn
1xOsmkNZaGnBg5lemQGXUKHqoxnqr7HFYszLf6aN9Hkc9EyqsQszQkzweM9ZBVF+
b5JWXdTgglBpF4bF4zywiHJYmsiCWlsZzmCBkDfKX0ZBrlSJIecAj51dOahd3EUE
tKSafVkzsv20uJSOIQb2z70J0CzZOrG5LQYPmPF9Dg3wn3wPH45cBaF5oW1xxJuq
q4sLV8Nny4pSzb9aUebfAn8gPMnvbqcTsx4I8x81/2+1r2tPXfzLjINupK26P9Si
uv4IUxvefPNus20/Bz4a9msuC4bgAKRmeuodTSeqa4MethvnU5MTYzvgn7/iP4P1
ifzvMTcsgPRkrKVilRLHwZDL0effE81ETdgQAS+qTN7ahN1oFv2kdrgxtvw44bQ3
1jP52O0Vv8k6yLqgKpkL0aN/Gddp/JeroVe6eodeOmTSY9BoqW/gOflvY6r820+0
YMeS3bB+P9+yPxmQn0ej70TQIcUtx6g0x1jP4EtuXnoClSxYjgjb4PJixvM/OPcL
QEelZJ6VeqfROkzGQm9h3it5Wh30q9hwiXO6CXXwbP3v2Umh8h7lgOJS7tRCnEFC
uBMZ7gH3uZHzBwHOaPgiMgR33BykM27NlrbuuLT8OVS8+chdX6BDgldjSKTArsL4
PV7G54Tu8Vvc5vBJTR1iJgZ9Bsp26oMjgy3X8bPfKfKJN3Ppt0Ig4NCgB98Qt4jT
7yxsqGyX9G7oePftO932nKoVbQPDdVZvNb+LWqQTZJxdkcmin6XV2gdy7+KurpG9
TqMDWsZTDUR0m0uutJe7qlgN66gQsNG3eKqR4evpL6gqTbBaDKKssnX7KcCGPQfM
N5iHo/AZC3VCosM4CdfURxTxnPn7mrHPbhWVkexM2PbWJqPD7aNfk4K9pRt5xQ+h
D99aPzaG0gtI/x0F8MrPebtwQOxB89vxoq4mqBAGyJSHAd6xV69YUlyCVHm0Wqdk
Pb58OSvexKp2N+6beOMUYHRf38CwFeVOD3hNXT+XNb5fzrnGeknv/eGXUEFLMJFq
b7egFssHlXI70BAIv5rRLtuz+Y6iuekTZCwy7rqa73J3eWMwqfuj18KtiJa0y8MY
k2jjuzHwbWh5IR5Vvs3CLD+y+tH3G6PY8u/1nd8yHmEy9MCo/hUn0tYT1LQ7VaIB
PsS5c8TKPMx5Qz6FDbrAvsYIm1eXz+eKNslR+c5ZEo/N8XQTkdeVfPu3DK/t2uIy
f2a3e/EqFtaAcNpn3N0LI2moyhCHaRh7O+xK66XR5SZV/fBwRKaz5Bf6/uLIPlBH
rmoElWtgloaOBaUa2ITOGqO/2poPE8T+FT+Jg/mN8azapKDdqDw9mI4Rp6/+QsdW
CgpLtdxG+E0h2ii5VKfsB6RQp5YyS5DlKI62Y0ZbXBRsVjAK/L/6geujBfcyX6cI
OOynlHSn4Ykeyn+ZaShW6vsFQijWPRVdEjkmoR1R+wmji6xr5DCS0d/hy5tuHXlV
r1NzwZ76HwWGZEIFb/sV8FkEJvChLivQnN9GFjzt+B0Xbp0y2DOklOHN7Gu547tu
uPjyQhdygVAUqKZQKVAoHG3MAPjxcmM3BTCCaL9NC6gZ6IwrXT4QmzkI/h+N9PIK
oY9PyD07s9akCutdA2rriiAA3xyfHKAVupnvjf46DgwWkh+iNwEg7C9bKd08cqfg
LFawicowCZ80Bq7pmiDcRs3e/Xf2MOh/UT5KW3xwoFZ/AJvalvhRp1fqCzeTrgkm
mpxVaiWcvS7ALuOfy4YhtJGbtEen3IDt8SQXkFW79QNysF6fm8sCrF/o3O84LtYb
t7Z3FeY5B4xyhbzfkPK6CSVXkGefAi2Bb9DvEz0SG6lQ4MzSs/SGastQsqrqLLcU
2EfVnbqANwf2Sd0YJ54p+pxC0RhdZU8/S9372b65vSf9PGhKadUBM2p5gR10l2KD
VXA2I3PkmpsHc+fl59l7QqMVEV2TTK85eX1Fdh0S18mb0i9a/apt7+nuyxBwV6lP
9Pvvzkawab8uaBIDW+/BCzogOPKCYqkcvZSMa902QP9pU/a2wG+6QFuCnJ7kxSYt
ym8UYWH7WAmBZuThGxuZgHITczK43/wvAdLJMMHDbuBqf7sSmFe5PItfPYeUoyJw
KAXkPVbSdN4ny+RzjIUfIyESZj9RSqaCfib82W5oY3eC6PhJTn5DipcNIzTQ60LF
zdyFilVjkqS5SWN+FrIxqucTA/ABXKwPUvfAddJlJ9z8SsOfvDGn8OwP5pFra1Xx
XPgVuV+weKuO3UWrTEsKBnVsPOdXEUt9HsF3jl+S5HHEEl9IwhW6YSm/7vJDQ/+u
RCVdC/d9/8LjCiw6vX0h2lOMyYyrsBvy5ZxZQe318eNle/4OBdIHhf0UUqnSCpwu
5jDER+CdvvWdDzVBWGefJ7ClIiv1SK59QxYfnG0cYRPEJxyiLjNsxuIc/XEUtGcw
gvmQYJ+l8rLtfAYubYNZwf37zaVh55rwNcsF8OydcVTj2iIffgqMLzkRATrpW5+k
8Ofjcj8h+wNaqJdCVnRoUXWEiSAofAJB6MORabcAReb+NqKmb2x9cZt3Av73dlx9
Gwr/3LfJntNP1OcE7Gn7j42LT4R5/AReMnbK0C+/TYojA+cTOcGIsv5xa9/OcbM7
itAsR9ubGIcMtC9EhJT3/FeYEoJkrqTUB5E5cGtIuLBypgnEwXGu85LGKRzPm5UN
ZUQ9j71CDcFtv9AYeyx5yqcHsyBw3AmLCmH0PqkIslvjTToDvewRLcYZUMEsHq5G
q+A2skhmlPRQLouZFi9srCojOtBurGeS6AEUeZvr1YEcNo1r5dhigczqW7upsqYI
X3pE6BcRpdHcUME4ZAQFrpgGNszLZaPBM7ByC+3+DIcMed446SzA60DFXHt0MSTP
Y/pQ+YiOob8lL89fn2zZjKfBnRJBBnuKoDLGprsoEAWoxFgpseNVxKh0o3c+zMBf
0JrER/wzXgiDkfdEu/8BnAJOgLm3Yn3cLMnRB4kGr6+UarQo1GLqttt3cq6J3sra
XdX1hakpZs7+ZXT5M/IDmOok7mQenkBo35QPkgUKWu+mEDg47Q8gE9OTAkON4jbS
7UT26XZPQVFyJpTN/8AgGbudDFiwL+1SoPqfzbMPGx8cpXZrMXh623PPuYm3HhmJ
asHf6nqXgCZozNb40zWjOr3vcOnnSQupC27ffBeOHDCBHnC+rqQsX1FHjJAfAgt9
T8sDo9cupCBmAzpto5/S+obWN1soi9hCdlMo5rj9dNtcbvFqFqQx+mRE802FYaDr
7HzzKhlbDmXy89bfWZ4E1NnufOn8OsnNp+2PE1S1i7LDiNiLXTZPMSI3Pv3pVclP
d+uwTVCBdd6CspBjTqSbha61W+WaXHgB1SiOwMaipf939YqlGbo2IPsrgBmhcNpJ
HWxXTTumXo83hxP9+k3bwSXMs7fuNt+Qh2xx+ctCzOjZkiFk6F+Y1OMaFAwnFVMK
OvpXbE8fP+fYk09/rubQWK1DMx8RgmZyUvqBCuglANj64yC2/imrrDtdFqymN39R
SUSKkVdaLzscGYD2dIMwCb2vkjfOKMH+CQmH2ks7efDjAH6R2B6D6gwEOGjn5xq7
c4JjEyZqeXVdIGsK61H2OeDTQBHSGhMkkmAeX8RZmKqSax5H8V4FITgTZKd8t5ee
moZ1R1wJA9mkKM2sBACuZHMIbwbtSQbJt4nC3GeV/ENY/+HHoj3SSZo8G9iS+s/y
OY+s4fJtTHuoPdolmZ5fOVMFqy6h1KeE20jP892S/9auJ3e4+YhfR/DL3zf2ZDOS
nGgYCdhZTV5bUDHouW8PFk22XIkgEVXzhWB+H8LAi44Z4VLT9mHNyuLnWJy/ZXxd
L4Bcxf9OdqOBo5Mb7nfLcGiJcwe2Sbwp2gdenkuNEdbVFEi2YABZ02SpIXdu1ipq
mitHdnqHtBJjJwHnvq3tS50MLusIP8pYBBZG7ysRt6Lhf2qytVElidfodEYcWCb6
ITfbRCSJv7IsLYyauO5oWMq0qI+KhrP9jloVfH3YI/CQMQlGBddKZxXEzcW/2SOj
DR2uGq/FAONXpjHI77dZ6Q1pC5q4dH7HhjK5y5d9k3l+jvgJz8Z1Jxql/hxSNEQ9
bVhEIXpMWy22j4KPzm6T3gkRgxFJFiS0S7PZBsR5cmChoi5Y2cPOPIECRXCukynS
bBAHPW3prO+LTW1LtpXOSwTXF7EKsUOr/PT/FJd15iIJhgwKnDpz5X1KLnMNQMTk
QQ+P5glWVEcAqOZy+QfZttfCdWVrQgg/M1s1Z6lGpxwulnWzafhwBfMVSBoC0UUK
FiHSL+LJdBoXXkDQM1H7aczzxsOFyymyHIBbrc1+Y8G3skknpN/zoBGj7EeqxM3N
SNudz9HQWtioOTAV8k3Fkomjyr/lqY9FNTS4K7n/VyDILIjpeaIXtFApI1jmO10G
pNw2xt+ZLnTp5QrhA8izU4VLoszdFSeHTKwzOpqKOabxtNRbgvvonyJIfABldgAT
AIIUGQ/h+hwp7C4czgn1xDWa2ycaUyEh6+KA1x3FRJTDkAhGapgRq0mIo6bDE5TD
qhpVyba2eS8ukGKK3AjObiGMQkCO/cvCy5PFxxylSH1ZTvvMfNrtIVLoXiZRXUoy
LPfEy4G7yOTbYaiWdbLs9qS+IKpfIpBEwN2bc2TKZocofv+R4SgT17s/7+IrFeDC
yyF6Rk5iP/jyWA0oOZlP/8Qj7gTbhkHpjcZxqJS6J32g2pJS6KNga6dEfesF/qk6
OcdZ3RiMzW+YgscBRY56hW847yVcdEdP8uKB5ygWFHaW4YThjrOSk7LjMZ7SrgK7
cYI57d5+nWYoyDI2k4SZi6f4wP3GC+rmRteuN347jnEouYYLzo791UxASU3a637S
soztPkhRI5Y950+yjJhvIO8vgcB2ffwNTndOUuu6bK5Ul71RNwao+z53M8HYduRB
bLWXwfHyYnbX+lpbKkW6/OagxhdvcugFNmXl4Akd0v6C7Jj9GM2AnLAs43acsrdp
seRyLy1HBf2nZed2lvc+VRPq2ntSl5crG+mQrV5cyK1BGbOu4VyXMrzyCHO/StNo
eycaTphLNPZqVoDdpoV4HNi6+cHdplwPdyM3ngSBTVMgHzZiQXHjpLAjw9YyndU2
pthZTYUAupXUp901r0YsQxOam53n8rIX1rpO4WIPGJ1fpgvmqR0WPtCFSoXFCB5V
mNdbSqY1Zk2bSIfTqB7b1J+QL+ZKmbiBFEYg9i/PGw5ID7kJ+tdJ0YUVbqDp5l4w
/G7+a2spuhMB7n3p7qf1fwmvyKs2+Lv9vwcuYYIUi/P0zxSY5+YDhHmx+W/hHiV1
gdk+wTfUm6teaft0oYsB3m8t+T3DR9HdATRzAAh+zJd4XYTyXLFFaaw5DgJqdsFr
nLLQr1JLITjS6XRBrRJHIA4ODMEaiCPyaG3hEwG6dNa36CpD1xWpDsAvrdKv03ep
B0DAiBHmeRj3jvY8hs+rIDliCKOg902otGigpOy4b3ELdZMiGYaUso3h5y+6FvWm
xUj+6LFVJqXH2f6fcnBTtktj7oDt6IIeCvRXMSyjNm6uvwGF7G5hZiJc6LT9CflT
5liM1w3+OZx4DnR93RTdwGWzcd4NlWRn5ZJ8gwW/3GK93C9RQrARyb1UDxBAZVMJ
98JVhMXja5ZQADSSdYk0apzVVGBlz8w5vEYLONzjh4vjcclCXhhh8VDEG/XAsHOS
6nhqkgsBtPrqzRtc6Hvnc1yxYqYaNgZp8OHCEw/8XGKctPmS1oa/RXqfQ0QQPFuC
+Cy51d4TCWy8SgbmmITOhIqgzh7LAzj44E1pm1NAVlT4gOb8sYhRuGXVWK3+S/wF
YUBJj+D1ehMa9OzHh4myEuGQIYL48EdHsbQC3rRYWUo5WsnsFJZRoUxNsE7BntSQ
ibgRlMbvLWoOIva9JpZJsfv3yBSQworTBP3f2cRrH+mZm8z5mhWVfn8YPuD2FpcR
euR507btNU8v/cpuHx8qBksTMzbaCsjs3FzDPxWf6yMUx7FPJOhZtwKRqSwaKEPo
FJaUcoTiclD2Vka1LYoBik0lM2lFbs2WCxkHwkyIVeYjt2E27knwFJPsNjs+Ppl6
YQjGZ61JMhYr0yCjdQ3NvQ3r373aTOAK6iOI1Y5cGfwo8fi+hgQ1MGhfYyV5zKMz
+dmnGu/WKe0rS+sKyShQK8zKgHTuHeugjq4Vab0Zii/l12dSDlNdhRCb7YAttG7r
UWOtDXO7Tw2So9RM/EjFDpGe3JsDn4t2tS5WzfLjxTgh4iWwsHOMl5biPTlcDOXR
bcRf7d5v+WtQRtyFeNrQUCCBgNQG26WdypVop7JdaicfCnvNwMT8f1lYdZGokNLM
epvlFq1IDLkcrZ4fxR81GJ+IzM9T+aV8TqI9DkRPYNIzxcjKBgU6fRwz6jZ1ebbI
UYhdzLVKoT0S6WI08AxzXyY4YBf7irO5kvk/WGGsqCgbLZRHqNcE8hK7JxygjUt9
AyVY2MspkE+xswEnRRt4nwSfY8BQAf7J/1rns+uPJdbDPvPJR0hYq4fe4OFnmkr9
wr+U5Jit4wFXfD/rzS7wtY5y7L7BwqlP0cWasFbW/l868bWRxj5AttZVbwH4rmbe
/QAFqGHxLj7jgLEPIHNx7g6uAqvOyX7AbgIP1CuNAAfgijqKrOhR4BSMZ7Z9b3CL
OfHNFbNuFWlt9ICLBDsqhf9kpNciDb7AF41E5bEMWXvhpJ0IBVzX18lYKgVy01ND
nidViZYOVvZ4+nISegl/GmUnb44iVpuhIcCvlWSNWZg9DRIHv3kq8jC/Upezv7zS
TXg7GSZU0KHWGD2Z9wWkri8+Bu7Kk5efJqtDzDWxjR4GyQ3RyAERYzKBT3+y1dq7
YeS5/tBGgiQy3+hZFuMjSnq88WwxbPSqmauxTnkxLUynQKtaVIsudY7eBLgy561/
q+XpfI3Wl1w08IIyhEGi71nJWFzY5kSi+xiLyaSV+T536mOvfh2hNFUwyztUv0UY
vmiJizJgAQXPlGVr9ihXMWoor0KByO5/nUGZSiu/grpWIwLQutpEQYZigtCxnaba
9nsHCp0IXYzyUfGnavneAGQDNQbgtFKNHedMz2f9pbyflzd9hKudDSX9Y2bn1ZrA
dACH3JxeKsBrqXdKHyWya6TgMLBG8tJwM/BRGox8ELRNMnuvLej2ggXcd6q22b/s
2QJGFRfFCtkqxw7a8hDtj6RH91Mmv4ppaPsIQlOIohpmpihQyqU9VnTQZhf0F65m
nKFACUDfN6wgD1J/nhcI2i7eD5enJ94qijPH6dXnRWMw21DZ7kZ7Mz3p3dzEj00i
+Sb0YBop/C/N2hKfI0abCiWLGLC9sNh9yOFDmSVYpNRwS7rjjYEnAD4FOhWb3e40
p+Owqn0Y97KBldFuHndfmYNn7FwN1MCWjkADQ4Wagp7XBJTRU6U2WxSjYu7xAGtC
bBw3uYpPR3VCKv1xOHnRq77OrfGpekdNQiRjSrWg46t5mKeuyoGpMvGVwQVB4tj7
B3xdKQhzOv8ZxMNoltp+2PG9shPg/7kTLEsWo9TcrrhrLEPMQ6TWsr1dupQ5gBa2
xoPzVdDUHodpU4D58gVVBrvV2RZLJDDGnh8PFBZBBVHp0rPu31Onm/zGjtydrOTo
/SC4b71hPQ6h6plXQsGBo/ULSS/VwadFfDfn4Eg0kGx4Q7bKPZNxIKqY5B+uoqDq
+rn1TUzdV/Pd8G16pnGFJlIF6QNsabGmRk9wJUGi7+JNOK/XhSjZfr4XBl/dgUXt
o/GvAsdF8gqK4ytYh7g9AwjeB0amocWAWqYpSV2jgd+c6ERouPA6cfVzuiAHM2tl
Fy812ZmK2JaVL7shMHAfy5xO1nBTVV3+xXDIn3emKeYD8FO5yCp/XCU2fjccNgP2
YzFSQJKw7z0C9/x0knxDqrbPSTneDjhVTnGdkVTIAc2mfybsoIVLcmRuUmeZRcEJ
fcvCmM0w2XllW7w9QUxjtvyLweM44tqeFM8wG8Q8RoATATRIq5OcnhSWdLuRjFOS
jhFWj0fGx0L7qvw5wTqn9Gs7DPlwJWEUJUcYi0qfVLbF1ODsS86OZ/rwcI2jWNML
V8opLn4IJlVSZEDC3SKWuB800TFSUxh7m9Yy4ShLUgxHF+nmEKB3CuhZlEqzj2/Q
2gg0O3rK/1T3IqrWt4zsjl5pwF6XF79F1L09aNM5xygB/echDDlEm3dLfl1UGAbC
q+TxWHiB2EokF4Y7kudF2Yl7ons7qzOvgHCxgKqunQphi5D8gGAKla2rjLwnBuEz
PiPeReLzQskbiHyCgfqzEnNEYoShJSRVcw4jPdE30uN/HEuQIuN+M5PlVB9pH6tq
REs8e9HQDREGWHaRakpW6W+UohMcR1RmEfZkhJTZewl8jE+jmJcNnTH/aHdr6LVO
ODiaUArRvF7pRLJb0RZaGDauVGfng2upFRzGBxOSMb+8PrKetTwVOBwfLi8qiqrd
L5OpcFRmRzkg4J7gUc5Z9iU0Pn1ZbDbuJoRSyo6xRK/ALSeTUeVbJnIpwFxEFsNG
9gtAUW1LRo70oHeO2L1tahgAa0p5O2tmrIM6NcvnqO1rzKlCm7ooi9+AzavmeiWO
sJoMR2LJCicnGmAlZWwzqDegsVhqyavfMnKCSv1RcUv/YnTcML5d0CrC2KZUaSYl
L+FPH0mtfE/HafvijkSa/QxDcEWtxjsgzWAZJuxM08O1WbIv5K8WMpCf7vSH9rfH
1qv9xvQnAJ8Pv6F+RcL5IJbP2+xy/VZ/Pv1rZQraKYF3b3HbD4YlGJ7n4ne/XreJ
D4iF3xlE8Pz5bTBz4HuUnVb9+m3vRMEg+/giict5MMRxKIBC7tz/7QB5SFTeit6x
rBYwatnmUPs0aqbyETiNoj0hwN+slzQzrqeCrN6iDALH3KG+oqQ5TJ/TasPs0YXT
IOzP4JbkWhzQRSEw61k+YDaXv3vQfOZ2q3fWwFsZA1ybIx6ZusPu+uJnz+SpcUK0
0Cy/fftQXi7AjNZGMc2jtYia7pK9UrOrsjb0O9fV1UfFPsp6l4bSW9yE6RR7gyEL
8uznr6QwZQ/ctwzKw8His0hqoOYzU6jzcae8lNuGRvBsgQ4N0Uofv5NoFTttUtDl
lIel8aYiFyGxKqYlC6zlCBqGEIIvKp0Tz0i1SKa1DQfMfjviANPuyBt2Ztojm1SG
bK+0qTEypLVgVt0KY/rfCfJ11XPcGVpqhm5e3z2FAqrexGIaM89ytMdI349Iubbe
GysHLQOspWX+ydq5To5P/Kcykh+VPxb7HS3g0uXJ3qJNJNQnQSnjn4rqmNdcMrgl
V5qLG6BBXluSuZLw6TMP2BMRXdwb7Jmmio9JeLIju64arnv/CukeEdPovc15139h
+fM0tsTqsPkM+rkyUTXxo+nJXTI6Pa6smn7J5bCV1uu8TzuAnmCLNU+h1f+2jOYC
0h+XS+shGF7vdfpCUvzTpzBb+YMih4X21kq1pOPdQY0WA5O6YKsvaGVH9N4Hpc/w
0VBJ6n/idPu0rN/34g4N+TYcyJXLlV7DfWQ55Fa9VDXSIzoJRqfOFD/Pd6pTIO/8
sNZ52Y79nnm0Q/7jFG5lTVNb4ZmBdUZUX8g+nPwhiLsibAnxO2sTuFQDwv1Efsbw
hFkPXHC/zc4P7tgmvnLukPHQqoZeyDRJpisxm8as/C86/0TgdP1x7+prhKF1iv3y
drruzeElIBihEyk14IsLX0lmJO/RdNwTGT0CkaY45aS0mCqSvJEmlztsZQy6Vwac
In7JPDh3A4IEz9J3F5xN4dZU0T2PzUcpNs1O0y4qr71KdkT1dM82mUu6MLH0OSjX
IfMlexIdv+TyBdomdZJkuNUWS8axe1wiBeMx9J2Y4Vd3IQwjs/9pXuz1DNeZV1/m
mA46r/KGD+mW84gk60TAgjKCtu6nbWwv3uzTRrn9Cku7cDzJgGh2NhjBB7OAVMj4
71ZDpfbDefW+5UGGOoCO0h9nHWETDG4ef2l5dGobJY+yjGa3fuUeUXPDWGCgSw/F
U65+lXL9/PSQD+ZE1f8Zd8uIoY6bNsVJIpqT6Vcc7YB5tCn6Ddtuzm9mR2sdo/02
ii5lpFqt+D0gGxQx5ImNp7UigFOstgy+4txl73n2SsgIk8VjdBqnVkJU73XGzARa
Yu5uM8s+MV+Q9lmPPw/KMUu0EZq22wNtPvIiT8njXMT9vXK96E8rnBcVwaf+u7mO
pl9yymZLQDFoMT1bHojdwMhv7COcaWc1fqaSZP5JiOHUUUHYWdnv2bxeKUpLVsXC
1Lk7k8RHmaREqpvVSIJQMfhZ5dNKyZSlmBcmrw+dZMfTQNn64Igu5nnA951lavLe
bPeFihzPAyWqY51dK0vMJmPoaZ5Ylin+/2aCgsUO36RCVaGFr/+XCyGKUTQROIii
S2oR1xI1qDdFy1H0AOlRYtyvlWNdLMUt9mlu0lkfaUMtq7Kp285+iRwNOibOC8Et
qxfG+/cK4P55xfx65nuT7Ft0h40zxIunm6zhyRO26LnwVxRY0QR8yZ8zgCvLoMxU
MWDLUE8+FhI/tzCBXKaK+si4Y6KdEPqv1JE4k6INrn6SEACQv8j8rwCpqq2Sa6IL
aTqS8lvw+qK/8sc/TSMulKZxZ2mEorIzBfPI7JRHi+pbwQX/9yVFai/7m7fWEeuZ
zweMeN5dankYuU2Uj2JPfWwx2kU+ZPzGvPxSVQY7epmxVVFVVWrMnoMi9O/5AIID
qttkwYLoos4wrqpCMrL/oNnshy17XTZl3Por3dZ+9Z953BRXFdMjMlLxgmHGSlvO
6ABDL2XqwgzlGi0r0l4wazOETF2OTQLzHoLExyQIN3CvOrjw32lFUnPaUHZEXuuv
GIOwzRNqfdFOgDnrNctXb6GDHWqRVZYA3iRdM1X7j0mu2rqiDf3/yC3fK8a6Dtxz
KOoVSrNP/DFLFQgVnBnggMlKFExcTrbqO9YiV98w8nChprX6quVvQRQGKwCnlnEU
M0oi7MngGfKOQLO67c0a1qALSpUM0EBi3M0V7EECZ5KM+MYRPjseIuUxD7wu3AYH
MyiaqoMe2EEPYHuk+UjkaU9KYkeYzO1mLgUzUGAjl3dO3GqtXChxJizNGl31sM9H
Y+gwm6LQdhyg5M/PHI0e8ZrkPTWO7JOnUzrWoitz6dxgRWmbt5X7KY07IX1E/tx5
zTAhL9n8zgu6jo5cZvlk3m1YwkC19IxjIDVD74ucAW44VO4+dqc74Nbe+alMgDHA
f7S6aC0hi5mwPTSDLxqicsJK0lSGFovb5fF8Zjx9zSSNYsRiLNSSoQC8gSEWCgCi
OAvodHKrIfkb1UCy7794ZTqK5nXLvkfoEjY5rLXWvupK//y0MkuzRZ+WqFLbsF03
2JPPUG1Zykuf7MQpTRsDUa0tTYa3InlYcKN6LbEttupwb9dQBeF27OF35AHPrrfs
p4be2K1FuE36ANNYY4lwE7h/w632EjiSEkJxBybA+Zo6DREwTZRmLB8QtqcREGj6
9UQnX+K0jOavOVlZxrgcSpLvNz9g4l/9eB7aZk6xtSEhanY8A/5Mku5NsYYprlgL
0y5XLW61L201uPSxxkdcaYmFn8VshOIXH4mnszhfmOPj1x1+H+t2EMhGaCGKtaQR
wVfXunB0aWVgpY1U2joKuK9R77rVtJZdde28KJ9VCs5pdlKLLsmDDF4DCkjJHtVf
0Vxp661rhktz9p+SzY5pn4G+564DrWsjb4kO++5V4gtF1qoOkJQ4agQfqHpsn8tb
KVXxcUhxYucpA1otC9tqFesd5g/F8/oR1KKEpQyQ4sT/CmHg0hX16HyE9IaOTset
HV0e5zP+XaPCtad/iXWctjSxudFmPvRIsDO/ZnpcqzsrU/vhSrkTzJcxz7R+m0Lf
mMLThf/CI3SwzR6icwi8HZiG25yKKMYEqDtRLhnEiuQgFEheL2zpp5Oe90X2BCCi
+08fyHWQIN+MgaNDF6LrJ+6hPcCB+Ynhu8g/9L2d9Zd0k6cy5PzuS3buUW0Lkfk5
35pBAVwixHWO27pLIysNZhEZzevjrvR19m0L1+6WBC397IbywQRmFvsDT3EbTnQJ
AMaTYh1OdiZInVXxVgpgZG0Vf1t6P3c5l29MSBKKxm63aEuzwk79XtN0ge+C00eF
YUyFvLAWyc0hHr/tjas93/dm/QOIjD3iAWXnc13BPPQ/X6EHYR0DFL3Ow4RYm/Tk
7Fja8R386i5v/KYL38Mwye06aRN/ugYq1iVdOjmd8yuVEJURAmkiwIO6SOtdhdwj
e6R+EEthmKZFTczX20KFflDz1PPU0W9D5Z0JR4ynC5/vFLOCvPivSZc71/jEO/mk
GeDAxW0TfAZf54raxC3ncmYMtpwQONhQRJvEx6hpgIche1zR0vLaYszNSYu1byeZ
XU6GT2G4TREHKkfT7IfEp9Jq+ItjdcHRvWVJcrRd+yyq8TUOsOHs0MhoPqpWytGU
yITniTnS47xWLzwstXjQT233FpHDTJWjmtQy2Pwgam30i1uJ+uGgX4vOfTksBOZk
oSud/3GtOkoUGlwRoULXsaCUhu/618YgLo0YWEpR1tksmalqyGtjmLPQyUS6DHc2
BkYuqQBtjc6UBLBNLNMwXp3s7SjsdkXkjLRI07RznkNCA169FJtx6AD8k/0sv8Hx
EiTTGhWNrYl5tmO0lz4zWbFiZdiv+BxF1MJKng5lFzo0Q+SHOCbVKEFbDr/FPR/f
uwBLsS7UBFzEVEZD9QM69MZYiYzl6Vxu1mWbuOsj2Fng8cYKQQx3r1EtWGjAeyJs
wA8LDbrkTfdOqxt565jiEE4dpjBFsDYJqT+OWBgRh1ThsQ1eUulmQ+9Cmi57Gduv
M3l8yuWsLuD7E2nr7BrwCQMTa0ibIKK5I9yoDiv2/mbDP0y8nbXi7zmWGKI2EJvW
HwvXgdiLDHDWT0CGv2QAgS/FJ9ka7CV4NAOfmhUT7a03bdmoSQPVceodbtuaaSdJ
h2xnAKp+92x9Xdgem99HeggwFFCnx3RtPsUL7EcZo9krGz6byAB3TO3VOVxUiRbD
earth6AaPtH7RRwyfnI/Yf8dAI34v1uPLs4W4q7fHmDcyKcLzuGg5pc83W5Qti53
wj+omB8+j0x8P8d4BCb/pKhXzu0ksjBcnaY6aKk+aEcs+WgxuChyBICekccs6Y1n
1NS1rXJcr/NEAm2dyWL81CPtjflHzpcUGx2zHoyAHD8+1aVOUD6koA3pAZV5YMR3
pb/6qh+uPy45Hfj2E+ED2BgGjSTwKegN44iWf++ClpznBPpGLpOa5yhrnp5iNyFY
SA18XdCvrZApXukhl3W1NqcfgOqKo4+ioYQtWTgPivPBwxn2aOpMEaSHc8tG01UP
WBoqS9edoC6mM1t52lDFXcqv7HwqMPKqKOq6DK0HiiUYu1RG43JwX3fvHTG5t4a/
j2IfmmZznS8+apmEKbHzKE3p+QyBdNaADSaiEdCrSKD7OOn4b2pukxtOL21g5YQi
KAEYg0l5ytpWqDd3X27XxtZFfafvgAYoLkq9sfxJkBs2IS8Ijy3OBZwMyLrqxbTQ
cOp7U9MZC3a+I/xBBJZfzxj7sPOOIaQ71kwBuHeaP6sP1BQyUrmDKJlEdwBtTVwp
MO1+RJI6MJbzeNEqthYwZpHGRwWbjmMc+F6J6MhqClt+V7rmeCnr7qkONJURVdUa
aUiCI2Pl4XXPwirbQ7NdYAn2uy63fnXuv+WjMd3vl3xvEVYu83hE6D9BqWbxBpg2
zKxYPnahIdgigh0DF27AOIK7gIqgseGTF0lXS9AwD8b8x/bRGL/Yr0Jc0Y0UxiFW
7IljshI04EKI3xLWr30gRsaj2rpGrOQk2nO4VDzvMQy7/YoAa/aAUbZpT4jkHOuF
rv31L0UBoj3o8WPWLnt3OegbdfP+DW57uysBokkceHv3FpAClYkMkosBgpBj7I03
sUpZC4N/KIe26aJJyG7dJwdNcnYal3EHaPg8E87SdZPno3DvlR2STMuvrhew2GO+
/NdT0D9m8C34JqEXo0UUSFPfwFqwELW1mWYVYzIXRAB4JNMj3r/Tbl5zM5zraPy9
3SWsLRJ7jBrIlwJmdmkeIy1N6hczZG+Xhxff4oiSmp0C2ivfJUXlvzp3xmotxxEd
ZqBKTlMEPnSxyjRfXpnnZpwFGto0HUH2Wq/G2Jq1D8/aZYGQingsTlaQxeMEgHAx
RB3QDTtC85rkXOFZUrzvVTfcewNpc1RQO0B8mLSjaRFAebUfK0ZLmUoOsl7A/NTd
/JjsVGXWDtaSYSh/ffeMOAD8YihLzfuP5ZLoAW0hpbBGkEFhhTdqxW59P5Kghe/H
lya/wnfG/KCw6QfsBnWVRzCsAQeC6lZ3GSkl/mDVd7A3pIB/qm0wSR5FekhgItAo
iaVZ0VrohpacThSc5Za36BXS30PTZPwrgPD/Gd2zkHSg0gc3yrRmr1Et+sb8ogE+
NyzBKX+GWe32X7/gRsazc4m+LfC5M/UdLxTv2dIBgbuhPOjDjOLIjMljQhymAIXc
XlG9DT1rKubk93sQDuziJNUBNl8ducLsvP5avjR8jJf00niNyacVQSdVJ3mQGWDs
CZCLuf8y3fxni2yCJQmZt1iBsFI2xh+UVtHiPFfqtzRrC41uoP/tEQDxXGRRV9y2
yXmab/bwFzXcqAnA4eLg7UGRjdMXwBrYqgHkA0EXcHXll/XoJleMjk++638p7/S4
1OS9//cQxV2d80dkS1ykwIGzdBYgDHe/Rd4gPmEPsKe3LWtRF4YK7QaGlWLwmnRX
CjCnmzjN0YNqDy6Hn3MrITFbmsq0ztPfpVAsex4ZXY00AkXEM4fnIA5F51t3Trd/
ocZiH8Y8NbEm67rkHy/R2hndX0ggOk/9pHH+BsoyBsErzcMUv/Z6N9gtQPCpVFe7
spUvKinZJbMvR3iFD9cH/8uONdkQq8sbeemSm2IdLXAH/oaZHVoqGlZ5bTTiWKge
QWR0Gt/jGhn69/SegbM2HW/b70YycpJXh589UtjPUOiA+e9UlkY7iNuCiP1KXRuT
vZFVcxEMw/oMmMtLdTnIT2mIo9eVAYvFRboWxC4KxOd1brFgMkmKpzu1yZPrLKjC
4jY3d6qT462q93Um3wMqgQ1CjOpE+ijJ3Yw+1Jy91+P0FNaOoqKb3AwhnGCIbEtq
FX3HeOgHVvbHeMl4eUUjnGazP5FPX+gcLsGmLhNb+WndfdHe+Do9dZUpgA7jTi/N
gt2HhyIEeAbFfL4R01EAdR4GiF5xMlZkBF3x4X91d8KSOjnhHDK2AG4RQp0gUAL5
XbP9MJ0yP5s6KOEKiuoFyfQVicBAQeGKZqA5Ux4dzyjdtQkeWxd+fTrJOVtjShte
DB5uZ1YoImsmsbvRoecz/lDO5lSUUl48UkbeRLiNBeBzZW4w76W8UE/mJSSePYcz
CexMbPl2nSpRZ2mbY5plVSuGhu0CS41ob/CCHAmH3tdotDPTJ43gi5mOjZI4fwft
3yPXvo3N3jvxmpb+c8GtmQy6gAbygF2m8JgmWoM5p9hXYd4xEKmaNITY5bfDXkQj
l671ukdxS8dRcNmSqL7JY7aPct4aK7xJhGAbXlgl9DWYtfT8gyRZnt+gfdCRHBqD
d4YmSm6MmKk498Xk9Mr55fq76RHf69VN+WCM1qesbZaEWbuPiXArPfRyXGzG8xNY
SyWxJG+TPxAgC0EXJfFJpTMl7dQfxSEUJ2+7rHxJifP7anXi5EyZOYbdvBMS12SB
HrbzuzBgoSmY7YDZpkNiznWoe4j8Ykxajk56nr2P6uw9vdY5smZaf0Up+AtPRv9L
ZR0HitHO+QvLfmBgg/ml7dDVJaNIF79yNwoFoavWreO18+W7oHTY+zlyq9WOC2j1
ubk26vWK8trm/+MYuztHo1yCeoS14OPGmE3OJHlccdVqGCFm1aLqFU36W9TwKKOz
c834tpLh1ZTcJDGGWqpAPKWrEKm8DwXAVfyFhoDByKkR+SucjwKvu05lhchapnJD
BbM75ooObt8cu/oAtEnQni5WK4luyC8Gu5M+tm1HrqzoF2t5moJe7IQnx2ih1xf+
28f8pAzClGsjam2+tmW8Y8lo+bWAMrMDJTR8aAD5infRIQCx8aswkl+r6l18v55y
pHWOllwShS/pCGnJ7Aq0+HbB/T6XcsZAFwuUxHcWnGqpI3nrKIRj8UWIrJUb0d1Z
/t3F0oYZLtMemB7xUu7XOHX0t2MSCnf64WGXQVcSpjwsAPT5qzI847FyTH57t19V
2konNy7pskqcVLWc6ge7hkHwYoXBd5Wq/fWxBYl00/bTaNJ3CyvUlDRdDHQFmb+N
jX19ZhXhe0v8CNWCpsjemeA/RciZDsVg47YO33nP7dHu/NmwHCWHiuhsraMg69hT
3aP1XUojxrmZD6SNxeAbsoysCkzXzuk4n5TWk8ck1yi0itIeUwd1crGjJiuMqIUN
A5t9ssjBBRxBl13MhjcSmglxkmkoorzGfWV7E9VJkoNDnhqmd01IFJ/+DYOQ4cOT
5AOmo0iDGjQ4S3SyIgz1kZYlB3PWhny9wFr3zi3lpRk04lnYF6NlrUZtNO01whqd
4C4r0ji4N261zjHndXa49bAMyvQKgmsS99sAeJyfK25OnRUAkkhP8go2o/Svg4l9
E5NgRZXrx/agEH2LfAqs3J/jILQ5tKcgKJANv6tByu5YuvD/semkDZ2nW2OLm+Iw
SIYu6ImYJDFoJ/rZWmLpR7SFEPBcKTRonDk6h35uWLrSSJbVS5LdblwYtuJsreyW
ry46sd2TP/jh0BEKZORupGrZLe7DbQ+a63Wcsbbfxw9/Wvrdng86ROMTbSXfP5Dm
nkzBWQaDj93JGqPbcv9ThBH6ZM6n7lXIf2ZZ/cAN+4WFt7HHNKBjsUM/583jdR7D
g7ilV4f8iMzvrXXo6I7L7CJWf9Gmdca4HpR9NzSXx53Rn5/Yu7LoHv1V4Vj4QKfJ
+kjMkT9WZD4ONZP0R/XbzQPNgSgO3urfFoe0B0z86duwwHh7+O1yE4Q0Ta2mYvoA
SO7ItNCMV+ulgEyF7n4jqsD6l37TtZhn/QXS7q7hS259noEuDXK3JT4tYlMsivSh
QFSpv4M/BJfkGFcwSFjHJvATrwN2hTk4pW4q07ndytaixpRaopTc3KqrzLwe7f9e
8GxsC2NZzPkl1ScOBUZwTU/J8AsQFjMLywuMaioaA7a5jeIwYLEru8QlhAUIOIOF
d9b8JXSRfX3Tt8AoNduRtGYR7jq7QRlSsEiv62DMzy1R6okykaAnwlfgw2l1qVAx
MRVDyrzKs/LWtw0Aw/T4egjbv1yDNBX6j96ciyZKtnKdzBehUnzrW/FSwZiqCBPO
RjPgLzYf7mu7A8ZdyaTqMPpIwSDKRx3w21HvQvjgi5UjEbjojtSqxkpWPR00ki7U
LKPAYh69ddee8jP1aWPeqDrsyFrkzgUSRmTZbM4kSzWKtS8LnMYcNaRqmw/JwmbU
bP2upPXpOzpaYoNmBhGobeCl0VKDlwy4RI343PejyVBlnS9RqnHmTZpI4pKf0L62
RG7e25YWndPW5OcJDqIuCVesuG8561yyZSnHHxxf32pkJLVLpJT7kV2OgtPnu14H
Cb8DApPxiRMHajGjGxyJGmK0ZRqHAuF4ysG8E0mAJyQLn8NDXJ18s8uaTi9+fMVJ
I7AEDg26NdPYpYaFiGVujfJ5r8pmbdKFiTuW4W8yFRa1lg9eXLC8G3rRg+UHv9n0
2e+lbWjs/7hWOS2JgvAISk2xD1EuDO1s/6Jvg/bzUYNP7etTM4KPzt0rydNy5sCb
QErUZn090Cg1tEbdzrh2dkKN1TdTVIgcxC++QDOAthNMDwlQYTc61iaf8dfL6e9b
gQwCx30+22nch0oQEUntcVwydnVkqzTWENMzSIGvT+M9LtKpRtdnp7tgw82uf7Zb
NYLhsu2AvypuCNRz1lKfE0toLxS1QS2iV8Of163WIjnZorZphuRoKvU/JCZteIA4
RbBu+kUprTox0yg38aP8awONRpjDX2dlTgf9cxN7JsNlfyeMKr90CuvT+90SJA5c
XTnnrSU5GOr4Uq5dR17YR5icBLgRkdUsvAazDNIdRGKVZU3HVpbevSP1A2sqIt1O
W+3B5BVhhPV5+1VOFGWNCaTywNpot8uADy6j8t2BnwQ79xAIFXsu8B8ofa4oBF0I
pjHJ6F6+zFdaBaxe4hnI4ICTtdmnh/UbytyN8PmwehhHh751frrtfZ5TFNa/EKgG
sN1MmB1hZnGi/1HTEd0zNb7MiaCNBi87oYCPf8BfIKG+rzDgezEZf6MXhERFeIxY
+0zX5JFDjog62kuFGZvSvK2vBqt++Rs62bgSRzCrGc84EvyZi5od6ImI0W5khUup
pmfkacv28KVaZnk/xPasIttwRQim7tUdPUFU9FOlbZ0GP3ztZXX5uW2ubzEbhmGf
es6bBa6Io/LjhvfabVRPCaU8F1pZsSkDXwZlZYdTb+/uYqx/mC9oEnRAkn1o05zS
pc1E0YDXAom6RHjKz1J/iE7Jsz3SJHeT/O6j0kl6S36XFSVb4y0/7KT8O9ARh6Fj
x/Az865rLVGZejIMq96Gscw0IcQWpscieSh85+cqCsU8BAGNR5ELnVJAqSZ6W0Kj
pzvqpxkdmz+1kwCDzTGVkkAuB4d8ZZzOKFa2Ead02gRIqCgo3Kks90sK6cQOt0EJ
67FBqntOAZqhGxml0E4K4iWEnUajCQ64weTpdi/YziHSl69DZ+LwdxaQ6JOD9ywm
+GWdjDA9yS6SB2Va0KPCTvZA4gTNg/0z4ctcLrwygLWaReO/RJXgBbuTUZ7WYNDG
IcskTrFs70T0ZgCmMHuq4avdX9j1oERdtsD3SrYzuuf6B40LlyrC9HtfJWf/JpOn
2e2NpkrPDkRC5vNlqK6kEt+I379KPfxZfRwS6yOBFMv9ANTT3LgqQ5pSwAkiJNKu
Ld6D7+88r2fU3XmpHYVUaBwMzL7HbdC2b80/IO7mBJp3EGkYU8FhiSpRC3fWEk22
VGxI4FySG36F7VrRK0fb93E+ZKh18/Mr7zQ41TwNw5aBc3hFqSC6eHPEFWIpBVil
4tq0u8U7S4eNDeBHQNe2BLowEppdBwgVT8fhWMqEyaRBbp+TsMPxooqTPfHpFaSD
4vFHro1Spb6D5hCKMGBuENvYnQnLTvwzKfm4SpwX5Jzpe59yy/2U457a5CBZrZh/
gli84tknMGZ7BdrbB8E0mudriH8JYtMa/htSZqHx9Onjh97G/nWKzfzbMSeiFsKy
fuSO7tULqaO59l+5IZ4QEvvI3b3/y7VL1C4g1+s26j6b0T62fD4t8A/2QK3H5eIK
yH0OCI1f4YtbL44atdAsSQzVWai+EcCrT9a0D5ZVbrv/Pi69wCys3UTugTS8Kino
6jeKWwKB3G6reEOha2I+6wwK7vxean4uZnudWFDWfnX75p40DnvOfGN9KEgfYhXc
hcA9osGFJMlF93SFqfWE2E+XD40BEYZaYoDWV0jsxWAVmaU22yPKGK0ui7lQQQm2
KQUKv26owaxZHPX7RQY3Ru0cNmLksxRpot1kF9eZkKXDBXAeG/0ty/01V/SonQoo
0UY7hVTTpVloAnvx7H2lQx/1FL9cClKVdwThAUdHSV0GA3eY+WCgCYR5T8Hwfwgx
brwJg78ISPsEv/ufgGAxIE872yJBRCV9GPHW2WoxQkuqm/liVkKsDVTEVsR4dDY8
0/DuJHucBKAqXTwmy5vehZDXqXkuWPLut2nUTE8V7McpjXzVtOrFRzjuszF3AfWe
YLssi5wSdL29osdGr6yEU/+Bn4m7MwdxnyyvI1gt9rIFSjPhpgvLpvBf152IXYO2
0HHdv5b6n4Evf8voQ1LLKIKLp+S02f2mimtuZlpy9uUjhj/Fp8syUCb8iJXGlkss
D7L/aQ29zAqEVTov5N0RjxU+CTk70Y4XilsYsaSwWlT2z67k+r4Lp3L2qqnw8oWi
cktr2b5/H3xuzSh+0i7uRyMy2A15M2XlQTjNe1w8V69nBqYSlLEfZcHW6xBdzYAI
TqRlm8iW4ZkuTtKWAsehqJGVBD2fZv5Gh+NeMLHbwjKs87i8MVemaPjjqwzJkAVB
EOT6BKeo2eY8G6MeObnY6dRkiH3AqR5vSFe1JycENaJF2StlRMYai6YxQRfgvolu
cO1O7KwahYMUigI8AARkVmjwCn3YRhW+XOSwnrzA//3LrZRLFNDwr1QgjKqjCODg
bYgUb6gryQ4k2XwLfo0rlTgoAT2DPSuiMVZ6nQ/fB10nRPc5D0+wFE45R1DSYhL5
00+j8hEhMmxPl0fcd5WfPHC61BAJcq1mcNqJekJTEXUSAFH0Z1l82uvTSYIDacqF
bFzNuFcNFWXKqFgxeA06H2ZU59izO7mk7gmdji/7xeZftiU9kl7WK8cZoQpJACtM
X6lX4BMm+xAjJ6X04aGcUMNkH7uCIDy+2RN3h2dPrJ7rgp5ZRcjom8e3AJYkWj0O
PlMnXPbGO3YksLnptfunD8o73fU9R7oAA4J213iaSfYhLlkV/+oZeGn44sDt7sD8
ijL5o8HQYjLtGMuWQTpaKKD68iqd16c6X7LdbLGxOjPuD8TDI2Q5P+Aa55X6rWzQ
1fIbErvrzenC2qHiywTZGiyUIQvV6434BOuqIK4nqSSVlLBsbMLQd0sas88JcLsW
9cJWAQyOzuxDfkSGFXcFmN3er1wQ/z94MTHlowira9036rRfpXGBoHkR0jPbQ88O
JsM/psNb/q+8G5VlUfVOxy5vUbx/rptwlhto1eGF3jaN1PgKNvY3L07xn+thl9xI
S68a+xkWrJt0E7/5piqJtychGvVGYAPyItlVHa2LFBvhZcEYf4bZ9sivhIU9Bevh
bgmvkFzFWeQWqo04IFeKVWyPnasjl0KVWrDm03ugHSpg0Te5SLec40hjiQeOuvKK
Yil+2h7334ZtSxupn3rwk5hL31O7PwnC7DPTzVDufzQ+79BnhkBWV2O5IfokGbtJ
2H5IBooRB0Q0jAi1z83FNRVmoUYLXAglUTWKI910se91AQbzvMoFzZc8rIbGLfrz
RntS1uCAZHjQQZdPnn3j8QGgFBIRh4pk2mHuzqcIvmbKRoIQ5WbU/lPm4rrxuVxq
j+eXzD30tqKSHPeoUM87c6XUF50kfT+eGl5eh0ACxTxu+7yGld9IFmPUAkAd3tFA
sr4rfuGzT5MJxsJLjKKP2fTctEKZOXLhEAe/J3jkYKTS1csQE6SulIp46xJaU+HC
ik5TZkLGJBJvXl47fjHoPiwFPkz9GTQ/EPj8OU5kkrEgj5eeBcpBmg8PtxPMW28P
H7viBbGLEUcURKeKItvaahdxw67ndmCdlVPhnneaI6PM+blb3ZaaNODVAWZWdM8k
ZuW3Ht6vLf67FApEitnFKJVm0O30IzORjW67Abx4KYYU5fpcoyygnHsgZZVXS8aI
DA9s1e0ce8tjZVQ7VXNZ37VaF00Kt/u2FYPj2lqzFtMgrCck/jKredLPhB8LIEiy
v6mbp44YRY2R+MWeHh1/0ClGLFn7j7EUVfZstTM4xnCIg3BcjwGUeBvSxn7YWSiy
yPJYZnvR2zZ05TVFiRrVb5ides2K96ugjbgQ02gAW5AcKp2n9pitnKaiPzKLaQqj
biAk74BWdZLA5uKZw044PHY7lr9G5+UhH08wwLyBmDY/NmD5hNNJCKnKnrb6TNM6
9b/bnUB5xTzXWsysso3ZvJPh1V24L/D6r4WrFhi53jheUghzd2ZqX5k33VFvsKkP
GrpQgmI8PfZ86Nw9YYiapztCYrHQiDGbtcQUFljv1/szNRhFfrqtkXbBs2z3xZWJ
66Wf8BeeUHn+17AB12CddXJqgpF1Kx2YVuzMFAqDW0M05T9OWMoPwIgrQJcHV+Rz
v4boeld47dnUkoEHeLTSZuo8IGFfeMsVZXkoaYrnEKbd/cZvqH75xfvlXBIYvtf6
jQMT0AxMLK9f/s6Etk/kMFhOTpCijH7wwBMNXH2vyKuUoLicjqT9zzlLpWbZS83D
ilWdZ3JOV8tVKQJyQCsuSKDFJyFeAIYzS+/fHItVJ16P0YoAYL1RjkQqZgclxkV1
nO5E6H+F28WKo4mlKATS5tUZWE/v52kbJZZ4Rdxmbd7d9EwgefgVf/VZOYovAa60
L/u367EtCb6iO/1xs/PPiOLTsSIlsallc3x99ynq+vUjXz+O90qv1fYt7P4+//RT
2DX4pjtyCH2knc5Z78OmiarqdjroJ+9zbDqwaUxG1ePDTX/uv+uR/ahAHqi1LjFy
ZITNQanlWCsysGrIFtFWXPgtp2TJfP1KIngh2bQsQedPxt7YXCXCrUSNQSN25npN
QTKYdrv4SGqiHeiYQ31uxiZj0Y93eKm1KK/0JStq5y133zDOmjhU4EYRvCjvMS/K
cSDYsyx8yJ+SEG8zLJwz3URo+/5mSfBb4bLTq2arag7wF5hVIq4kV3BpZjOr4t55
fad2omOr73QjQW7ySRwSNWLz9sksvs/kW3f7ooaO7chzb/MAPF2Vjfj/FhFJvs3Q
Zo5BAZ7O1FnAoJvAQSzPlVAX0P68zdtbya099EsICrZScn5i10ekq1OvWrUjDOZB
pEAnE10qW78L72Ui0DpydRQqQUOwz2slGAMcVGUjjsWgT6XP+sViDxCNuvoSyxsF
ILo3lvODccn6pFakOgghTEYy66vVcMwL/bHQPE9PNGWc0FGRSLm4DzGb0L2Un31E
wEWl+lpmTVFgnfhS+xPbTXpzS3YMA0aqQxRIhFchrs3xnZc5F5Eq/tvfEHnPKTEm
dh4bF6qvnAawVOssuFZp3yUD6/jOPku9poVyRH65F5vt9J9nUBEnyalw9i3Xvbk5
ALI+5F82/TIiDUmsfWiCmC2RM7cXvkV1ltGQGDhI3aDQ+BEJc1dzsquyWsK6wfzE
ib9Z7nEVta3RH3VPG7fnMeUMG77zngw4K9wIxCfk+pIVZPzpGrtXuJVvly48bmgn
4w5YF8BWCXF+i7iFqNVSAKIrX8a5UStT6fSY/j8mPm45WSCxMcYwWDPIc7tGJAd0
Q9mus7MzCnXU+KCGSjoJpMo8qlf/8jOSBDDyeWDf0T6cNvfUEJavjGvkKubw/xgf
IIGGcmNFdJuhT2Stm16LcniLv0VLyVqZFatsx4oxm23SNdeOFGOFqX1EXBVDmlt7
ZAXSVv4TU2eoEFVCfw976zeBCEd+UaCUdZ7x7POGYzmt1Wc2H9DEpxwddyvJIrtP
ZmVU5tC9EBVEIgaEvpsOSZoXzFxml6H31lC/UWP1VCy/uNJrUb8Od8Fa/9nYCnNB
BEL705F2aZYrZr1TKpzuBEd1eCc8zcd+LBPmNr6SsPA667Vv2c6RDk5vNpM5QlVF
fypkwRF8nKJHeWMRdLzf4Ht2GItQxzCx2dKCV4/4Vqwf0xQfsWugVVJ7n/1+7lzV
KEcPKOZjX2ixh18itfe5dEEQJUnJ1haMTDNC914vzAjw//X9Kr1KHup0OE8SsNJy
MFAZGcBv8rbhI8QZlK8ymxp02dFI0XPkuk3UIfkXg7OLsLc4CwKRKCogVO7tMmlH
QSZqNBFUWE679FFLI0/tapkKkDNhIsGXyWZ70oySfhSq4j3J7EMHDiGl6zoaFi5E
SrgCH1R09leGGXSH70WW8CiHXNsngm17WPb0Jvo2G1Zno7X9tXFZpahOUDkIZVpg
4zBfYRDevyjS2QFbTHw9SPVTyMI346YJStSHUtZL1NRusOe7n5jXi1iwznmZHVoG
iWA1sBfEL1r/MuU7MinEiPqiPOIkkmoOlJeU1p9cOeoA2hwJOdTLOIUrwUYkUsnW
6snYDU6oZ26QNvXJ31ZycxiKpUNtH+cMKweufHOUhDpon+9sE2kxXEMkVz4HOWFz
bfe2c6c/SBcsxVxtIOHaaeLLgXR1Bt09ObFI3JkvW9SdQu6AoWbkK+s5dfAdTFHo
7Mt1XpsBibvzCKgM4xyEBe5z1BozcZKAG9kY/kaq1FyEpMvC5/xqJZLwAL+zFFel
52brfqP0BS6cNUZuy4NlphJf8DefYWjSA1JuLAHhqZjphMFPJAvXktaGhnqmDbTN
I9QOb1plcsF/z0QzEcj0kBdOmyHJvsxqis1njKPD3ulRrIXcvtPGh4H/V1hMetJl
J/wVrshPtUYG26ICXW02ZeQsPqRFEpKtDGjxmnR5aooyCYDJZEAPcgXcK7G8PGBn
ByvcTxVhMbBTMSuQzunP5fJTwAQ+NLlbS/s5M4Kb063lRj02nAY/x3PmL4nF9EBu
VeyKXdTK/N/O0iPuLKLmRv1eYEu94EZsNXU/oxMDM+HF3nRiFeEOx4eUe5KHmDGg
pHQFo7q8zPSYgmbjlTJcIDm39969le2xt93MBXUzqZ8bGPp4YaP+KTDVQdml9+Xv
a+VWbhocigl2hAUG1pExW8fiexW5Rj6kW39/JJDzdDWEvYdwk1mE1me3BkANKxnC
9dhwr/uJnD2mYmbohLaELCSK0vR9tyckjyM16culxdLB4Qpb+F6sW/2zVawtkFbo
ID26dbRrnsDZ9srgxy0++4g+Xq3bkO8WNYzC2E17Nz2LxK7dg5ksaGN5qdk3zMiZ
3e9LLqa52ylFVDGnzJl6cnXfAeAZ/nMtCNamAzEjZ0uEbaAvLkQwj1Wt7O0Ho9pj
wNu52r/csL8UxQRNzRGsl/OjLyemgS8MJnitZOThJHlf4rf0G1igwhCPCjiMqtrT
QcC+sf3rAUvtBtrPQyzz0PA+iQpL7wDyVnIU1r/PsjUcSbL36jS3rv90KSDew9up
oq/Z3suBbri/u5rKuPz+F4nKlCjNNr+kFPUntDXuv/wYz5CWJUopHrRJiUUxrMwc
4lciW1M0AwjdpOdabAashDzlh9rMVQvl5vRwuPbWWdVgr5zMffELeIQT30g0GAxK
be/YC/DdAOo4jZtu4GAcG7+MQioJsGR96hyykkziEfgrUAnhf372uiQNL6raoYte
BBaAASNz1wk/PAzY12RA2m94ZwJnw0kZq+Em7EpRZllvtI5gf7DMmF0UE3EsWyey
YSh8VvRxtaXFT4stGWGYce52FnJ9W9OIOzpHmI92hDm2h+xseSN6LsTAwI0/VQO0
v7OQIraHajco4V9TMHANiio3YoA+onrhv6QpIG8D15aBVA/6p0vM/2As1eyDtazm
Choux7ioILCTKqiSkcwOTGg0Zd+Z7uI2BSX0WWCore1g7X1PY/2uPflLPHvWzy9z
cLIKfXSZZqQaAHuCvVLjyx9/wP1NO3rC2D9QeOaYIwBqt6y4D3TQV7b7n3hJGhR2
KFzAWxdTFicVcpXPWJ1SFUbsdZogDqYzC0iAMJ6xlrQgtBKzdw+nDVQiDg0AEoiL
az8yExEnoAzHT3USWRJyAzcOj0LwhPmL/p5q1dv2HkP+VRVDwDHsrBnqhbc5dmi9
gHVemO0REhhtf24BAgYoAjIkDxcOiFK17045re3C7OfIInwJ8MMvoO0GWtpWESlc
HVTLCW0jr9SSewotbD3eDfgg0V+prL2XFzfGKPMA8ny49ImB6+O+OQ/9XuuLtHMI
7LGYynufWXvi5lBhcL4OdvKy+FnPB6uY5MkivnVP2+5xJFEozxRcTNix38iDKtuk
jQIC87rK+Rvd1DWMcLAqe7U5lnmxpl2PZk1pLgwrec7JRSSIO062Msn3ymXszyyl
uTVXyrpc3XUdOh8qhu/8yNvIjy5cm3s4pM6iDmB2gzeZxSlglv948bQpPMPumu6c
LuJlwSgbxEYi4s5kHU5uo5GmOOw3Gfnc9UqXS2MzcDgdy3oDYxHPmX4q0uKYMblt
qF0JCmR2lY7dph/Fj+G0scH7x575OM/NiI5rXEK7lRxTbp8kTz/dwqvtRH3j1ht6
SwLJYaSvu+U7irJfx7IpEGYPh7dmRTXEoP4L53RNIG2nGORz3Q7q/MIyLU+vcLHb
/TjO1DbA+7DK2knmDKGC11e0ggM2Mx0HHxFQx8jCAH10MV+tcEbmNmu7hoNU/50B
sxpk6cAnT5BRzYJBm37BB0HU1K2KoQQLDufJC4ThSCAZzEH6w9nmUUKLGUMHQnKq
8TKaIZqVSaOFSHLyZnIqjt66btEFJSjHD1qlR1fvaK/LheDarVmCM5/PtHuH4sRf
qIFECMRhHgpJt4BEiAg/smDLJwErjaAn5WNZeyWZc8Cjf8YSUTj4GK8ulgGctU4W
OuJG3+CErlMSmbvbqgTqndB7sL0aTZk4e5VrwRDfu6RRR9Ng64+9yFwPQ3KCr1oD
Xw7VDC2EXBPOGk0xCL1CAqA2XZikEzJ59nxIFfeFTIM8Z8ATpWEju1e5hPD/L5kS
Waf2qkVLiZdbhJ1hHYNHDEa9YJ+oMRv2y1/iiddYTacmqDoaboE+fo7N4fUV1g+I
AOqVU9RdAhDKPUSrM5WZj2pbstXb34PNl/KceuugidVf4qzPLMPVSSWEMLEEJk9x
aHCtFFo0bM7pP5ZyUO/ir0whegestpwg8/Kh7fjonolI+olcQoKEXm4m/Q1jbBu4
/cSMRo+ib4rirUAPBMeZItyxEVtReIEFWkmw0m+OXnFKvqHy9ZtG33X4bVyvNFGz
6jvL8it/BqFdbmy5pWPAng//JmlfjJVc1lKDaB5wcj9Qc0k7U6nffWOnF86gWnEL
vLpu8mp8EUCQRKRG0wuFU0VJ4lTn2Lh4tqnw4ekqzONwLcsZHWsYIfTdWnQw61yU
hViwuS3reAE0+/J9FimS+ah2gjlPXz2/vZOpAb9Ia1Gk4FB83INuXy+Qeyrh702U
Ugt/zQTvijlYNbW2kGWdfur01HUfD0E4VoSX69YBx0RYF1gvyHSt2R44PJftERRt
in7DxNQ1G0cle2J8L6eySjd6Q+9fJB+CVJExN0h9N62l6OcSBkC7fTM05S5nsoli
ug9O8Rq7B9BdofS0kq86RapJI6YLubDhRJzI030uiXxhYXVzbR5rQ21kqVjggnsy
bzdSEFHoRuL52KAOTEme08k6tlBWaGcqdizcI+Af17YwXVH45M82uoP5VZtxz3Ea
q/Y+eBkuttWN7qIzh6LZYMMPOJcMgQAab0mQKXGZ9jvmUUcuVtb3ojq3FwwZKtQ+
r5WhCmkTwpXdR+705VMEamEq2hQEO2yfPxeLIczsSblngwF5FohuAlDKjNVjcdlr
EcABndg8hke1e5sMD75pRCZ0EqqWkVukgQw1NEQeUcwP+meTGUukNsNL2fQpRp/b
p42K5t8aNT5tQc+T2D6dsI2OQw7Ai59P5CnQIH3CMBr3hmO3in+KmXzVGympOWqd
ash29JUYvIm4tPaAq4TzMB0Nwf6g6ClJHomzN8mR1z8kpTk2naZtOrTIu9GfOcFZ
Jx+Tx6abz2yXuAbAgQWtXQPyaVIQI0BEM3fhKezUkT0eXzveOFlEmtSyiuGyvuGw
s0Vi5RsDwfvMZ4ayezQqF/jFiQ1fUKhrIy8BfQ9GyWbCvxqnVCduWaYHsXVoWrS6
OqZqffMFVhTJhcMj+zGybr6zx/Sce7PW5pwtIHbt9hVtwa/H4Nd+b3e6hOX+BGWy
RRLZNVWLDEjmyyqeHod+2CzW0m/rukE2vpHucHKjiADlF4x1qqQ+R6pq9NqMa0Bs
rFYPIguFMGqk8UBoBWUjMn1eci5VPKezBALgcUf1zcDQe1zDcJOIHpkApM5yp/qt
HMx0AyRgaAOYdaYHqCRoej/dicJf8MQEEle4sw0VAa6ZYjHaOoxXN7qfY6VXEG28
TZ+c68rJMedppMoyjjXFWjvKOd7ZxzhSylcwyycNISDezipEkCMWxRB+Fb7D594y
ARjDQJOk91S9ic0eK+YzIMKmSuJAeVJCfV9zxIeNYriwwEsNCtVTDKLvZIIb4lqc
IJj1dZ0+NSJAWIbEOq56KRoMW2SH3X+oPjE3YrSXVdxKK9NGm9TYyTyK3ZOXffEq
OQ0u2Cc3LgUJvFYjooTjKhhkWuYuusJOuT7A5+n5KSUR+jMsCIBebJ9iz7ZtpCwr
0dcZNFPfYeuKWeo6Xva+x6gOcqB87fJjM/VEpiqNFijsnDOWYmAKqKZQMDLFwu58
hEPY0B/cNjFQRbHS/JWscXQShtdQkYLEWhgqG7TSkitUElValwD33C5jzdbIP4G4
sMb3SIZontrxz/IkOtaC7IWtX2/jf3XhZclZXjNKl7ZK+hs+aVTHA2x3jJl6jnTH
qF4waICfzSiiym4YK9h1JGuVk4uqUf0Gv+3PYloZxWA0hMcgZYvLV0vDFrDVG77k
wSMiLi8hkJuVn9k2pgPkNfILQ14MgUgVGhpD+o9N1Ygg4TPhf5qtzYruodqdayF+
5aNRvT/sa9qUfIcKpOCcGPCNEP4RsAY46XviJPzX0NmpaNimwK8/LhDNbVAt7iOP
vZBB1DZox9cfqPOQAe2KSCLBCoWnn+9bXgRpIsmdhYDatwdNsuPfvMWYcwXpcqly
EprImtc+DoMmBFKJZkbnoVBr4dxcO7BC0z8UMAQFl9QrdSr8JpkKeC0hzV4RFwn+
DYS/2Ub2Scwfattp+AdWF2MthLmUrUdHK8HgBFH+Y2sH1twV4ZoP5Vw7cyLU3spS
6WSoDhvbZF7dQmS5z8+lWrpYyz8fUKxo9ipjJ55SewQXsFYzAk/PdQSENFyto3Nk
aEyw7ChKH3Gr+je6lD3EIEOcsToi/Im1RXyZFI4Uemq/5xDecq+Pmf8c3VMQMeat
kAveXXTZK6dTzM8Jo2xo8nItRqEaKktWkwRHB+9oRr/tLFGf8VjQbp4DFC+Ha9Ov
OLVW60+B81Ex0Tea9eT5gbmcG0UeW9bCUIjMRG6XguPEl+2MAh5prxf+u8gdE7h1
KTWqp5VsEgiRcE4wQniRZw/Ks4WLiC9wTxErJpGg6j7YNXf22oivX3OqmNPqBdR/
5ewRRmoiUQ0VZ3xntWmAeDLXffhWz8oo6a7nGajJajWmxILvEmjtSM/6wqtenfQx
F25anqy2Lyj8DUMXOviNulupgLtNbxD8gWuWGfya03eZMszVnecAIP/EOVuMB30Y
K70M1wIXZSN2/KMxMyjTAm0GSBRXSmUgQwr5qMUCTuHLiNvZErSOdZzkGw6KbT9z
PCrXhlKhVwKpZm8m2Ak2OWkR68QctB5SWbOta4KgD0UtbMPgJD6Q38PIhDN4WjF/
YUJmrnXidwmpf5y3mu7PLvqTDHicKU4FCBSa5uZkAFEXjMw6UPVSuxq93C5WAaDx
pBjWG3zHpbfglj1xL4G3B+1+X/OTdjzoA8GGywdwhzOs/hUTRV/JgaqNpVfA+yXm
U9aGDJbekORvLj7DoMby8gC8Plwcq6htLzXKXszd9J+Mpec0RKLHql3eyFrLyfdP
HNaWCvR2LHrpIVJTqQCX15nxiUa9YdbwGxcCeGCKO3z9tSi1pRAbRvbOsvV/KDu7
+NADOGwaejrHo84AoXyIXDOu2q6gDz74QgoAtEvr2MZwtYWYNoYx1KKpBoIz31wA
fXpxAzO756ER4nhli0qmm+kneiX1ontuo9qOtM4S0YTjmKJwTVEPF6cDiFloE/bo
rBoKQyuF5FFFOOA4ku+znXONE3l3bYr0QbsRK81k0cFI7xJ+xU1b1zyfu18Wb942
qrDOu6yEGK2KF91t8MGwBx/e1kjbrU7XCMe760jajUcFiwvjWALfc1CIQwyLdtkJ
BtZ73f1qHzicdKKS2bf7uppWjOcYXeZ1SRR51lVBQKWN5q0T4BlvAsLOM0W3WEa/
HoWiet9wvDfSTFZwTHpkElWnP3dsHH4+YcnrXP5jSNPvgVhdxfYEtE3C4Q8coFHE
UvRHbgz0/UFazZX8IxxvISrPrr7orlz63Ndllrll3Q0TYEJrisvtzp0SEedZA2CA
rZqmONLCjVLB+vzOJiPDif6fv/Z/Kc4PazJmSE8g0041I7ArxweRCWkzVLM6lP+g
SVaNSPIBQTQYgJEs3XPZsFMHnu9DUuM64mXKoTOZZxoXV+1e1/pI5gfk/Vk8cV2s
E4OVOKbUgpfdf2zbuhglXzAzeGW86+r0xgwoyP7KDVN+T1pXPJzmNUuIh6CLlr9I
/7Hyfa24R+qoJbmIU9zneAywD1OpUAG2iwceRymqEagYO8EY/CM7pnY7cPF7U+I6
Lps4vbCP9plOCRlcqZuM1df4KYfa5K1bhb2cZCMP3UYq0eZLveTb2ebaewkYYZqQ
bWOtdk00/K3Gcb+rEcTaN6hMIVtRIk5uiAd7IyH+URKA5MtlTgZZTGo3/Z2yUV1H
Q4TtPtiVVUSG79AFJ8XH5VxmPGbIwUFHFOiRxvwkWLud4fzLnljJ3x2MWE04Z1IG
tqdfXaHMtbLxQdeX2pcufYyMRSLgfK0hwRNTB/7K+1ku7jInBr2o+bZvFIwRpokj
ZDa52OO926z5hbEs0DZuLApMhGYDI8IHgatmqoqJXsEU7A1ehB9t57G+lr9FKVsu
NRkFXnvMoOKDNLDphDFRGam/EQ5mtrZUxhYHdgVLqS/+ji/1Jh+q36JaZ8pNPLLN
D7ZkGLJCVhPpyAMCfkct6iiIjsEadVC338Ppn9f6xtdk7cZFuGWP677OVpajfmnI
em1vB9ADPQ/53KCv4nBwHJhXXN07dHlWOOKMnJ2DO/WfaDD/eCeDzi3o7swpqIuk
KtfisGu1U/B5c5qMNxA8QIHcoch670x/cmmW31AaRESAisgvhWU/2YLXixvb3CRg
WwSlDunVeWoFbVXcP/tV5qx4SfCc8ZZjM0L+P1V+Hs2WyeKrThrIpvQ19EW6FfoK
TypQV+r65f1t11yCH+q1ION1UQdnqMcSEY6idzVmmNLosLNkdZOMDRKyzLPVu3Fk
cVDKZWP2JidM4Eg3PRCHiEoygimWv1bvTrqVSp3FW6j6r8HLJlUaqhfrU8MDOEkM
bbH0VNT4pUxOFwk5kyJlchUlii/359q/sk3Vn32Cf0nUdsX2qX5wavavj7TPAYRh
0L4nvqx5JXwh0KGYpt4R8kKuybhdii0HVX4ebeiWdvvMbDiV0PhGEryVAnZDiAM9
yN6UVEPRtMfINbOtYP0ZjERfO9fLEoMm63gYLan8Sk2NEnqltOCM+hbd3at734w8
PVPWrKzU6NhJgbJHfCaJtznITlfdAK4pgp/419VIQyb4tI0QbwSn0Z2xFomjFBvw
ioxyt67Y/yYUlbOddA1ysp4AQpn4Al3Vs8nfWHUY+mXgizysye2TIdrg/Cjq1Whk
IB0g1PXep5/S2dqkv/h86DoCjkeQAxL92Ak2/e2yWtuy80PuQZnznUaNM2lXUw2y
N91f4XMVQZEDI4UgATSFF7he4S8m342ol/KoMQLmnvOQ7/UTmuVIOPcfopOEycEI
RiT9fDCh6JTf+hUVMTG4jLVJ3VrTw5ft+wImn+tcqvmJkJ2iuV11yJbdloud1iVJ
gupnkzRX8JiKKiWeVLjTDYiekh5azpHZfQabs3KN8GVB2kpCEGSQnau7G2kwid4a
IM5zkXYsI3O3WHI6Tr1imitST9XlcwxN0BmH1WavctXrX8yCVPINsK+2Tsg996DW
f9KUb8AbnXZSjH/ZHMCEa2oZ1NLh55c/DQeIXbvQhscLUV0ZNmMk70HDw8SSDfvj
TVGmIC4FjFTLVqUQzggm5+uGWVpx7FUO2sRmPh4YSHM5qmMZCEYlK4/VMsVOJVFz
rPGvEYFYgA3SHywg3ovXN4fmCHvhc2Ql4J9ZqqjGzq6ct7YNQeKU8L1NDUF2o7Bt
cPboD5tOrgWWV8bJynT8cHj4BKg/nhO/YnLo6bMDQbRX68dQ6ncKIvOQyryRYU6/
Lgnr+K776JTXy1NBSzvy+0vqVz92IS9b3mg0GbgYqKcd8QpmL2Sn4Wig5oXEAl8I
ewBfgcMuNHhhhKZDpcXM7xb7cGVvTjOLIo4Zey4QQDhpT6N4illBpBqVRmKsnFAj
yj7HdEJkVYQDb/LHJSd2faHYvanSO4r5CrOBaoDjrm8NN51Um7pMWn4FwY3aTK/t
SS47LxPb0lp6exxLiNeBE41r+ptDSxldNjAJfX5VEYh1gi5HMiQ47CEDiPyE9BtW
SZEEt/KTOORx257lTSB7s3lv6ke4LzZT7jKmYAEv2JuewHz3nPxVzjd+0zt0bcD3
NneNnz1kXe9SBIk2fvPqqQQg5PV9+wSpcrEb5/Y6VhUgJfZxSAOT+qZmW9vHuGkr
jlOd7eH1W8+VAI8bIW0fYD/Az1/VgVAo+yTNOUsvDdnE0wzK0EB/df32PsHHSLcE
TjvezxU5VwtOBlrB0aTFz2PVW8+zEAlaV1ehktqlty3GW0jXFmYbvDtXZ3uekBFE
+IUifGkLm6rRnXfu4c4DuIzDSOzDE0oCQCRcvfMTJMG3hz/mbT/r4xDy5C+r2u62
4voQAry5sC8/fPUZdewPvy9TtYx6+n8D0oWXU4zaJg2T+ZM3mDCnX8AQEo9Nvzp3
qTlRPT3isEz/j8dzs2igAuhBcVsZIDK3v9ahv5otZdjhSPvCxikRRtLBODSswFVD
yxlaaJaagOBkuCYAyDLOgpAHQ2W1ZPZPreUSb/Uc/ySvQJhZyipGYxie5Zj6IgpW
BuuVG5S9/dZgbA7Uu8XDn9Cyw2CwkDXUD+xHKagSze083aaiANBqmjpDbhspAPtS
sqzUvOFUnSdgqNmBLQDK9h7aLh6z6BD/66wV/XVI6q10dzL8Hsa4sa1FUWm5ERwx
6jXds9s+4p21ZGl0Qtp+s1p1h4aFRy6cpwl6bTZQPc+z569hNDqMH/3YDJn2De7x
qmh7IsILxoikNTtzZRdQRkgohaJiWzG0L00Vzq7Z2eAafCt+WudFCbcewdu/gtRn
B0l3hFKXGyWGsYsfiDnSijuCpXLFBJTfFinnmkkFmRNkSBOl7D3Y756BkcIQQtmH
ZAROP5P0/JOfeX5hQRp6fYw04Kkj7/y5aRHFmxS6vwcl3uCh66HeVDP2Ig5l6cAG
3QotFCEdkePKgm7SBa3Lwz4HCERu4wh8IOa7/vjJutAIMmp/4lgGnZRXE1OGyj4O
kjDrOh+JBY1gPwNBT4X3MvRogU1O1S/vfhBUr+HK8aHX5z65fmmcD2a5OwOS7wi+
zo2r65E57uxMBlqPdJladc64gT7UmbqF4nf11Mfgnyy31siQd8iLgt1GUrKqYMGt
szqUDHaJRBel5UwjXiXRc0pcNis+jQ8cCLnvRQjRiK4BelN3Tdu1VHtbsf4ml6Il
UEse1q4pVaPxT/bDztFja1It84W4nm6zwsuIsRAUNOtBFDIDf0AGgMB9Pww+TqsR
Smb4Ki3snzCBweUlKyZqDdqc91b9O4rMWyw6TJUVgRCgBNnjYvMUmAtjs75HINSD
71OIsPYB741klABogtcbN2oh9xcj0BjOl9h8Ond0K+/0aemT0Ucq3m0hI20+QhEn
+1IcR4JqUKBN3Oyn09wtSQ0ut53hE3FGt+oTeT7be+VU78Mh6KTtzNFML3DwG5qS
8RMTYyQ2EQGBU2BEgSWF08Aros7ak7iTQirmj226sItSLciT6SexgPn1GhGcs+ci
Un3GRME06xNCLFOSPmAHIiR/mF3PXvkf5CHeeAfkvCFOPCFECr8AuEDq2mwLRKl0
Tr+gfn73hXTh99esYQdyzpfUB2AbrERpLF+EK2wD2ULz2QJ9W9sWahcKjIQg5tab
N2YXVdLovSobY7kaY+FEE2lqbrZ1r/COJ2bX435qhee5eApYRpLJ2cDGuVmWF2ik
gmcO08V1vTDxUtyr/XcWsM4x6JLAJrfP6srhp/S54i1fcGD0zGMVwYlh/IuLPDf/
v0AaEYy5wUcl36/8xs+1EuZOuu8FI/LPc6j3RZ4mOZRPz4DfCQp9vU0BExExpTXZ
9IQQ0v9jUZiQSy3e31Mq7MGMqkgdc4lPLSkArDOorRLmmPsK3uy9CPnvw5Odl03G
I714Lqxc7U166yJAS3GDD9FGp9QQe6ivfc301C3thWEsV8umTTMUy3+E2WP/PCJi
pkmn4otgwxXMa8n8ptX/IReGtRIj8kuox9R5bId7vxdeJ15ZBSbjSODUj4B7eXyC
OT1ZbMxIyBxys8gTUYxWSD4VEOluwLpLTzzqwdzbV4wZsO02EDp0DlB7Yczg9cni
U/+EVgku6dLgJINCpljWuiUjS1hOrO5VweVjougWo06Tu79vpFoZ4iRrxervuvkc
6cMh/g72Sbz4Q1NlSQ57rVDg8J+RVAqMk4hwLL6CmhL9j2py6nUDXPTxBtbSzNGc
qcB4od+UOoiVzbCo5TbrANh8guBnIkhwhhwQjVV4QYo2xNP0vtgvhM7FJ1L5trhR
j13nuZkIzHgVd+2E6UpQQkFYRR2u4bXikgh8lEsLqC4qkkvh4DMAr8tBmVcIj1I6
Ql+CptV9AmZzhg99UhscvqKUDZkDL0jylPan5C0ga2J9KXPk38wClTTUMszBTiu9
eTVP60ymfHnCMK9LUivCRP+KWzjFqQQ90HovuWGk+MDe0ZP01kib1HJwn99/N5x5
Adjfk6sFGXQqi8x6M9r+ecixuw/qw6xqP8AUHCrTyg6sG4SrS+BViO/Ksm/rEd4t
kiAoskEGyZHBzzstg3Nq0rKVPe32hCBHPUxI1/njYBjzENl9JayZ6rjF0GL5SiZg
v0wK9/0lJo+BcBnoEZjjS9mHp5xss94KO0uMr9cdzst/zkhXxEwfqUv0+ebCwRLk
Jdc+SQHcZf5ve8vplOaFGY1UWuNKYQeV+/AIELx8SMOefVbMEnYeKoUgfefu3RZA
4viBlIyDWaUt8TS2Fbdpri6sJK8BmDkVNVh3mXRonhiAQ0azVkFO+C5KWncfes8a
KGXwEQXa5dh1i/Pya7af/9Ktzx1bitZ1/ZobyZ2T4OoSQxKb7WlfTzv2UNAup0Xw
YhU1Qr3YUkeJBYTa14FAqE4ks6H6CMceGxjLX1tmVYCEuCiPZiK1sNM4b+YXQBPv
toYMtU4Z2csnOysKPhObmk7HUwcs7BVVwiXyz7IMwqr4KbvqpSdgwY5aJ5+0Pcs0
aUVjnqpQjN+TLLsuAiBjChZLvKxCWxr7ik7eeOUGjvaISqT+x+BkN/hIkAedyWTj
IvmkqLbmx1JrXKUhcQjcWozZXJ7Csu3QxDHpL+7W1zXwPVswb1euAH2Cgc2kWc/e
3WEeQrEIMG29uHuuPsDjF4x0EU4u1BZ+MURoUCZz1KlFnv0mlyzDC/YXj7n56Pis
SBkcfQzI3wugTSlGUjLOnthbbYbIlQh0Q3Wd2FqnJ5AaWsSJKi4cJA4stt21BnfO
n+9L7W42xFQUVUXHUmh0HjeKLQqi/uWDt4Xlqrvp/nBB4QufB/97TcBf68HHLZ53
1uZCUJcRAI0e/64tR4MkzJo2CmSfJj4oC+GA3ejqesdI7pLBTXmKePNG8fc0tDyE
vj/4wIJljackDrnZjmaKFntpnKJ7C0s30XGj8d6vKmdoCBOsA2BWKGOuay5kikGI
cu6BkqamKFbtOrVhQ9+4YichrU9rIwril3eR4Omy+Ltzs4/9P4wBwvQlUE8Kgqrj
yRehw5Dm9StxAXqjM+wnsvrf72G+v82wTCcJNYmlKRV9pYcDW96JDwADmrNDWXFz
t6GILpxKBilAao9JlaxygA/V3+/9ccaYQnMHyxZg7UcFEg0qcBFQRj2dKld1rHye
nL8pJgZhucRnvjw3BxSO04LgNiOEzcqpwttVenwRzLCmnJqIIOjxC8hYctBjfZW2
dyMEhNNU+JlcS7bUSy2Mo1WvLGN/qjclKFe5Vttx1/7yruwy4NWdWbFE6GOuu+nR
Rqoub0jh+rmiyFOjvcg5QGiGYvuyeFNYY3qEFGnXkVc44ggDhivKBpR+TL1B0zeV
yfcUJ3PLbA/7Q75JRyX2LlzvlEZjiigaGXufvmjMYev8jabHIChayFG2vd7CoZWs
iUsuB7YWupFqy1i+ICM30vfhhS4o+eVTcGcdLSkCwCBugnH0AiG8mX1IrXtL6tL+
gTCVZ3r0fRa6QLwLeePL3EMSpeeFlFTLt3OovGf7hjXZd3zbdDEprYak+X4BEgNw
f4W/Vh7fu0yFGO1zjAKWEvj9RIUBrEAHiZhLzZi0XJ+CA7xn8VoHmSXSKRvFi1te
U0IDUUr/oY+op/MCpxn21XUH+7key12HGLbX+YE06XCtwGFl3M8GinpMECYIR+y5
nLQaPBSdwGU2ycZ3vVIZnOjC/8LrglCYNRR4ddRCo+JbMMsOhNs3CTzUbq6ZubAR
S7iJVgJeJ99JriGJZzumY5aiXgS/njJrpPX0W0H8yIWizp4gqx4edLbnJKnfuEgh
ezi5FksBo236vvBYz/HvldprfT6NoURWK+XYJWjqeRNbVwub3JL8FdoEaP8ogzv9
lVLtYkVg2Q5p4B9axu9BWctYsjrJn7tI2l5UQbGWR9rOFu2EZ9hTJr2/i+/onLH8
e3Va6gbWtPpzjhE6JdJWnFtei+RhAKQEBIZ5crIOONA/zTXDLj3AsnQhr7m5gQ+x
KPYeGed3yyH2ZwfcaaJFre1Lb2j2hILbs1tUInbHMbOMNMPLAsE7UKo/OH+ssw8t
O0rzO8ouzPcSEwwuYbaZEvYVHyahKUKhM8dE83xsBNWJT3FwUeJ8f5W6mC16zA2C
+VIIo6VYiF03RgIzAKfTyfq8t6YnKBqdoJgQtHnLQFTBoZloC2zFa8JtgxgD0aXa
Q7Y3xv4qCn0Qn1SO6VE8UCiCO7yakOerUEOFpl4ZFx7TbVbYwtmKOcw0TYvzk3K7
kqn6oO4+v9DK3HxvIlrWFxUdKcwsNtCF1LAfdOrf1sqrdZnxvRjX4/EtAfvyMUSO
qY7ioqBC04Wiq4QieGEZM+MDc8RrqR9IZ7DS2EES2kZQo3sIUovJYNoaguk8BN4z
LdOD0/ALHhxhwv8sm887gFBzeKFoePN5s7vt10uADa9ooB0jE1PE5dIW+3ST/HmC
Q8ctw3surpl98nJMXAtQjrLy4bPnemhj4JV8B4JSMUMRUvEiol+6FTVcs7PGLCHk
jHRcfJV9BS6IgYTRnzY3Ye9XbjmaHMBk2Yb0Aab7VzCW+yX8BRJ+8J1FKmf+yMLY
1FrJI1sdjPaF/rg8NsmkJA116Nc5jdgcwzsyza2VmQchf7EthwCzIPtW4c1EKHAC
G+lT90hxLdImAnodv6QrpUQj2hbIeHaCFGlvXr8AB7eKio8vpKHnHALHz/d8CCYV
wh8P/tQ1R0HQw+KvuuFXpR7Suf0XE9p9VeajpVHINL2XHFN68jePSZ7GpISoBePV
NJSGw8/LyRiCmy/XRD+wEr0LWfHChMOMfAI6BmJD+3V8/q4BdWGpLJpbvnr4yyDV
tLBdTlrmWR9FrCmP/8O61MF21Yml0Zn9yngGh6r3AXgDIgH3hyQVUUVBCghjWNAB
H525/EFI0hbfWFGBp1GI+/YKaqaVQn7dhQNJXUOm/x4SgSqaLA53uTamoNKDCjIE
P0fP3arRBoenmES+j0rd5kFrQZmVJTnmRnerc+1ledzWaHLv6zgkUSkPSjf89YHn
olPYPBIQci0Ua4Q8lMh8nhcbX0vkf5d9hJEWbucpSuohYnm8X98TzR/6tAvbHboi
zSgL/J12XvwviWtfkoiHts9yJd3+tVE6RUEaDQcDX8r20BbUo4EZFu8jMp2SYznU
qcPfAHnFHrwKKzi2mdxcrbzjkTGULF025AcUPJdutt/hofKo7sIvEsCsOzWaf0Mv
58lK/0KpWiDcUipLFd29t8Bl/mJZHP5ZmkB/hJMfqAwj5p8pbw9CHDI5KtPf4CFw
Zw37Hc2XgDKrsURpkkECwMklHb/8/dFyN0vYpt3rju0ExpnTzcX6OHYMySD9PHlb
NXI3V2b/Er6NZM4FlYAQoXavw2I7T+nn+q7oGQP9xmTZ7xX8VHy8d9+KIEL7s0yZ
UU4dmABfMa0uvud2fWnD5EDHjwVqIqzaGBJvhOPn6uxqdaqAsMD0GJKzhEaPNbzI
R8ymO40AHGOsqtX9dwkPk8NUJQorfnYYLM02sPVOiqNXNPj/HbdOQFqhT7ibVEb2
wP/sutILJryqwED16AZlMrfnnl02NARVEdGJlZBidaSm87xWbyge+39JLkP/1Xbb
5kRoWAgJjG6LnSKzwD1jCRrCP1r8eppWcoWXdL1gx0ul5MYaIrZtyl9TKy/XaB2e
rboI8hSQqkqWAC0fTraCWUrVuroHp0U7mtKk4NvkexZ3NyqMjfd5fLDnH9vjK5Z2
Hp8lm3/Bf6Cnsb2XmMmZ8oZaFhv3EbqCNtPDb+CRmj5pZAVfxk38VEQT7XlRm0sJ
85ez2kMR0PzaCRoOK3FGwxhAAAP4zxfEQYdJz5iGS9HCGw9T0L7fxZP1xT2wbYuY
JXYwXmmzLA0Xo7E4tVUmrzONDxz+b2uqE9RswpX6yRYGg2U+/KScTHypn8nTSQ0/
ARiDAeHkLj/Z2eP4tKpvOUDckxDnnY9wGCwUiK4neCk3CeDlC9noPUh99O+crkiD
tDQjF44ql3KgQXmeEJt5OWHwP5Ew8rlJHBWIMfmYKLCyYJWVNANMjUewbW4wLZBi
YXG0iaihj2Psv64hQ4LuJSOPMwR6VIw3R0hHPGKMyfVkWemvsJM05h94jfy2pOHN
NfFPOwQHBmRo9QVcgFtFS6PFBIS8T5xSK+JxqUgiEf1DP949n+tZyMHSEul3y0MB
1F4yKe0VzD7B5TgQzGU1Yfu5eO5rK/0SERMvTHdv0JT9+d9nE3K57/qPSZQU6UYd
xDbt1Jvhz7IQGkkhIrV0tRJeRpkw3cfodLoo2Fkn+bcdfJFYQOuPlTsSVSu79ufI
/Nsm23s+EU9xOsQUkcbfBNUjuqD8fdx0LbtbjBsO5g3INOJR4rqPpfXs/AjZ29gV
WlHuaQRBmzGnsIbL0MIw/jHWhGc7I8yr904ox+JEngisk4z21zSdVjYEoXC8iMg0
oSV+yV3SfRWgcWVpV5ckCylcp7CJRTbxl7Th073kHDsljmwhBdQCSygPKSF2RKRD
cQiCG7536FY7JMZ++OQrY1X4hcyrD7Ho9qG7PXNyyRhPJUE5WPG2Tjv1s5hyR65a
7oSIB4z0cWNyr1THAIwn11XOS9k1z6cje2DgLH8QJ+RhKNiRe1F1jc9YDN/ObSBn
cWUtMdfvM7AIgxM3inbA+k9Z3ppPMSrnujMG+Iw0GXZy64yXmcfESOwJ+iazJswZ
ly6hRg/6UwDEuAMatCBmFWjcIK6uaVwNR9dP4wQkn/9uZw7zV7ZSdEjLs4DKLGvw
d75fxm5iDGNCpkeBKVB27QunG+LEfsow4OfgCRQdrAhBqIEpzaGzW+1Y2JcmB78g
XNtapRX6DWEDbA5FlbgLLes+DQARlu+VTwijoZonsU/Y5EjZYogqmq5X4w7xVlj/
t5iOiglxSItPkeIMI3ovz+8GiVwAhKRD8w+24FfL6InS07cbwvAnEZCOOBIRQKgn
X65jR1DqwKjvTiw5L6ss1kWphE0hU4sHY6EvJj++GHtDf0Jj7pWS2iGhQUfax4Zl
59HkBX5eQQCP+7/tZ+cw/3d9BWOWlS7MophQ6WbcWkFejaD7TuW8xmeeW7SjmPvR
x8IuhQbCHXx9QTuiLtSbpA95wX9cyfcp5kaTHpWpsBwE9rTjhNNjb5Pn52yNquyQ
yh1dbJl2ZlxZ3zapuXR3/Jv9TuISMcRQjNRNmSP/BedYtk5IKtxEs/NebOdwixVD
2gIJRGB0sDjLozeeA1iL0v2d0kLEpUN6VRRtdjB64e2oeJb2Fwv92Z6lWEpavHuK
L43bwYe6miceJwpgRWyNAHcslzP1+onH4WoV65gfH/PyJj/NcEFx1YEgiKEYYM0w
g3a4RCiOX0fFOLpYSTppbmdXWS74TKc3F0GLbvJ83M/V1RuP68i1YSlJo4OWb5x+
VCJC7bNUB5lxS7HN1AnniN/CobNONvETYTkRZ1tYMbggJIAbYnoIMS2Zg8mUdCrN
3Y1QZQOxX/5h7XnZIwm6ijlcGYVIMCfiy4DJVGzf7fMZuqjiY66xLuaG1tR9wnWB
9CrP9o+2t1eMgl0oGcOQCgkXLGSizjxswo2OXSySFjm12q0Ox8R4pYdDt2vDvAsf
8ae82WT6BjE2J9kqvu7qEM4YAEZIAMr04UTwif4Jibs4ygXmW/MJJK1GtqQwn1z5
LsSzdGTh3wOrMoldq7nccm8HOXEJDouj08EsSxdBTTVzWPCMaAWBwcCUoNbou6BW
/nF0JJczLJY8OoN80QafrptNFLOb/LgCRaMvzOMZDlH7zc7HZt4S6dorgVF11ml9
BxKNKnZNdluBlsNKICEaSk+OBU6ospMi+ifonP+zFyMJDI/dVK+e2+n+yFKGMlRv
/vnnzT6amaiu8GtBwCFxQbD2UFZHIVLXsTNAnOx6ANB/JDyhmk8GlAQO96dJbs7Y
tZucTwKvW6P/pOUXcjKVL8k15NNcXsO0NXxfLaqWjVzrK5xMYA7gAaa4CPHXMA/v
DkojH2A+C3XRnywg6HA3z1spTydKlBgxJ5v79pnVd74gaFFp4KDjrGUq1PXv4axS
WDuc64gM/JjccrmuL935pAn4j/sqjdOeIJpnnjTEX0ek0aiP9NsZTThbM/b0mFiV
iK/KWOn7uMA/S21RXjPgtOjGVHZBN2nWe0fyMv03E92jKd8mtfwZhh9YdCVtN5vm
Q2D89VhvQDurKcjO+8Ls+bqvxoS+vLWWccJtgM5vjW/tGl3ZXbE/i1RHJ9qpwwwA
tmba+VisDDt+Zr8hWTeSwP5v3OpqFDiSGaPoqkUG6DbVFf3WcGwrHmFQHIckpJNO
WhwtdqwVV3d9Ybju+SI5AjiG/Vvqs8JxA4wCwQ0BHgdFV/Wbes9/y/Zmn+G7Hj0U
+ymI1Ne5JD1Y92PQHzhTY727KYJr9ModwDQZsd082y8u0c37Y8fyt1QJRrxi46F9
U7PTYIQbsfCQt9HPlTfmrASsJkNZEjXSeBRQyraoqdfMZxf5qml3h7uh4WMxfFrT
arozkT+PVrmlUlMQRtL1iJU5aKdXkIcHBRukqCV1uOIEuMfyXuflKTLuuui+OsZn
3gSCyZpNILWhDJ6IzFiWUkxBunvQHMFzxLjNs4S7dxYV3Q+ZKqaVzEbuTbwZAkVA
pQY/4sjYZ0pQgPcgCxp4wGqa5v/02oIYglZtjA261uV1m/iDBDIeuAcRCdsP5MLK
ru1/iZuAONz6NQScQ53XCHwo4fKBVKd+HTsyPK+XkvEmLKxOevC/Q16fDjWDkyAi
ph/8+9xaHDHrDe15gmMOt6cNPp7/Ea5/zT4ixQIvIG8gHGe5co+y8mjZOMygDoLj
4lkrxYedqdjHzv6ktGUoK9MVnXldLBkzOMol2VRU/NJ510yl97qGOYPLAG8UJQtj
D6G736qKyzHfO6fsgoAZ9xM6P+xxQ2pzBf00bkZ5hhdHQ/oaHgaek4pbeBok340x
7JKfvFKLkTvHfwD2lwPFGd70VQh7O+TaFxY0EVsq8Ss7PcwrXcj8MeHJ3A2CFbte
Sxyp8+DizROavwfakLRJFcyKwQ/F2b8Reni+zz4F/llfd1mJ7f2NR9afxVctb/7Q
RcdlU7adNGsr3/uksVza5BiwoStTtzhPCdpAHPgWL/GUXYX636/FgA6NuAG7npwD
zvko4rEYzfEu0Yva41SVsAHCYXzBRZaONkZcHk7kU1L+aBOH3ThtmxPkF2l6RGcq
kCfxA96xpi9zfSL1gnl3CWrI8ow78gWo1i8jcNEJhQE033bkNvr2/DNHnoF5LwBi
cTgLFxaVk6T5ErwStWegUB9hydo2TzWSBd1D32ZnsQ1Bw4N+jPgJk6KZlOJAVNh+
AH3opFnk4cdNL3vttvuOf881DTKQwUFCoZr7k8REZRP0VaDZ96fHMH7LzP0SNPyj
aAc4vWQsTEbjJV1TJYd9V4Gx1mFymSVOjwvw67cuGP/K/an4mJucmcNBET2lUh/0
sBnKHmpshmvBKHs8P5lIOvOtO11XW03E7Rdjo4wvOBuvPfRRbI6JmcVkce84hHBB
/b9FDRou0R7wDOYYesUgIX4ZQ5gHBNpneX4s1AjmXpRaE/CgbiY6Y+lNcNyGpr0O
CJjv74957KvYpWN2Y8zi6pXIoqw+vDliFSy9Ob+komq6t6DsM1IetTWUjtl5lF1Z
Uxp2M9QEzgmPayrPg2QDzlNQTUibDv6hSaQhrBUU9+O73xFGFwzdW9bH/kXfy+0P
zKCPl4nPCarDXnaea3NIfFCo6HEx4Owy52BULlllGOclfxF+kXlqYPIkSnjIxY5/
EoS5yF/U3ShynBiQHn62M3iFC8j7jN0kVoBDKtxRUXGuiB7lMLUmDbCKCKdOzeoz
0y99WHfM+2wQw2UuI8W4FTvfLWBHc8nNYWGIeCWBNQeyrV+fnGdVOTAtzY8Ehnbf
yA/q3xrmWS4+ow3xv/qg6L9lsYTWi/l5E6fJYHEy3dSMH83BqLe12+khEl3dIkDb
1uDgg7ZF+2QGP1qaQC6SZsFtjuqDBnmgtHZW1Exk1yKI4yln+fYOC6CUar0P8TfJ
+8otLA3KpE0KbRMBEwJ9bcB9AONyZcQLABNthTAYqRMkaMX+qkZqm/bLVA+UC+F3
YI0Y2lQ7YMtyRFB5iLvGaefYNM9aBVVd3/VIkLT9poVhIeZxdeFFf1wQMxI4J/pI
5Et1ib/ZU4NW/JMH7bajhR6gWBvLnNPBhcyjtorhKcW0Ou49P7A+2oROnBRD0T/4
6FfyuSiPBNe3aGrrgHIslUcb3AMh5kXIM7nLOUYDbD0UEzYgEa5La9ihg7zGh4BT
CdQCdCqeqEdX6wo/y/HDU0YTagBtlma4mHLZHahjM/5OqAoBzYK/K4s4MsX3VMwZ
hnQl7cpJc2m/CaeAnq89ZrUmWDIogvEsrIUI6U6jRRWbhHCujp/UlyjZmmKszVRh
xFM8eB4/JoZ80BRAyjOpSEdmrLN8yZgZD13E2663EDzHwcu8RtlotyGvD7+IIa3n
mfa2aIsSkY7jr7CVso6IiFEOVrDijRbm+iuVMbkkZPxm+KctEeozsmIjpIRqsEb8
jQoj7pjFtXUHtOxrf54t27oep2dsbtSEBAdK4X3AQtY2xJ6JibqEg490iXbqB5L2
+Vh6Ic22C4KpLs7zwYyobyHg1ed0SHfrhiq83+cn+eDradwi/xoTPtzeTcysWqRL
lwqtQH+ZYa261+X7VB7b0vK34qU22C70cR+ptvc0MoRK1MoZszL9uMJI2T5NYbU7
9t6in8vsj7YEYklO+mqN3PqPIkIpU0dftD7Fi60B9WBa1SyOufSIKyQE9wx8/L2b
Ms9MSdY7NkXzFBxnkmcgDE3LY5uvWuepgs0qH7blLDYt5Jix2Wx4H79iECEH0foV
+UodlgFKlFXVSORIKRaPkgCifKIM/bsAwk3BeED3Q+MISdNQzbrnBlqgRyEhZBtg
ZMkXc7S0GGxfBYN37uXsj658UtD3SFCqt/c+QZMM1hHkhIwPJ1RQsTjTwW9ODzj0
Vb5+gDQTfPgoss5tSkjuHQUEjOzP3hrtDqVv689uhi3sCsZM9WkO5uOjcJXkfPHH
ntI/jLXPBZXhdVHyKeWekVMvSCgX8EQEyeKGlnYu9bXcTFJWxtyw4x0XUBdm+Mzb
a2Pk4HvQ+0yFLyUgROZ1/6Suo8krgJtUdkmGd/4sjupbBtGDkOoEg0Z7NOr/KTRP
5ZSF7v5J6ThSWBj0TjE8LFr9Gu5zwfOikvIs3gW6WKXZoI+YP887wEXV6T9GLA2D
59kvSIBcmnvQpqn2/SYIHoSBVdDEMkx4pc7B/10BSA5IgQrMKcybA9z38rsVBnfD
L0dLFkER3v6Qsl5xCDq1KSNeAXqXueSak30F0lhJqsv2rYxSC1j8wW2GyN4cbpfm
8/asaLwEJMo1JJWd9UDOrNDZ4AnNQ5DuXDkmxs4DzvMZN7R+ukFy9aCiHnxBtp48
L1yzXejfJhMsqVD2Q898PAgcznBag2wIlT6E3qUB1Dog+zREiFlktYWksqQlSDRn
jQyUFTfXAdWnvQbGrMW3jnDoAbf/WJv5H3verFlpUkIdVMBDxtjIidPbdBRRFuD3
eZnTr7k74skpf35MX3LosO8xOEn/PJtUcX1AadxRAms6XPl5aXF7IGOz1lnNzmYc
Eay4QTv9+HFb07IOEx+UWCaQm4FUI6uzsXX6iYt3HN/hgHlf0Eh1UCeBWk2hVj/j
aQUZ2HjeA4gmDx0xZLq2F4FUuhp9ETaDSHjF1BD1eoec9MVBwkrymm3JTqEG7onI
VN7nhRuvsMPEX4cZL6Zv9+IX9/KZ14i/B1e1BvwRp1pQdDE0Y9+SdQTujvNfq6VC
rAmjyva/u9lm+XuWoIiJ0GNWOm/i3e/WPALMDC5KiYjt33M2RrlQwvt1iQCLe3pb
cWzkBo8tdbFcUhf+tbyK7M+OWUiD07aexRMK+8wC+NWjV/xLnd9Ufz8LNUJ7tWfK
IydOZw+YHmBnOQxV0VssF8gNJPitobE4z7IwrWx5beZ4xGKNPTGRq+sZ3P4fKheB
vds8rStZKPv2VcmMa6St3rBLNHvSdXCpIH9QoAjIaqNPzBYdQZ3y8KLn4g648Tlj
7oS7mFwr6FlAWq4dRvYW6b6dhHHFym1/cy9Zl5jsqSj4x/ku0MC7OqCbx7lfd6T7
9oTsxP6+1XrHwlKibsxKJjNKZdXHm0TW6tkpKgsaaZb5EzxdmguYejaZVkSc6IS+
ZjVKUDv1ZNAgAGKr9PEBJrc951Swz1RloubJ78YAXFMiJytXy1qKBW3MLPEjtduy
vX61T397UrJhEjCFeaGekZqrC1wsfjYbHFKDpqXUNorF8D5g6Tx/dE4cH67fKwv9
cZABKHAABHGVeAqkULNgIyfFmDzQcwNcQJdrLMnp5/NrZm3bMb001BQ17ufwttzu
I79F+m3E0C+YrS9lv/Rgvfkw4mQ24VciK5mkEVieNi/wq8BsIBW/Sg2d2HEQm9gd
kqmHqLX1RO7juJb54wwloVGjXT3In3X8SR+y5LpZxN3IEjcqtxPD+PoUtkWVD1rj
crgHovDrM1jZ6/4SHW/0aSbEn/EUiKqyNrbwjM/gkENLdC3EUKARN0CkISgIQ0LL
xmVZ2bU+6nV4wQ70ttmYWrR62lGp8jfvLFNRqjvBOOkPdkN0FvJI8Hyi+FXmoU+P
a0+7h9s/WsPR+zvSr8Lmbd0rxMjLkEMs1zbqwHkcYynu8ab+1/dprOh9PhVrdvJk
wbyhLDbv7uGOe32nthk7PzBTeQaFHxEkoHB0gs3qhYEfL/zuTKPqt6EMj4hCLLz9
b2GSxJf3jkWpmshgW95gBcxOnWbyXdLgR2OlDloeLg45OWeKHfOpQoGETQmYZh8Q
n8Ajm22W+hXoCfr/7u0VDYgrizp29FZWLdnhajkUQNQvDsL4sT6R2haQPzGuUFjM
SLdPddl9Et9gWBxYI35hJYTalQb7tup0duXsgiAF5nrGCVxntF8pX0QgTbQUb4b+
kttXOhVYb1WlTK9YCOB7nlrrrylEcYRevP2/BZMrI4mul35IwMA4VsuuPVrbIOiD
GO+K+7x9q8no8obavReDKBJh+mmmUU0gjahZGUsEXSiVHHlS1Y+p1+Okm3M4y5lw
7RZrqFhX3nGWIbRcuksML37fuMDsym3FVk7aCl6rsFKIeg5yy+wgBllnNQ3Gqvoa
zwTbHP2dpUY0GNoJHXUO/J8Nq+FITfVVS/vJE8LD1/SKFwzdQMfMhFaIaYbU3UtD
znzo5DNni5dsQZ91eWCRfralbF7EhfYnXi/twkZC4f1cmPbF/vZCQKCog4AiiTXw
1aUs5qqiCv4qwBW28YEjqrrapxLL40D+a7bMTRnHO7ABoFvXeuucxntLjVPzlCWt
R9h7cqHRJrgnaEtcwEum0oO0WJh2KdSPWsPgvxfw/O0jzI2JvfzqjRsWtiJVEy4G
p3Y6YnWbtf/bSESLFLKPn8N4BnsricDA3NBhje2uxjJ7M1K7m+ic5jcZNg6VOt4R
8RCgXy4MO6rPvZS+mU31ybsiKzpJhk5h2SvkJuXqTs756gbf7o9gWYWq247SVvpB
5WvmiXKbhUYYRlEKcf8iGY6ha1LSYU+o9Sdgzk8hQygE4nCMkbLQwLqy+83Xm10t
HvlshLm/bZyXqu8elQJHgcacmNigpxX80pUMvcbhpy1pq8gPqaGe4gUv1idl2f+w
jxxBDRWPUKRanxOgWc72HiFQOm0AxrqbLKun53GaVLMCOWDBCfAfTBuw+AbkOC8r
XdA9bhuKi0vBtp+69uIxmjVs6DdiG40oFDVCvhaQJiJGow5xDTNr9rxx28dZ/FeC
jI370rrEeN6TJyZlPB9u9KWylSmQnaQNbdBwYgvTjySJTOz4knxByxl5vIjkaT0d
lVrVaUfgUqQKJfJdkVcucR+/WP36AXKxREgw4xi5ROr/duA3b44d+B7ORp2xgqYh
nLCYaskCL5duZ53Yjf8HpvI8tHb4RfYpsjb8rOlrMAx8TiGHHpInRSuo6e080F8V
WyzvDcCkjn2/hrDpmZqZbZ4+XQMGxA0FUiMrsi+Q3SgBxWFOXvHzEJGixj9IseSh
Ydq9N796rKxLDdGKymoezvVi+nfYX8kounk/O/3mTpotbBF8dnil/BUIcSaetbKq
MLJK4heYTWNIBaYtKx3oW/sDPZ373gPFobVp89hzSmRBgnbXAAnJJLrGqGDEGzlc
LUb+b1WiYUTvUbuQ3ACHRofwziE7v07KpVERw1nU5XdJXMFwKPmCpFkt4/uPA2AL
Fk4WsWxT6dWsAjVPJcCsu4zGrxmdyHe6p+quhldOZhvdSbSnQ0xWkA1KFv9bKed3
95nOAPPeJLxdeDFuvmykmc52q6IByEi22V0USqlmFHUiLFTqDUzvZ+Xwj9ZJIaIF
/1l2rL7Twy4k9b6lNdB8HKcEgd74dCIp5NwvEmjCLe1x5xOsxyExY5KwKhCI2IJg
106gfOuSZUqF/JCnLSh/6DfBtZvLJ7VjEgwT+37ovLIirJFuV/ZL4vXuKK7tRBf9
263jeDxadblITEQ1TDUqpt0kWvBguN3EZlzH6/qoqExbrlhhDDR3Z9XZjGe3iP6s
Q21RGxhaKfpb+hpYAa1xQHp1bjSTOsdpi/Q8wvs6t1yqFdXX8rBdCHJkie3K1aBY
jbwXrqLaJ57F1Mz5raT87hFk/ZKVY11WauKKAyWnme1Re8ggbjhtuS4ts4ZcWj4v
beUqHFmQzFzs4C/coGe5VAOHP01xWMmIWbEh64odajwsBmCQ09bwIhEnxdKIORQk
AzwuW4oRldzfCpIUHOAOi14hdL8ZdqbpA9aVELYCOCrFGBCnAXECSK/x9WSdhsJJ
24bDlEIr7W04EhAlrCHr3MLm2T9mi6JkRoNI0hKD7HRxi1jSi/C6mncD1hVlsnbm
14bJ7mRrErrfWjCkAQHudElfZYQ6PzpNluuHoH4ga4NgFFNI92lqaC1ZWSRMPKDg
NuITl7PdKHcuyVTIjNGzxX/+K/otePBUWW9X6Qv7O7If+INvbH7I6gT2a84SDgGo
TVEUFSdc9ezsiCTCKJ0695bUHlnk0xpDXJuy1dnnKrUlI0gn7VPpok2lZsNYlGT6
oTskecu5ApxZDmiBm8Gx5MvlWBNxB2oft2HdBqiVkEqLHn/50qOmOljV2vXhFZ7u
JDbmD/HszEj93SYTyzAdSkRbYt+VlbodeyZYil9W7sHAIIjOZeGnui8iaqmRC4qT
NerthpsWuQEnEHkGZM7RUihLkZdtaBBOEIUYZ/4JZ3gsnXMn9xmxK2aGxp9qU2OP
IF1F2d81cogdiwm5JS1sON7KnVYy8AWDy1sFvFUZrRIc7NEat+Fs/L1SGnG2s+TM
7ZQx4XNbZOCVpwFSYHeU/5uCPkGt62W9qUCcH7Uim4hKO1aPdzUp16loTuqVeVU/
2aV5hV6ysVix1vg+DgcpNUUZY0+IoPiBgLePQIUtI2EPu5gp3G6u5a2wXAjFqFLP
i+Sr/asVMSRkNrOcjvV8xO8D7vYzW+NEtu9870El0EA/Ce1/xlUsCmPH0sHSRYH3
e/pISstgbW78LW/eQ5v0nZrVMThyjbBt0Np2xCARvVLQKFyfNL+b992L4N5rRzUh
UImuAP1VJ/ryk8sYhK/XJ4JO9ukcK5k7hgQrhDH1or/9/6cMJmY3MjgM36Aq5+Im
Y1xRNlApzVNEz6va5MlV2wyqBJlq91KIoGosU76cOXLnhWaG+8FJf8vZ+2AHDyRl
FSc5C6LWWnNvdrFct0D4XL8SK5U09ZKbWE74dW3w/BkxQwj31vj8Gcs/8jzIBlEA
hshaKeAG9m9MpNr8to25meViNwHXw0EXg+4kFNqcv3q/53F5hiW0vwRmlSdf4RQh
DcAR/RJs6Fg0RBAtS+hz7aXZrBTt2S15Fo34siYASdcLfcTkzsjw6FSjU605lx98
27L6xYKu8D++qWnMLEVZnTiwNWHbbTPwkWRWElPbGZhr8TsqKfjf0ma61qT088RQ
sCQKnUC48bAj+i89spKjNRww2zVh0u78kgmycV/Kee4C8Gmc+o5UJk8zFY9FEOwn
quApYERnjLMxrXI2e19HKJhwUFrgb0O4wRoL/VOtGtDpzH+Yvg4vKUdsdN7JHade
DR+39octJ5eLTfjifWQoL89Lk51Il4qz4DOJ35ENteR5ZMCiyW3QeND3Eod0X5ie
TCPo1Yia2aygyGIQfrCCn0DF6ofjMltTATCrpn8yGUaYcwGPS/urpMMQKykhqe6x
vPvetzaa10/RtZtlEMYdvvY8DvfLYoIanpsrSJ8+d7lBqhqeKtEG7e8Viyq9s8cX
zt5s3QhYTULvATFn1bLGQxv7FRXAbNn6fc56D8mcC1ii5m9ptyHpwBDIkoCJ0rYf
peVjmvoxLmDNAjC7gesSheFuHf6rvtmJePAcwQDq8tbOy0tsZYOH7dMBA+w4X4dF
63kRrw+hfvU5oxCO4Yank2sxVGZ6itjrhdrRGXe2PGzHTLhJCPMYFdbf9WmjW++U
n7AuCtbCvTkjc9J2ca9eZb7LrBE0RNg8sn8LIVXhSyioETUl8DbVHUy5xysZT6Ix
+hmcMfKXDJuHcZFFOcTFwu3FLsA7iuYQz3Rbq2tIUmWD5zgHoo2FDMrmm1dyPdv9
D2I34ppAlJGGocKp4YEihKFttfwJ+khZ/JnmGR/Xcw1IXJnJOWWyAeppoOrmQhiL
81Q4mFBECWSv1I0YAezFZBa4iGBwcmYmlk6ykpiRz1+tu237+7+1ct9f7jhBz63D
0wo403MyUBWNdiFMRpEKfRdJ3M8mWoSQe0uDQ+kjEIsk/MBnJNwuoTpyEnuE6Vau
wedz6qMBG75d2LZUuTLTvNcp2tEVB0ZJacfHkWTViYBR0Qly7Uy6jRIKMN6iilGo
96SOA7PPtm2j1VYaVlH416ky3XvMO16hVeGjVjSJ55nKruUsFDMp7sQZsr/7inPe
mqIRCwtePEI2hIoR0Z7SgrkzkHhWTOFDd1Db5NhB+mzsuF3MNqWkZR2jCWiZFqxq
3ds3w7zWCELcO540UrV2JlKRv7JiECX1a9RJRKIobgB+95HT1/hg9nekNlw/quaP
byhjI6uJmLigMELuiejrckpXfkZ5fwBuWRSTwOxVnuSsILjW30NuqOCUC1pqK3s7
4BID5xli/pdWrxN6u3yCG8VkaIZ3D/VOl+GxtYDCD95yVCeneD2hgzbf/zqn0paT
4MHaae1j9ATOC9FW8UDTfRtJ2Aya2T3loBt8f2l5AHugwI3svmlr6HhZNs0w+b4l
tJUT047EDEtc+COW8j1X5SnYXNe5T3VA27qojQjyNqHk1+wFbiL6p6F5IbkPmV+G
wXmuz6jLXbwv/jJA71xvlOnfMK2qpUrlbPWMZJ4/ucbTb1JFho6hwVaobpCS1K3L
Gb/Fia49YlLHd0Z4H6EpBqZplujNViO+mbyr99+FNCq+GOpbIKPJf1yLAYlFDS36
9oy2LDPAjM71T+7JPwL67yiAaLMb89632oibWtT84S3JuC+Aw76jaDJbmJVcwPmf
C6/prnf9Yvuq8PHNT3oM/RfC/bE/1eqyBLpqrCieHylwnq+wF4Kj72/E0zgCSMxq
kkcAxK9KhPJYY/hd6vx9AwSLPGOC55kiubU1HacpnDXGsR2wLwUwnTIizs3T7Lo2
h+niib1Ek16BmI5K0/QTJLhnIL1sTgKuXstIplYCUqn2JE+A08uJFWHhD0dH0n6B
Z2O0rGdOzkyQ6X0h4MHA3DF99cnwlgJMTy28S2zumczDV3z5kAEywTuNiULke9it
pZ++5aOQhqjOav4GHgkucct9E294RF/p7VQ6Mcr5JuFy4UftMCoXMfWu5xhCzgj6
o6SLonSXQQyFX7/NaEocSahfLyv9t24Q44mZKUvRk0gnEVUhVTjPmjtSH+QSaVHD
te9aylqk61OSU2/B09idlkXeqXxyRr3kkGXFsLSm6r+VYAt6LHcPudJt0L/4ccy8
OY8TM4X3PiKVPgOblHv2+jFBAa8vRK+c5+kzte0mALQ717gsY+t6rDzeAOhIPMNj
+L7TkenTAykZbqOp6zRPSOMGVP7/qTC/h5LWBtu5TDI/WEHpj3/hHwWwPqrFI+7n
P1Y5pQkrEvAS7Pvj8UqyCGKTTDFRXKcQnYph2IjLHf9MAYxLfSTY/+LhHJaMzfpu
N+eeWbWaV3TSvmEdlI5CBpm3B5udkK/0yavfUh0ENM2YVcFFFMNiFNksfYUGxJGg
oh/Vvs5ab46T6lx2britUoFyB+O4KpeRNTGT8Xe00Lo+ARJ7/JJmmTqC5ocUmMhR
MOsAf+PMUEGBcCGo4BX3xtYsnl5qxKIhZS8liUlAujGQdW5pycgXqMLxB/rUN3hz
CsvsNZD93dm6WYMgb2giqdNpoKhPG0wUv9oua82o/cLTiluclfN7xbVQAuU6chJA
Bl7AGbo8KKWQUPiER4b8yP1aHSXWi1p3U4IdvTTa9S3pZM3B78PljJ1i8TLZiVAB
sNG+/IbDGqQQ1HwoFKGNcm1xhexgu41bv8ChvCL4UMkEHColEUaxH7QQ52btcOwW
X6JcMVLK4XRyohlAZ5wQfktONAScUU7w89NjM5cig6bnGXGD58zPqVq2eP8tVUeB
uBG3JozfkwhtkP/2rPcK/42ijvRsTrhzb4PG1f66lo190gqnP/kUrOT2PVC/r4aS
KJII79kUk0xmk9lkUMV8wboxQY6LfHxSCzAzP1T0BrGzOM3gUXacOPQYcCzQ8/MO
YCLg1ejCWuyg0yp3yc5pYRC3g2vvYbudcpg4+1Z9UHlDQ4x0GLjNQvs69urUv6B4
dQW6bRpdJUBDgItH+oDseTDjUyYufD1o+zSwIwLfg8MKdsOWbx6BVRx6eoZh+PEu
XKkqvlA3Jg9HtvElHCikGxvgWBQkK+8LilmZrU6Dx3f39Jyh1IXN75QVp5AbbgSt
F6b0nIHGq5f0vvv+CULR2F577FBKFMLaNCrCJvK9XVVXo4il3zpPPQe9RerR1wWv
ZmAK97D5uvJQ/DPTE+8caDirU3bvjq4KYMvEKHr46I27UwgsQZLzMHeaKKVmjGrL
eamoFn0mxTPsacO2j/If6yWWlbYy4g9YSEr8aDfDGeELEpzCi1s0A2yOnVBIBk8y
6YLm0RKN/WhU6pGbLQMdyYCNWYyT9/0/dBKIZ7Juk67zo16dLZXFdObk7R09oEhI
PYg/dA7cTvorU6A7TdljXtEvFJsUoXQjN69E+GqJz5BVwaNY5cZERVKcfl92q+mg
ikZakHzYH1z5HYDKnxJE/i1qwynrE76AVmsbFw3xAqf7bKfaahVi4EBXTk2ElMo8
McSYlMsOWY9OnSYyU7QVeKvHRn9GdORLNB9Nz6F9dDA3IPpOeX25G90dN507l+uF
9fBMpI+d3nhD4LZFwyW7bvdor/eel9T949bTgSwsSuyScMBJchv70OkJ93/hX0Rp
0xWbD8U6jz38FXKvvnv974voOURXNNaG2Eeid0ox0oiv89F5cc21pqtMpFphCwSs
fuuK0qPvuvfUtFGEXjBny/e+6h74DTbY7M5TPdKhuQuJ8hyxDRuw/SkJTHDZHDNt
6cI2mx63MsoZa7n5CB/gKbm0hBxSr/mmDa4inOPgoZFWCSJ2lcKqtNyHtLLwOgLx
sB4d3a/o5Pq4dy8JQQuTUZQb8AmrEQ8b1z4awYdSplpGPMf8PxFojqCrnmI/Wz5o
sKXYCmMVoFAFPt5enlk6oGwS8aHa/OQwY00/UVlF9c4HaW1zbL/e0r53L9Iqml0h
i17U/pnhf3fn29wZf/+204UY1HQJBVlWh0vassXhvj0naaCMaUrEZuaj1zn5H9sB
7oxGG3AFtg9D1+cN/PkYYcztWIdH+ukk+cvaud9Q0bvm7wHQNsOJKq7k7RjBl0kt
tpqVM7uc+JDUIijcWEWLfbrBWmSrapIscOxUnmdhq1UYpXr7WXr7xoAYhTHlFzR9
Xa0WFS+f75vD7qWdpZcxKYHRnUPzT6ho26pRXkAK3sJO5BI2IW4k3i15HWWu30qC
BFtVscZrEketbJmgVY+hRNR0vrQxie0qL070HX1XfbArfQ66L2boHB9Ul9cdFn6P
sTw8FWXlsFsGLQjySJd6PJJ716CYU0A2nINAZiS8IzqurjepUFRN3jAHH4CXZrmc
UPsTZIrKCf2TcJgwZ6V6IkItWV3OPSOCjWeP0ImoKJ3qI8g57fV1Hnu4mwpFZGIq
rIRiSiuxL79khYASk7zrPBhIfq9devCQjBRJ1bK344qeQnRumYkoggWCH6EFtz5X
XH0P8//FyeBRvuhKYH6EotUSGrs/WMCDBFASHp5b2oPO1OEE//VypNeIPvxUS8zY
Q/rmaY1oUHRkM7O+T9VmPZi1l6chAx7CtXNZMP7N+jAh6kTD8JmOE47hovzMMPlB
sGCJtFU8CrRQO67W83N3GcNB/W1Pam2ay7SHLDOmodatzo70mmd7w/3oiUxi+NaS
hIUTo5ODeZ3+dKF86588mSGk969KTyUQVdUVNmmiZ3MRU1j6t86Oejq2ZRQzTZIz
AregjcDe+y80sp0KL1ASpuy0QOO5j2zh+0b7OoChLafUKHGQMRoDf/1OvllsesI7
VMH48YkmGalQI1DKRXWIK1tmmySWnErK0vLHx8Y9zlXVwvrPYQbpOk/tHS7t6gw3
1DaRbSINV5++n8Fx6GCz6IHgia4+uSt9d7wJeXbq+gh36tEa+OlUXt0Ia8zHbmQN
HC4IMBEcSvoj504jNtzbfJ+POVIIICvBx2m62frEuYCIjMX9j6M7LdcxcwTERaEP
IX/EHvZZpMDGeVo36mTLoxM1GYyG4no3whJjykThJHEXghecG0ocVpazlcLSvNOJ
EhUk01iu5ZQP0WwweEUHQj4nm++ELvIQk4PfVhDyFgsTBEQoripsGH/bRDeTsX0O
wvmCiqRRRU5M8TQKduBkmBNj/Y7m5Wvesh/cVDkl77WpxTW/QFpslV5hF5ttdQDP
tJEzVkmrG558SX9rsEMOvAf+NDst7oFpJrZq1HhdqnJBA59ilhgvCw7CH8thjhEZ
DefF18iAwrtxonHmTWOQFnA5phzafI13mSBQvccUOof2Duhqf9HovLNoYK3B8Kxu
UHsCso4JLZ+fpjSRbcz3Miwb0agpjUVqFRDhHTVr1uXZ9WhNvDVzbCE0iPrsAd/9
LojLJoVqPa+GjJf39mHv/UG5cvBLIgBnRmZ8JIAAqP6gS02/tayiuyZYK3db9KHx
gyRgys21QI+GlyHJ9xpx8pl6JtQ0Yx/mxJ47gs/V2fd6RJcUnjIshKv/Z/7vMVt4
m95GjEFnkd9wzdmEyOlo3YS7qPMGYhCoP5s7RkFBnEQtQgW7rorgHHiQxPdhoY4m
ZG4/SRPUaHBfZwBTmo6QBvtQNA2So5Rdizox5AEabc2wEQ0kaDcVMIY56ZU7Vjdw
/6Ae7QqCAVqXIZOg9N6taR9/mfJFzJCdGXaJ1uLbB8U6lte6j3Dymr/chI/IMfUM
MGnGD/SB2+kBVBejWqnywo5tlnF75b1CtACFKY4ckPpNpmkoT2MWYpXDVTsP/HJT
vESBkW6ISaNhYouLsgPzF7tli7AYrMnDSXjqXI2at4Pzp+HeF7cE8vgdsuuAnTes
ON+yhuJDsunYhtYSmB/AqyC4tNgaWlUR+jDIlNcHM0x+webrYTu1vgV1dNZ6zq7B
6X/U5lemIbI+ecZRTnhDsUwZoyOuN3OpLs4X/Qc67xXdAugXJ0qPZbG8YX/Sa7HZ
V7MQBOlstizIjpVdjkiJh3KzU5PPhhFdno9IKcbl4wRSAav7enliCPI2SNOM9ThP
QdXigdlLRxqrwZq1khBuU9CzYLY5rS5jaL9dNXUpqk4T9oW3qP35+9Np8CCBRHAD
9SVbPEvmMqOIlDntct8IBP0hJQ9RmY5iKBO5/pWAGelg1UqhHITkfPHEAaPisZQn
ALa/9w0FuatEsRziRoEdDzAjdwfO2QTndW87UMTcaHJMyM9+IWS5X3pW1rrlFm7W
qX7wOF0jQF8SSPv9nOuBlKmFB7g5I5lrCIgpSrvLN44FMxlmPmcP3yYlocL1g6d9
2M1gjAITJ+2KqD8ne9KW51H/TXYiG2OFE886Yumf8jEB0yyjVTjB+BHNysM/DsFp
DnB3LMjaXK0jLzuKnrHbZZeDnft6zMikCosCk3L/ewYbQbdXyFXLTVymujjkTMRM
81c+UAncAfzFYEdIF9KlVKxOLiVhllQuZz0dfUF51NxdzjkqXQ9sB95aZW5W8rCw
hhZnWlpktIGguU2HFMkzmhtIkm/chwGMlfy8ThtRzBbWM/LgHYNWzxRrGvpk4D05
Kck3tLNZ9bt/ZjJl19tzWvZZySx8wvKC2jBo3JmQswmZkB0anCPZSPLEQ2lEb1Zg
HODuIpb5x3mgpGJKBw/kVakwaUOB0Rri2yFW8EoWQqKdES3EHCqCr1luVCcIO1tb
CTdnnvCYJgmihlEi7BgtINE/5C/84XTLgRcz576NDvp/Mvcs7haO8G8vXiYkHvlm
p6FAzH4l+q2XNGKh+itSX2VhT/xH+FAFMxw2sknJtQVx1q83TUZw9koUyK7mD6WB
9gFgU6uRnJOde4qGNa86hI1OSa+df22HTuG276y9Lws2zwm4QoRuUIv8L/3TH3YN
Vgks1DSnAx/UHvypEQAA8vtOHdvaQ3cgcDZNHBuj7Kb5i5VTvC4YcAdS023obYSP
09T+7sKzNghkt2h0gBC8Ysaf8b084sZZ+nnrnpPXRwv3rfueAFUeuwtR0quGWNs5
akUTPXD4mxuEv4VIo1kWbmR0g8Ti2Zvjpq1PgP/ScthuJ59N9noMHGqmBXAs/vwx
SVEmwhVGH5lJQGqTgffqEJhRot9siumnwmNc1Oc9mttk80fgay8jejeaQfod0Lpy
aPlZcniYbbrxYREz+aH7iDq+SAiCnN01VXCk8HVPUtvw/QSmP/KTcfBI9WSWO0JV
3vEHGjIufxwh75pKj32UzzXu4MQXDy7d5CBHJB1ZtE0OjCFiNOIG1lXqI7wvYVHk
CqmYHG5nkXSuM0weceXfRN1+amW79Wa57v662t8dAB3ogObaWe3bXIuLeXOOmD+A
FvPoiK64drOacww+nQK58I7fu45kUuw2+X58W5D5zJWWwNLCgNl5PsU5KgiW/Tcx
7fVkgiBLnQdoLfv1fS2heIMEzZQwZNJ80XbTtlL0QKcks25J2RSmzLs8nU+nESQB
fwTpbQWDSJUXjaR0jNO/3ZNYr3kNQz9BscfeFj01/IpV3WczX+Ys8xY7vuBiF8Af
hqWcMlm+jLyQ2HQipPwgwAuTY1CUz7QTYMYtJi0W5wC7R+kga+VmzczI3X1Po6us
ywcLJRZk4cZWAC8W+HQW6Wc3CnEMIc509gSvEy7vIyGkMe8S+t5UocoLH+a6vWwX
soLgWNGtYIcbhZkcsTDQMiEdLgafFAZxluaElxA2jMOkA6ZTyfMQ9pzEd8XLjLJi
q9bZflBg3YjrBvwAdU5+NXxJgzVkfJcILwI/RRiyww8cuYeV/xrwlfFSD8mg0YJl
VphcQNZFUqWDKBt+BhsVPPyAMFaBiUKWBG/FPwXyuANWF+MkGLz8MsmG8jLZsZmy
WOE3TrtQGFHGdMH7+xwNc8kzvNutfBIpV6gB8XksRV8z4CBfabRWlfA+3yt/725S
RxbUx1O/piTiN9+0UAcyMATE5zq78EeZiGygJ6EuVnLK5zPluVr+2x1S2aBfJdR2
KL5OaVnEJZ+mL3cTNbe8Pw5h9b97rtRuISIti7lrWKJz1JfN1h/917+LWfH8WKsu
WNWSQsgm2KdorIAEh8WDI1sx4PxydOjLQC9vwLXJv3/OYvZxjdS+qTRnrksSuOiI
njRnJ1+H2jDhuhwr//mZkKtBDkSL4ur075jWzQS4YPv5ymoMYPQGGXVf0kOD5IYl
xl4xUJqK3TwkPOoatzMWtWSxxfTPyIB32xmzG+Xr6RTzcnz4xL9H+GsI6VWZBaUj
p8KLIEW83aBi78K1zKzdROXYRJ0kS0F95OVJYAeBoMpCMDzsXdxCPkMms7lKjLJI
+ms72uzosQ/7b9+Cv1rq395mWJDPtHEoau9uYwBS3jCUmcKuP8FHElumkHg3qzur
DaBSD2GuWVzNOVdPXY1/vjIBYtlRFOp3AXFOUO3TpHY9cdVOxGZi32TpgbyTSsuO
ZmggqPGbGDKYFhZ50M5te9Fatd05DASnVOfwC0C7Q+KwSH4t4qdwFiV9ScKNanyR
SyO1J0zaoxzKHma/ntAZ7Dxi9R2+owzYu7aUmv7d54hOjXYYgUoXgISsgJ4/zEjk
iKk7Quq4UWPKKuKWLE5oL/3gZcxPFoOZM8qY+uRW5Avt4shA0o8kmTtqZR3p83cK
o21EFCOR6eKiGEYC3TCQKhmwsimiskTCrWMcDdVS+IJbRlF5TYjV1YJaaT99bB1E
jeNk2zr1NCRBWFAccpUn5cuWbQJzXBeLnl0vH2lk/ronwWKdqaXU2f7DxABSNHtp
1bXO3r8jlqlODmYtppUI4Ftn5jNPkot416tkCZ3qdCaHMAiSyYCap8Q8MzG6h+Rh
hhb8PuAskcPsORrz4lmuB+0QbdNtdUMhWZvwWH/DwjAU4eZgphhiwD1SGsO+dAVD
CjIPJ6HZJ+kVygRCh9+WUP5Wwg22hnvzts0lJ6IAI6SYm2w0d9PQu4QGsz4YSkj8
e+ifUGdDDX8S4c3u1CqVquvgPmJrPMMn+B1aaR1AFjVbeZyVC+fW/MnxNeM4nH3P
Rz1aV8nH9hoTAw8hX7KeXy3ho6USKx3Fo16h6qdyKdxHVA0b2HxvaRAokuueyxHv
QJWv1VQaDI4OYsCXUEu3i3hBjWDpFeyKqM4nJvR07WLcKbFewEWIVNW098bEIcGg
oIwRFy1V//FGnsnNpllxsWXPi/jtGis30E2fXdibc4Fe355mCxEjz4S38NArw9dX
SoIX37htF/gU8PdgE7RaJkQRqjf/pR/PKqc1rmACPfqu/c9dq7ljJxYevmdYOxOo
xwIGbivkBXSgMAkwaKL1JXoDG0yKiQhiH7PP7CheHxbQ8FRCLMzwzoc0zEZcEAww
qEPJo778cVMIijs8IYiYDiEM5LD+KD1Uk6ZWN5H7defgNA8vB67DBtrLw4WBNWSA
oo4JhAB4uFKucuu+RajDhrM7LY6BJDu22YWUyicxLz7WpTwLBXLDRZolW7PQ5Nwr
sn6DAdaaFaLQHNM3RgYnDW3wv1LyJ27PXos3tfXIg9z0zH1xXFs/2c616Q6u614h
KlYlaUt5ni4xsy/6wvcerSyJg+/9KFLgEBD+5qe82Ql19ylO7kPvGFzxI/xFbYQ+
lkOM0H0+bZ+tPfgTAlG6gVLsh5jdMWeHkXGC7yWEcYJHGL9HZJrxkGP9pttb8mH1
AiSe6r0LrjTf35QO+rzP1kThU3K5mq2o9HN2UOWlai27LBQ9O0oqkxQJh3wR/JhF
4vp+wm7OBpH0+Ei06iMklIxTe5202iYztIFugQOFPxH0LifZEaLxNYYWyGuC/8yq
TBGgby56enANWRkRi78ZXydzZYf0xEwtT+sLh8pcLxSHYtoF1CBleeUP4f17SFuA
FWDOwb2TE8CeqdaT8l49yyPgkQ6QypDkmwxuj8HuYqo826ZLZneIv7YtqsLgbeeS
nS4D3CkQRxs+QnkQOmims2r7iAXuzmFkQYeRrMnOlfBhgqxEe58Vz7qPilqN2075
YYOZ1Ox2VvQlzdyM+W3/26qm4YTxX7NSmb//cdNJmMTxVhLU8eJX0eEGaNTGhS3U
9W8jKnpoF6UixFK/QobXXY3ADXFj/aWk6A/k/7cLUzTLxQ5g1iF7Zs7rH6+xMjF+
/vEAOjWDDgIuXjwlWtnsbUXdPnwdnIVexoC+Mu7zaXDhF//1Zm8ZTvEtzDZ2uvL0
S7jATdAGscPfpOYOgksNSj26Yl9eqSuNaleTaaT5H6FNktp6XlylhDW7LSTC5WOH
fR5g0YktxWkFndehsVgAT8NY6iDKnAFxEAo9WpK3oGZ/yLEpaZ1iLHmFqzvUxz8P
AyvZ/tOnK1rRgwl26jVRea7N0n3Er8mrYSO0Q5KY+VQpLB9CrxGLJZg+aQQW32zr
3V098TUvE0cd+CiATNr/Air1m95jEjOiDtTfj3ohQ4L1JsY/Obz5KMtYy56YF88b
z0ts+cWhb4aK2GBnJNqPLqTI67guZWB8MNcfb+Kc3medN5Lg9ob8ZNO/zbt/Vua9
D2Df7XpszoVeUdtfoebLRQ+omDRcVwR9hmGfYW6kPTo49mNl4t0IK6n8Z4/FqIqR
9lgItCc6mEP71XDGUYa+EuFOv29LIXzEBmK7kpdnfF8h4BQfM4oXuTiH3NRCrHea
SlWZCoiX4hspcO6rPC/iIpspluScvTdOyHBtKwkntJYEd4u+SRg0nG40yFNMCiRt
9+17jSAMxTgTD1XR/zSPlqavdTCFgbv5qSqK8OcNgNaPn3J7qSAG7yftfU/zxMaH
6ZQQ3ZeHXZJbG9bv0wHZu86q0RM/SgZ+PlbdCL5koj4OXpyNDWCJW6xqNdO8MPfs
fxyrMLlMOJILEHc+xMcDclMkardaX4xnmeuURXCzhQp6zcARVlqnDX/rTIcHNLmj
n/X89kvZbKcDOgMzGpcRn4mz5b9K9dlLIsJz82Wnyy2rnmFvKjzxNv1uIseDBand
sXeZqi/mxlh9nW/70CFtt/L5uxCjd0KkGuYQowfI6Fiuu6vNz6vvBKnpmStadin1
rSo4PZg1q99GYLV8l5eOJsIQX3h9mv275ZrKXASmjrdZhjJAivHCWc7Sc6egdl5k
qWLCY1208vdi8IRyHjkHbsVMn14+ok2PBpB4l86jkypHrHEzcBQzGLB9oDNC4oSj
YTZbH9jNBRXsWuhc8k7DeiBfRiz4d6grJZfAN7HDfuKQd+1DH5xSraDi8OTkdb8U
qp2XXSdSMlEPPmywaGjHAvpVD4FvFfdqdTJooicjBM3soVV4sRu0FbK/fEeVY3Tt
YCbDQyUFxx7kmWTZbskJAVDPDGtiaczOUHYjBSnoWzl4fOfMgwMV5Drvzf7nvH2G
9Ga2IUSAaQ/emM7lTinXY/ANtJ6Ki2IQAnRzytca+9xN+nKBoeCNcF5lBgowaI6l
i9MReog4NCQdZ8myqDy+3e9j6McRzRjpGuwt28/Rj7DvgqzkzPnhkcHR2ciGOK9J
7LQRt1QeQHSxm3duizzKV45lVEOfXFRSkUPP2Ir8Ngb2yEBkgtEkdbi7K+v30+4/
IQsNfnEbW3/KNNeJgjJRD7gj6yo/TkBrG1tBrOcsH/vT5Tp3ZTN3qPiHeUuOcx1b
aCDgDIDwvs5J+8ZcBO3Cf2wiXB4sT+iL2s8h1If958j/z27XGOb99jS6bfa6avAd
UbSY+dJYm9abEmL8QZ89txPdQLOu++Y6MM50Am7h65O0ov5HCZYhoMdRlTzjieNY
K00pbqiDpKaIewvJBB669HeOFE+oi2mV8GgoJRp55+AEOThptZpTHXItpC6VyuSB
t2FaGnglF4O5gG9KvJPlouyduNHuRI/0LQFWmuaIVKXH3xGIexlZbzQvpWDFhwgZ
SeeLsxWAxh7fi95b4dFnlsLj3dg52nxisnMIkZAeESYiZETcTleqOuPv9UmZXqCc
jlEBqnimYRjZLEFs2vHmIMzKVnTLRXivh+hXBVRcnkkt+hyPnzxG0jJbgfiXBPmd
Ei5OxbrgNQbG2sHwc+QuW88Ove/U4Vhb2FY7Ql4gBOJTwtNZ2xAsAtAVwo2lPcW3
VTcA/9U0GgqxX9LRCusI89wu+CCbYGSY9SzVKEmeQ7YeNRhWpuMuIFoxGAqPgQ0g
hvr8lcv2Tbv68+31S969F/Awst3WG2mra5VbA+OtTRhmNWkZ7MAmbY662cm/J4sL
i0UWqgAf5JkzToQvAkbx3GjcrxWfhcdG2aSrfqXEzDL7aESqXRpFWS1b50OtnDg+
661vJ2id0+guT2Ggas4Z4Cn2HZP94Jm6h/SgbLiiedipF7mOii94/rdv1c4PaIDj
hyRxqgqWIVXA9UGpw+sH7eQpRns/COFo60cL31l6qJwyrZaABzwgOMs4dkFi7rf1
Lu1AQyGoqyBpj2HaJVrfvq/vSA5Tlariy78OQtX9eCzy8g4JsIZY+osUAcRd44Lp
ic7QvLH03LJccwVh/o9/4VsYgtI+7Y34+INRUOFBOzzpT60ktOf9E9RWRuDnMq6Y
ODAtBs9b+LIdxVfaZqJ1LGeUc9D+UDeyqN3TCTdaoevUXMVUHbSiw5SfPKbHECDR
mzDZwdMl0+uTYdMh5kZQsbsLojzxECPycSh+S5PGyI+L8Ac30bYmu0Z5EMYqqRTe
TXOPNiH3hX2LnjosieySGcvFPfWa4xXPDsMr7Zfl76DN8Ew8dhtVNuJvDed+M6iN
LIfRCFCOMhslm++jFCMBylStYWULPf1/7SrlesSfzFY90WqZOca25If3uyjkVSXc
F4M2lGEKqtkT+dd1obJJi3YEcpeW6gigNtWP7W3MBylAnD03aJlXi8Yvi68QDYza
SbTRyhOdweRIqxIls2G2LRuEIhXDjoOVaMxHKULH4UqUWsQSURjdScR8nUDgLkD1
m51VXbLEdG1bPNcTo1PymNml1sTv0TJ0yccSj/rrMWsI6yr9SuXQap3AVjMnAO5z
LMNvMePB3N6YmEaRgDjk1w4mHawslkTRYcCTHTU0rrzTtg3jDVUcEwhawfG00Vox
riu/gm4WYKl9n7nIuneUh3ctVfpsliQJHgVge7MRp92co/grlWoDDhFNqJD6zZhV
GcUXKMhgTasSICwCm2AI45rnrdf+mwmtoUuT976PfNSx/qOtIUhIa30+ctAdor2E
n0iR+oBhtOPKHLTUdYDhl0hBt+Oii5pA/YdQWroXHILDMwiyJYnNXsUbP2WY1j0H
Izvj1q9Sa15ytlBJHtkP5UYqHbXdXnmBY1veX1A9r3pTZrlL0b9WIvNSFIqXkLbm
YGeN9AXG8MiFatni1SWgapiQl6yMpyc59rnXqRjmlgTV1NeLa6sHha7nAzI8oHOF
Eqr0hzLQa/DEwrCB8yVDxvSYpON0Tb6b+p5qiNBa3cm7LCc5crJX5x2QbdQKwhq5
f5jEPaY1woF6X4zXSSFcbzBhbbfU4XEOovD2Erl4Q1pwdr4tbX0/gILBeJrgmSYR
O5CMDSRKNdpI5Qv4+9B6hyZIHF7WMD8nSPLlmECNxqlsYodhj68ReJKsJJStT2AF
XNM4pYOjnsGxFkbC4G01ilMXMizgK8ALp+qX8CEW3T6Ms12dq8ZelgoUEF/Ll0lO
0yy2NZxTWixYLKHencR842yzdDIGmxDEkdKW86v4Nw8Sc7Po8TzZ2hHoT6QA9f3h
L3pI5C3u4vejP4Q/CzKXyFeaPghUXFSGxDtkFe0CfeLrEd6VXfftW8GB5NaVs82K
mbT8IJG1Z/DKkZu9ZKSxaIMDP11CPhUu0w9676XqiXobjbG7IneBLzg6kNklEYZ7
C18LL5Chs39Qhv9N4oEuYm7YDTmL2god3sI3yGEM5/jvcyUHHIcRHSN/pPOUZCZO
GiSkV7mw0xqPGMgk2q6h7uhl7wItzGS+dsPqvXiBNKctvPGkDJnBurOspgdaBU16
zthvM05w6sKd63mhhe44xtBdz0yAfLClmAvvqkcFiJT3AKVcEjeSZDGaBHF0ZMA2
zLsuOvbktZ+leM9/N04jn1QeNCRHbRBsEBtFqYzJHyLoMKxWELsvAlGeYde3WcSc
L3/zo6zWYFUe+NLCGQbEVWarD7iQVRlnuyIyigTAXEE9IUezr8H4XYTupzwrqsbE
lx+v9s9qqO7XoQCyqiXXC1VLE9kVFQyyXeohZ08qkExp1TQhMfSawk6mnVPBZlXB
u5ytswAJOlPC8IXzPStWgdEmRbjowkuzavwQgZ4JIxo34s8U4GlVAe+fwTOxqkwd
Tcob6vSwd8NMzdGL744jgQuDSF+5KgeBCl2bSg7/eYmgAZ59xcvAboB2HZzQQ4S9
/Pf3rr87DujW8JUXAmqTyKf/6TGz2hwlHesJDW+suuSb+YaHCxWkJ6bjvrWCFfv0
50dt+ntZyTbxItF6JEfJGTwLrLgiTN7tTOFlxVHCKN1KQdThnZ33AG/bb7aGpqDw
d4v3sz6X7kH7yokoxH4KmTOD0FMLKwBxZcvqGBd5wK80Fewp8aaUJ+d4GLssXT1q
WyIwbnbZHD47H8Zk4t/snEFaVTUFtSdLMzetbOBFsSHIbxipetWM2dNrSe94C9u8
BNkyB3QEzQdfqoklIYr6clyqhIDNN7PWb+1mDzSpuV9X53X4aAXZnwAMoHEAGCmU
32Lnzxhuye3TILTjPmotTe5uH1P8tCygQbILiTUXkuwh9+mbhBnBZbA3/ZNq7YdV
3XGa77/a2EwlQezJHrwsYGAFTtl4/dI4xnOs7PSk7OKH5RaLguJcV1Ea7ghq5R5k
pa1aXtUT/NcmOGzFyF9QN704k0U227sm+mCLLraBep9Y6UbQs0AysCD/4f8BnFUw
cXqs7xJ4fMzJM5qGl7+51dRMANaaPm6zOINXNOMSeadouSh18LuqhTrEo1N07dCH
WDz6mTuGAGDLu7OyUgjRjxm+nS5l72CtRTuk6RMNF6q95+S2Hq6Hk7PDfih+lexR
yV68/4V+8hzkae7PypD6nf2LaUndZzfaRSU4aaVNt/FFW7lhwdBedq5SXEqzx4PD
nmPOhWOoE6p6HVdfP9ihdfFkZhfAN3fyU6CiOc0hxHfQYV191/ZUM0WVi8LMh5CU
Cu+r375PzqYuRBmU6nwQ8SZ1F3TwrKZO5Pk+Mie7JOuV6Dm0+8nuKLyQx7aebxlv
EIuoT+JLPE8vHenqV/xxwUHI9aUvgarq1fAPXF7PiC2MBvZpwOJma7JLRpKku2hG
v764sr70X2cG6cQpKv6UOziFynR/KxZR3iyvNYgszVxw4s4dLX34hWQuETNYkb2x
90ENZ5t7RJp2tBSo6wM7HRLWy2SS4+BCXC8z2b0LmbIiNTauqq73DMZiuf4US8e5
6P1yKIeKVmmBkS1sGmGfqNL3I1OsUN76DBqjb5pJLdflJx26fmVe1N2JLu7fvsV1
JutWuH8CiB4eJ3FNQo7ABojjQXw/3mp9On+8nYTleKDzEy6tOJLyGU7eXDMfS/wG
zy1jJ+LYQo8cn9K4JP7iGotd9MTlX5WKT8E2S17/cV+TKq5mi4fQaZGHWOXg0Dc0
oRrZ4wWj0jZyEx7FoWQpd7/ftco6P1xT1gXsLf+6kzVAbrGAP/USlccIaPz58Obv
qdk7pq4t0XaFrp73E9giq5Dmjfbjpr6fv9+ybRqiiBBf+uHhTZ4M9S7zoyWSLOZ7
Rhvnlv/WsXn7XFy9ZePxgCRKez1s9B9EjltnJb/qMOcVPvuKCcTYk7x1lZd6apVn
wrrUcJMnvGXVNjxYnluxuZUaCZ8rCGNHuh6HgfmrUhbBtWyF+Vr44KHNK+rET613
4xPfYUYD8qENeHyFaftGfNOKEa0WO/DaIiXLQeW/QUEQGCzN3RaqlbVGb1DVWWll
+hTceO4SNeTDotGbCZA3QOHb092+2MiCERZS3jd5h90GTADpd2njT40kWjoGyeUS
RsHVKD/2pCKUPoh1/q0QA2GuTTHILcIP+uhhFDGPPRR7VFWptfap8eNP6WFA+4rY
Avpf8TMUi1+bU3+w51XQieGJbPhPMT4GhiFBz1peU+UPddlX9eyesuHnygUzIpfc
DKPNbqfZjhVNci0uH3GoFXZ1DXvo3ToMbpGcL1dM+s4ybaiQh/ux1E7dZ1dBdPgz
/+WpvAzw3UP9jLDiyp2XCoROTSP4vjAvI8dyGTM+wdQHyr9LvGtVJ0g5HkkDk6mL
/4uhPwpGwGiokmhPK6TxnqJZbxTTfpxikjJBH5SzYCU8XpX3iQKEEeky2FyXVRoW
FYYdxZ/OxIyfgGXZfitAgQqZI9MoBtQa0NC9T5plpL8RqMbP9YPhRZoIMdycyNjB
JSvvuibvsMPxi3Q32QgxAlL5NOcZnG3vevWnLJNYhV7VRujrSqnZ+fSvVydJg0Bu
ESse5gmZBmnQgwDBioeW0llxumwJ7D9sKLp9K+R2XRjI7HervRjWgjG59woMArVh
1MlM1sgnJoP2USFVTuQd5h3aQEuUV7cbqtnmf5NaxpVrCd/Xgdj4+HKDkFAJpkRY
3Q0GjDev9BGPrHp6ws7X0oy4+bvoaeFupCbXZr3uF0Nf/H5wDVpsIq3T9yWlMc8K
wbUqKTHaxIKiY/6gwynsQET6vcPbK41nONDMghnthHRGy0Kc1Um34QJAYTM+eNZG
/oNQuyHhqfjHoaI2WXK1k1SABDTJWffH+gt99gOP/p+dme88GnRwkj6HfQD6+qOa
I5+8vguNMgfOaCW+652CD5qZV3ZTDX03Q9zZF6P/b4K2oWw8fvq+Aub2v5Y94lVc
G8Em/F2ibSjwH4fBbpQoN2bpaZ69bD+tge4xOoSMqssHsmMPiR0OTIaOKFI5/DTD
/i6ts4BFeAotFY0qs+tPKDly5bs56SmbVES0PL1w+/4Qj2qLrNm/fFIAYrW/LdNJ
CeXDx/G3qW6DthAiN7SWKy6lq93dW6pTQCpPonp98v8EYS/lVgwR1J9NunJlY+Zu
Etd6waflXJb9wwZBYkbTFNavq+ivu/lMhpkKveMUen/WjHLya1NiFlFRX4c8PzvG
ronDRAw7Jk8dpi9/Qva+ytgqlb/SSVtUm2dX/EO/kx+z68XkaKvOYDGTubyVDngo
cw4mSJiF+WIsB22jgMaFnfgHffQHZ5dlCZ7/c2VNbGsWP4CmSD2PDHQls4jy0b/g
ocdN9DXiTsTUWorQrw7cVR0Ar7XV+whtq4jAkgSPSiTFfVFntcz5uifcTdEWiS2+
YoGgTaPOmJEQ1I9gz0qgsGBLZVF+3wPraYq4b4JNOlp7LremwgM+q4g7HxZc8aqz
c+UxxJwInOL52sDo7WtaEz/sPUgVpgtv7X2kiuhghyCCHK2ktsFn8Z4nWd2kggU8
188hgpahnQy7ea0vr23phWH4jDv050e6JMeMZbSwzBWzZnTlGElGE1Q7R1DPM0W6
EvP7HUoPgYyUC7m/gUrTYUyd2DXpIh/dVaLOHT2Wd8ZJNvDxl5n/jvP8cpaSBPl7
YhcSo5xAI33WlPN40lhCBGcGD62T94inAy3Xq/cewbf6bgOuZqtVfk8bZb7DzhOa
cHuptoXdBeubENvGq0NT3+FeZmz1riqkhLrIpdrI1drapgaaqbo5XazRYraILPe+
IHbVYR4QG9CeSDdrnCRcmEu4odtgQ8XjPupn6/iRXRVblLKZ0psNMjw8IvAp9Mvu
X+Jf+0ANN/tfAiDc5UHfK8XqGoMEplNYpy3jSpHqFe5GClHTd4ianKgCRjpq3AAk
QhJtYiV4zCMhN7T74segxD0p85yk6nMpq2QnY106owBp8nFYd9hbxg4IcSd7hf8G
wmlBXNXB9NG7YeON6Nw8kkKLZv3Zdmu2N4LxG4huT4uFs67C+xBCTq1SBh3CLiBV
wDP5U0WglG4nG9/Cq4tc75IwffHtHXrh6p8z9YeL3XkfMWG0W2yVhjlCrC3DCSqX
xx1+sDGwXHb9jhFJVEsqIjGCWXXYFYtZTTKhBTWIvEtO7FCmPW3eO95z054aJ1w6
/KfA/KLo6q+Vft8dVKQNSTlbDwX1mZC+hZpE2P36EPaM7/DDrzhd2QegtEftha9L
cOusuFjXYRVg06gzTa3Mk2Gn+IVfL/xlyIwYbFcQJvyKs3ANsv9cR7+epjksKV+1
ZGknsSdaFuC7BJyMspUb5UBz/65D8sA4N7AVEatJytafUjAICXLPQaJG4pFqFSCD
Rzhx8mHkn6MKWMXLmhKeTc2Qh4325ywPmG7R7Z8vdvas5nI+Hxic78ABQo6MnTNi
u1wgxYazrGMsoOm0vSa8KoGCShPxPEh1DdxR7H9H8wSLYnAQYoil9JgYfJNg1gU+
JI3ZA+n9Oqs1wGkx9ehtw8jmwXBsNqRqzNS+mGJBNIqutWn63hDHXldcAvHhrgDR
tBwKH66CfmwUQuylfYmxDWI+GUum0fEgH7CE0AVErjYYg8ZsRJPJX+kMf00JBBjL
Tvy2fdayEXvum/VLVHalcXIJNWfFh9tGjgWze50AUVUD9OS8XioczZaqzAwEm/ey
nFIqiWayjWWKvQNxjm/nzgdaELBdU4yNHKPQwitFZ+yinSJNynQ0hrBAkHf1xik6
NrBfgVqQdpMv52DVIKyK8EfaplIEJtWhorQ6Qrn7P8c54eEHc7Xcrejd2Q760gw8
pDk7H7WKRfURNu+ASO499MWjD6HkIwhzokzpZz9nefsxxyE189HYvE4DylNRWZPy
RUXsjSRbm2R1Edi+2bAbECJRj7udLZpCmVXv590655At+1hkt1DFxPB7ltSviFtk
hruk/nIxHJIrNY1uSaZIqcoVojiaSVk5Fv4V18b7G1l9A/UpH18HFRdGMmgt1h56
7IBGtJMDvlTLX+5yBgeXQnrTOEbAMo7gHKxfj6EGbLV46FhAGOpBaxO26raf9DJV
mdqeor8M7/W+9A2LXi37MCjRahOEiT7R067hUYGMOPHahWlNAzSX7hg6431peh0a
QSrEOtkgAEEiPIRAp0flgdybUdbDrE/uYpjGCzeamXB8R3z2s/pfkDVIU0rV2y8T
XHKWVi94mIvQUnVAl4mOmKPmfZfudR8CDui8sHXcdQCVpV9e89c/n84/CBm8NDQU
Bgmh2kSBl/TonugbuvtDl3PdiONCkWI6UkpYAYDFV23cGL0TCBYM2kU2hN5NS5EI
wtHnVL2nBCzA3lvEj4Qz0r6L2pFzrmd5QAo0aAKgRXM08zsNVsGPTJ6GeHVlfS4C
sH+89kl+YxcgWGe38gI3ty0vKm+/vD6oJ/Hdpz6bPqrElnCvMCLUXLSxG/Dib7g8
8esvqrD637sacYRanevz4mKf80xew1+OkCp7LP6p7veBPmBMHS7gJD0aJAOxhshX
xb84a0RARxB8M3fSimOgfYCeS276sQqDPVprs5cDEedJs1MfHYw5HB5moe4mE+XY
obxHWnjTm16LJYDVnRZSxgmbLsCB6ZwRUBAqwq4N2RlWbAUPxyc/V7izy5giH8RY
BEWXw7tx8OR0ZjxtBiQb19ms69ipoPLsXOEIs1PXciPArXVabNyuhdTPgGuelSmk
qGhnbfoM0o4MWWMtVPqGuY8Q8L+rmg96bPDDIsVrTMnPirSt1BTS/fvJQYkLr3R6
Js3pMDsP9ugOep/DSKS5Q4NCpuCbaPtL9b+qZYwgmwHCbNwUKnbMnoSE4FgB+TwV
EJKet7fIZ2NyLgXidvk9YDt0z47a7t0M+7hlt4/VVJLTEnHoMAN4nB/zIhv+ccRo
WRPwUfc69P94TuvN6C8ZIPemr04wkR5jOL6U43uuc4CVW0SxB0N+ETCRXbrhmPYp
avD73sG31vA2hPfCyR5uTngD8jd9WeeMLAKHCCoRKq2LrgvTKJXVDhcXplMWWJYj
H8Zyzc9is3KLqqoU0WeafkcYZ0DJ7chrl6hVPjkgQierduUiE8XA1pzIba8V9sSb
ed+M7KjexIA6wgYgNqd0fsdEXrJskZs1NHR7yypp7QIJ6CWoiy+TvQaSKqVmBZ4a
oxBkzmUVrBXateMtUbjv1NN1jCdQWZ3mPo7L0DeHx8g6sewKSiBVBa7L1y2w0w8j
lpcFKrRl/GgGlKh+PYRRoNQxAykJc0Bb2j+J5kOUPrLd6DWm8nqMps5Jy9m1+qvF
N5EYWu7sa31mmGnkHs6xXPYFuKqBc4wp/p17wGWxvuQ95x8aCRANUfVYXUPSliF9
RCncil54zNoYz84U70cC6/6rmDuvAS33tRgMHX6xtyFPcOLf4cR6Z5zYGlntni4v
N2is6f24swqmRQ/r0CEw9OdnxS/lPJwdBPxJv13yZFSbgboc3dVEki5rJxj8+Q97
7fCVeFmd9hwUvENvm4ji3c76pimYsqMXvWcJCV5/hMlMAnMNBB007mLpq2KW1kDu
NZ0x0C29CRdIOI1Z3hmX+A1Vq71p95+LDqZjJlu6inHuMRhz3wJ+yrCM9xBmI3Sr
qhZWToZTVjxztIQ0ebMYDGLVufZ9rJ7uhZZiRd0V3WLCJQ7Ftsup3f4jdUCUXREv
ygBePOtso+8Ipp0xlwXHyFsv8xsZ3k2WqGr4XfhAqsXFaReMkpcoIejYLxEofDxp
V9XkP2UFqNFIPIodXv0AR9ucVIdXB0Pb4ySJHTpvfOt7wn92l2eZ29D7jzgY61Kk
QH+BxiL4cMsYnY8d+2lVWF26WCMEPlzf/yRfkmgTf9EyCQQQCWEFfjU96ARL//OH
Y2iViGDkWNuijrfmp5angbnMH3Efb3FR+9khkFSN4Zi0canXFfaGgvJCyQfdaKqg
ke6DkLeUoWLol/3kSFPMFJg5XifIHsRS9j8S2hbaVIVNkDn1yD+Ylu+fwJDZp7uv
Ngjya1n0zsrPy9aN3Qha5779X/OaNnGdFs7U49b/1ztL3Zbx82LXMezvAM6f7YZf
iLVuy2IBheoWVYGHQmenQzrCrW/q885z7yau+AGdOH5L74JuVwhwp20fOJCHRjTN
I0D4Akkz8VWG0a7NI57ubL8pwWdh0GLLk2GdRMtOb9ILAsyNv41DGqEpynnIPw15
07EgQJTku9C7GSLrU6MoiDwObk025ah3F6+/ITpdfYMaErTgjpWFgHF2xOKYpja6
VdOtogCoShtFrqj6GshDs5jIQeM3POBR6Vx2zikxb/L55loAr744XIRKbwWYJrdI
XF2Krie82AG3zhHYb5RO4EEd8WW1YY4HwAlw08cCs9IfvyE5qFszK88DPRkVpV4q
NHfVw5B2P44g90gwz9MT9ESRM2hh58iMR/jpcFAcnNhPZk0sYmKlRyN807NJyv3L
aF0STam35z1JaRbKNV2NWQ91fvtHUt704jThXpJoRpNTV427Ixtgy6me4WZMVroM
9h4An5Z4K1SpTI6l4HKVMLH9ghm6VFspoXuyS2y/N/T+0F9nO1vpI0OfodwrK+OE
18JbDLs2+m5DXtXKPVRk7pZXr8Wjoh4w5NsToxvt0EyI8xDKmtrfRyNcOjaE7CFX
dFZNc9BjiqLVMAkneFvLdBr6T3CoV9YJouEABySbicX1+6cOreJp20upP6/XOyeA
yMwZCD9Zla0P7eApPwIf8iZKSzUEcg8NwY9HLbSlgvDg+kMaosTo3L69+exI3UQm
RkA7xK6VbOQ4iER2VhI6lBecUvsNxLwV0FwIfHHrYQnE5OHaFApCIbOA07haAWgG
2ShxnzfBD+H7ugFSmmxpaUROF5sznMYb7rScr42JMeNa5fx6KPMiGup10dEvaKIn
OrDPqk1FqZLo/kkbnQElToQ7mB+wyFKHeYshBFU5HXjbxrfhvMk8H5b5U5y0MeKr
y0vWQibQEs8z6ynqlqHFtHzgpbRryzTnI4H5nrtk+LoJy4xWFtA9prBd3IhtC8P9
las5tWE25G6+gy7OB1a5t8vdtfpJ5fdqcQJIZmOPxmbMxoC0hEPFDSzIJsV4WF6a
lw9SAgWp3gf4jmXEbPcD52pEfvWEmHRgaTzg0mu25Q8tLTyMytFCnXJuZRB+YtDW
72vVqi7eNmKTz4f1zg/kxcmwztz0TPND3lheWKLGeH6eUJtZiVg8QBro37CqnXTG
q1IRQFyNbhxiyOO/N7MPqAUi5N+thovUql79waQhonPVXAtNaOPhXDFu/mxyhS/z
zBFZay0lGPNw3W4hqZHIGs/3ygxk+BGAOwTqXAytGeqwubvlQUYlTaNk7n7U7uks
+8QdX2R0uhMeKfo2FMk0Lyw//h44G8pRAvQkkcHkEfESM8QGoqZk9gxl/eupukM1
Ghq3oAK4zwcTZhzsAhC4xwgNtK+VPSl50u994eiljx1DWyhJM5EWKGnBxRKlNfGr
x1Ctb29d/WhtWgcQ2EGavA4YL+KCxsA04e8Gm7xaOrVtsoiiFXw/GKQX/j488Y1H
xVp1pF4TiHRQsA8qWRRqcESDeb2keF2BytDyo70H9T8t9+j/YN53MOKRXfhEzah8
xwn3ekq9+7pi1eTQvUw3BObrgT0W2auVjw4jrY/1pVDssuTKRvoZ3Vl5Tcz4tPoV
tGFvCdNnsxajWS3tVYxnd4UjqzRIFyGEK+kg2hFQHDEu6xH/Ml5JJDBn3AAD6DJR
HPoeRBbVy1p4/26Yj7YyHdKujW+4LjNjGjRZ2SWb0jeGrIiH57nVaEL4KG7M3HAd
ierUaqpi08HZHVGdUD60nKP7NAPtpABgtM9mYRSQDqZwfGT65TYR3J/1ST0YsVVI
upAc1uR8n2pm1rrpQbxLoo/PNLk/MwXXl7SjAXxt4Ksfpw1ZUoO+SQhmJj7zgpm3
FXsPZVYwxIkJWcsLqI2UhMzZstPEhYYw4dykh7X8hKgXG7hJK9dHTZvSzrx8DT3U
1ecB77hEaynGtZYQdJT5mCszVdG0lGPivb4ZJn09BGHjV8I5ErVRjgZMYl55Pe2v
n+GO2m2xlfcqb937DvCfzdR+OHKJN8PynDfFwneKz+5rmz3r5k5cKB7ToKizyFgw
1oa7MkdfPmFaFTpuywYlXW9uFdZ4sXJ3TMymOcH2G/BfOz6VMZX1gKt7cYw7NvEF
vgECIqso2RZqJDHfV92cXWbhw8AvjWWdZ3/FMkXy0Itw6xoMoKOYB8j32FOiac7e
JM1o3oHZAmIpflegC8nBsr9T5f3vTzCQrqk6RZP5vUvjr9iRr6W77kx+1l64sfW3
Pfs8qCnbQi/l7UlthXDVh0ZZPcVDL8qdQd3EJqBbpSC5LJRfenc4Hyw3u+Q45e7c
Sz/lalvxyJ75N5oeNTv8putsxscmPeSgdvJNHgbZ/gCzZSVUgfsgys5yWqx8bVRq
RCINUxGTCVNC7aDPmfkOVv4hiHEYbcWmFed48ngTq5e+LhSUplNcGW4Ks2+sBeiq
2NAvLRFB3CQSbaj0Y6oMoz892h4FNd9tnqgpgWVel2tt0THvhPRLnF7qQ6WF6nPZ
hngh56bu+kd/KbP/U3xnucERNfkOa2sZC0sLxSIn41TtMPLxd1ZquRcl+cck3pPX
RE5yfajidNa+tv26/14IJLZ4JHKzXmsYG/plyq3RUZsV3HSJG4rHaCE7iUHFzeNK
xlzZCk8dHIeuahpkVfrIMe+0VDfn2k9yHY/eaqiEy4nkrG5SLycsdZ82EeIDwFKH
jKN1fOUuVkqGIsIaXaGg5tDO+YZ9ZcDjJAbhbmfvM544X4f+SgpkHYM3g5jefqVX
Fjazgde5S3iVcU9ZGzsGWbMCwPEklFcfgayVBcoYhvNwFM+XS566j7806aJvi01r
0JzPqdURmLoNetgVfV8QWRqqG+oYQOcdd692imgN2XMOHoXFioIp470ltBh/fw7x
W4B4bk2QWmamXKHqZ9oqt2ESqPcDRguHAxA6fNp3CGav/CneOgdUZviV1oHUlNMb
aSMbN/zq90cZd/Ht1StaPB5AJBV4JEDvNnVZZ/fTi77UE4Ibud7ydLi6ZpASP/tA
k00cae9NS7Bqs4P1Xfle2ivIlCAps16J6DJqrtKgWjT/0HlODR4BkAzG4JeIpY9R
Cf9vH+hLPFi2cetB/gjIB0nmlDDvRnbd8pdXsk7NziX2Az8YGnEQrsG3q70hNQyO
xWDLgFBV9RROcIpk+l5sRV9jJ9x2bBv5HjAa9hRfqqxI82jrFs/aSwvSyAEOtR4A
KMU44iFSL/p+hjYtDbM+7TkNO6+Je8JA1Slr2ZTa4kD6lzBPpP+tBL/WZOW8a97d
/1RrdM039Z2QJOdK16JWFBIOAXfJee/OLCWc00StfDsbl6dUlLU7mhuOYBlcW9Xr
sImlxFhnHNgDFP4mWr1kDXb/meUsTGAQmif2gTBlMRaicaUmaTx7EWU/xYKwdlBd
QHOWDJH2pl9zSi19yA2bDi3QOGrf9HYBZL6B//UzjZjLAtw/08W4rQlnH/lFjE0i
QEhuz07zSx6NlPEGt/f3PhMaw8wpWrZuIo4ZTuyDed6+2Wh9Y5bew6X3qQ2mOJAr
A5j6G1wVIpplGmHGEWAgun1WUyekYUKXYThnQdG8qqUw6j20WSeBmYC4AWU+rvnJ
1lVZFovz27AafXH5tTifEy0kDEcv0giptDVRAj/XJmbvLjOdhEry4udTomp07QIe
/nXVw7lLj9tYvnce03/egoE5HtxIxAQdTIuZmnPWO6VF12mQXfYfRLLiKeieGaj/
pZUeGEFIc0y/c3h/9enwgI8jBYbDN9WqGXrt9kqxNihbJk8JOjpkvCbKt6LCPxyu
hR+OttN5+FduJZ6jv/wc/R+CdscDxkFuxYRtzB7o9edcCqB6y0u5GRkK5S1+2QkO
8iFaNlmsVEg2qUJVREBXw9MpoN2b8khs6eRr3dW7sJKo+6mgAjdlxaCCbnyR5jpB
goWuyeRylajJ+RQWzml3knMOYH+6n7hCTeRk5xxmBhl5K0CMw0SjxdXwXnYm6AZD
P0f02sslUYcZiDv/UILOQxRlYCnqy8/mLqNIDuzFjic7D7AWiBv8AxvtY9f+ygov
ULbYmY9zAfNgFw6tEoWmEcqnSX4Rwcmu4ajXRrT/B5tyG5OQZWquTHz95gsyv71Z
SZlH45aLW9u24recktzGHwVkVuZsipWzB/theVUKviVgSlWg6axKEQx1rzS8U9nY
C9KxMgVVJ4I2IedP52vZNmh4JO0Mc+x6Cf0fOI8XmmP2A1Qqu3/uhLDCcOP/UVWx
SirPW2Mif+3weVI90eWLk8fxyHO+6LWC74ZVBRL2Wn6cXW02Bcp9WJG6pTTAruMU
H9sYV/BOtz/0AO5PGWzsBuRKLRs9oCC5iPOxO0yFMxu1xiH4xGOxAeGMUfQbr9Os
9BT+esBZfuFsf4SP4itQ3AC8AI0C6Xm9lywFS3DolOmwmQlhwZMqmT5gTxHDqR2n
XkPJ+OzV8NPpXHJKaRavJSPvLtVc4HppJh8vzZNTRnB6SAirVh1a/hc0Rsp2s0ev
R8UX3d/IByxypWSzsiVec6TGNKlSo5P8dVub1iyPjEtm+eRyCFeFTuMUvVyJROC2
gGBqE1vExypTzo0he/H4Sr/1gjCdn/S+NzBgpegCjBU6BBnktUR6mEnLBECXNxlE
7s0Ma+NCmDWDNdO0hN6zviSeVb6zSSJmgbpJSqaoUBSIet05N4lWJr92MQywXCU9
asN5pbmgm1M28jLlF/1goSXcHPMhPbGkLXgWYG68VNfBq/EbGVBXaCw2XwrJUubQ
mCfKcykdoIFCpYk8ncXz96oK3BF+Vr62HhOKL7ERhVZJm8jipUk32lfT4/nNd4bV
W+Fixo0YCmfaLBZfi306Fvcef3vS6qtSHCnJLN4ifZxBmI2atl6/BW0f7xLIwu4D
W09/9ofnIMEkul173KqWi3ccui6mH/HyOVLzBL8XeznFrT30UBn9ix9s/66ijjrA
rAbKmmvXojysSE3TTZBfp95vQANq5En4bQ4S4HC1nnJ3fXj3+7S5TT0bzLdfSvZx
PiJAnpzvRFfAYBASElrUAUreZlJd+rag3B2VM5nLr3pre+dw1VTRlTI3Crv9wwa8
kDSIR1blKixuysQT12eNFeDVblQTsAgVm6vKhzovMiql5VkZ4K88E4m1sdEQhmSM
ahjDx7k9Fyqj6fNnyN9dvihF4dXE4tVqECxAIU65Q8k/L6GljBzyUQzOdq5vn79V
fG5lYJFVKtBgAwUMy5ume2zF8umjuEUzS/Y49OXHXM/lL+VDARjN1fqwSxcF35Un
3no9+O8yPXDKa7QJ0vVT4KLQQn8uFM00I2EP4pNt8mhbed9Et2j4adtBBkv6riLV
sQRotcfjaZvesd+q7bi6I8KBjPfewcA4Rq2+dnxn6O3ajvn9gJSRuuY5ybZw+ORz
HIyLv51SC/wUQ4cJ3X6oEwRyNdab8cy8y4O2IfQePV/SYwg38mbW0kgcNazKUL2d
mEhnwgxVNfiHenzXdbRnrGvPM2fPrQaZ0heKsTR9EIfXQJOkvBoNVLCPH4/ShL7u
WjYDfWl/3NbNr38/NursDjPT4sTN8BGkcmPOZkB7dMqbZfQQ+M12HchtiJ9BYmqs
Zfi/p5CKe+kgIsLbNoPP9FUZAmZHqbvGJH+X9naKyVLIKCFUiPNmJbP1aaSHmyw/
fDIXQZhdGpZ7wlJQL5NeFPooaEhmyDV5HcPCMuJy1P/ce+oJ2x+OvjMRaQ5/mqWr
jJmnLN7EzaxBcbKQ4vKiepVzWgMxCIG3FH+gbxk42HVDNh09gV1fsMHQlgFiZ6jc
8g4b5Msg5cffmFR3nNcdZ9dQtEtthfTvPzB9hISL+UFz3HtwndLB72tkSkiqguhB
PUp+gVo1YmoF8p0O1bjtY18vYlInBNNUT7AOiVi1LtyvWwZLvneP+zXisSFFg2/6
eQK/2yhiqcWXZh5jqm4CzHg1fL/+cU3t/8eF6M4dkTAUAQTp9EIAJdhz25m0uTOM
X+9pZrrKuOrMrA7TjuVZfVyB0ExOqA5rO7gGzmrbZHLqhZCiC6w6tbVC+LteCHrT
JBUgbLhvVR8bAqhymqbZh2vEC+h67rlaNhZBGMRfEaMavt9CmHgoD8pF+3injlTr
vh6uwrIwE1dd3dfXCdKIuHgeXsAeBo3AJiOtgsB47KhWZEYxNxEzklru914K3rSp
LRuidhosMsBUB/l7tqP6tVKdgrxsF4nRKs9gtuKUhhGjcnVO5qvvMWWF6h4EqB33
d0a+tAAMvkr4S6iu9LpoLSoTt419+9jwang3yFaSMIxMWdwIpnLJI7NiYXpD57bb
xyFOjBW5zOeP/ytRF/LbHk7ryd4vq+PXEBsHrujf2JOG1OHk5m2MsiexbKbiD29K
1TypJU9gP5z8FbxTR/ahSJaMN6b7zAzJd34osVAKOuD60EraxqAaWJASCCcIjIuT
JBLsWlKWRS71UHaV4q8zFN4XqtEWtPVVUtY+rx2qb+iUbyQjg9Rh0AWzo7NXAX98
QG5r+Qv2AT7ypDj6PZDR0ZEMwjpePTf03Jo456k8Og7MB+1QxCbE+UPqBI0tG+kH
7QE3vl1OcrQhYYneVuF0GmoD0WnPQ62HIVFqZyJEQgyJIfj4yOCDmF74AEA2KXMH
9WfIOmjNXSS4cs3fScq+8nXExpYqPY5JV2YIz3uLj3JUXgD8wI7c/47ksDPwfS5g
jCZY9FcjSbiTURqeUAutw7Hu5YEBDVz+E7aS12mhsijrUqEwE1et3ws+qi6osjw3
Qvf+uKMOZUwCftEy9Me+um8pustSulHtCoFfl7eqWnbSQ1iow9AcJaAiYEjIrNMw
YKq09zM3UXTdMyRYejm32zrURWibEgpo9MR4/jPGwIGAGR8vRDA+5pAANjctdlpD
wgV8QGEGcx9gp+kptBZ/JS4Yk9hiDgpRzRS88nTUS/Y1pvwGoQ0/WjghTWwvFIbf
moMwkZfGHYx1L2S60REK2Yc6eIsPR+9XdSWpEDqoYxJ8LuX1G+rUNlasELpVLj6B
1rx2j19onNExh/7Bs2YGkZJWoubV5hqXwnQezvsYTM5fOskUl4SHLtw75ttvEuY8
S1Sk9nWlIBLKHHD3SOX3D9N3+4Er79OF2oBywkseczkmb3T3dEEP8mmwTlKJxU0i
LjndJVSpJs/n+nPhzE1WKZWZR82cK+klDjaL6qj1aMHusLGLPqAmawsFWqtVHsfS
QqaeCILhWUEo0DKwA3H+ILiIjnViO6amWFnA2I8Q+VaL2LQc0hVt8E4yQy0pzHX6
XtfE3bRJ0vx9SmaW9iz43CD4Ze2PIys0ePdaPdofITJLlFKSBZ36NFWuxujmvFyQ
Fc5oqfc9MD0V3q723U0mcUExVm2VCYvrOFwNRYSLrDvf7jA0oJu5zE2DaA1yoZsr
E6AWAbsdTQb4R+XGMpgUj16P1EA5euBToC8GN2MLkyaL7hrYy/g+oEbAix9Qr2sn
wtrqvoEYa7oerFCmtqSf1Og5oVWgXEH3O6RORzV4QXwf86Na8EYHy1gspnf/+6ry
hK28B3o7U4pS2nHGdt+6F/PGGVn9Mo7t64KnjpQ+I5Zc9HvvJEsaqk5JwF8sQ2aE
5wrvdCyx1pjpYpRSlmv8E1dBIoyyTYzeSm29pYuPx/7xJWoe2H9nyo6M/xQyVM1F
vUlpBvLBawFhvhZZ7Qex6Uh58upQqjTVZTKfEUS/7aT20Mw01WrAxpt1vVoaIMZh
JJP0BE1f9PwzhYJqbmrLfAtqqcYP8tE/QQWUvkNySZ3dSJq+HEkNfBj0+oTsqyRr
2aH39Ddhs0ob0rbkJY2C8RsDJZZih+OMnulUWN8hC/t9ZFTWgNxRSU0+YXxMXm5e
NLYI+Oc6cpH0mh/tYQdzfiUSKP7jopk8JX8J/gMD+wuzmjbAJ54ZVwxMa5H+9idI
L9x35oIHBT+ZM9gLep5DLY5paKTeAB3ok23gp+YZkoYgy/fXx9seUai1Wq/XPC7i
GpRDRLK0gGm4nVgqbj5ma5EXqXYaiGKiFYt9hYddIkdF3yscW6/W8DyHaJsvKGv/
7I91CCF2HJg8HTKiB8NuKBweuXw318veae1nUNCaxUxgm39oAPy/EyyJYIRj8pD+
iaHdllqxL9HBWXFQgB4NGoqTxs4twwzLqd5Tb84RjkPvQb8vfCht1tyAuYgUeNgw
fLuWaBZU3320cHDZissIPoPlk8rm/n/+5IFwv3zT+eIKC8IdjOCX30g8wx4OZRCh
r7z/6XdIaPwZyu9IGPc+AkN9zsZh1RwfhE10bHBquT/iOAjbzXYwCEJSBUQfdiNh
i774i88XvQnmcT2oeULz75qUIWsgCoW92wDZ69YtyyQXAN62kaIvJ0p7EQ4JcBpZ
1ba6/HzG5LumIxo6xTparEso+oHZGF8B0Tt4K9yO7bwyeDmMjCgpz3o8E/ZBm0IL
KRuV65IJ82fPPrgam905dgUPaSby0hnQHQXyJu6LwfwzQqd9Ci/GCzv6kqeiSHk/
F98stzRB0aQgOLelxnv1PAPmTTycO5K+PhG917AiDiSfnpgFFmtqih+zY0e/yF/g
sq+tou27MKW5mJYfFWI4hThrE35KRtEvNRjKa5bh63YAKPKTvHXXwUSH5WWlxzNv
iuaaC954QshfWY0VDksgYQGccOxcolZ/fXraZgW2yes7sDcBAWkYenzs7EufXoRZ
BuAxNySQWvwJgxLNHrbwZi7GTQSsrJKuensqGAhJ2c/ATf9fNEh7oGN8ow3c0ubX
ExDDA1YJlLLgC9f4TWKbo7L6M68zGlhXHxFftNTA1Vh0fgLDaB+tNVhdQKs4TKFm
YtCP4e1dd36BT0cTmeXW2a3CBH+0YbDcRBdl2hFq/siMGhx9d874vFS91lqGcYhd
EeNS6PJclLqtMy59tn49O04eSftQU+EXZ5ZjwqtSCKaFgHFxGoTMW1rC2rZnzezn
xTODGPlJ3prrlUZ5cWv8n4Zmaiobye8vzGVKJ5cX+CiW27bEnu3R25atEgbdDNZm
nEa64kQa9mMw1Ef3aaL0WAyONbuWRF13ZwGyg/CLYFTN+iTvUgt7x/Jadgro5qdI
abnEXICyWCzghRSqQhUW8aIExI2XZSogvin+2V0BO5lDt46NetZh+XTntDyEdmfn
Bsnzivy4rM7wA/sZY7PD0H2UMuvIYBV8rMk/u1hldh4/y74lLALb5Up25f4jW0gu
yxRs4NFcE3w4IpPdVg95n7aQ6a2h64uEDF1GymHBdDzqNuKtii9r8GzVX6pqDQm3
XILC7NDcTAbdAEk9VHLy1M11YGmqrcNoKaFxQe4RiKgJg4nq7njTCbd1BUgOHonu
xTO6jnxpd9WknJxLlFIRAlYDfg/ed5YiwmUUDov3M7eL49V2JZUQ8+yNaIVv/YR4
P9vHCN9K6fcQRr6UtKSfgZ/4wvC95c/HXDZbqGUTY3K1SbawpRwQMspei0S3iRNC
YRkiRLnRXd5nNaK/hNuvxA==
`pragma protect end_protected
