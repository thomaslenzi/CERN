// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cNN77dsE2r6pdPorjk9Q6tvU1N/wW/N72mfW4Yf8eVPjPK/PpIo8K/iEMinDsJhB
C2IKOpR+PC9rfSYbRKqKEabEPJsT+PumnH/uGShAIz7jm9d7jBw5rNd6eisju74s
I3qHwH+pwE/jD1P9oSZbvMw43jA5CDr09MTdNWRj6u0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28640)
f5DnD/r1BwoRNDlXuJ4iFMwkBNqLRJadi6uaYRUQUYeyTOI1PLbDdgLlSMNnI5mS
2fhp34GW64X7odKGDo/ALd4HAilYkaenC0nGQMPbweUO63nb9bsQu93Ar9XY9MZk
ItZBJkFQurOD0Dcj7jCMnVwUUKHdqBuTSt7ROQWjOLG4u+OeJ8Z5CnBGTRGgQ1L1
NAM2NXVo6zs0ZJX39gGl2ksEVRwDx5dE+ZDPSCPJe5kHtWSroMRPkehitaPyNMkY
MT+rJPqJIRU5U2QQ/nBfFa5uql5A5sHdFN3mThZ/1+L2q3du5BnaBH8jGfhIYeYZ
TCXCVrvqnNxC0dAhkd6igtHGKsTejwV1tVixOv9dvu8h2MPtYWBNkKcRPWqScj6P
V3fKe5m03L3RvRZodEgrO9tS4Ox//aviA33a4cg+8A+9eHnLoFsr8MClI0agUjTA
pZ9kQzd50G40zG6ozAe0eI9Bc/lweEcurYqni+3AqrLgl8xFyO6njp5tsNv49iYm
L5iOST0j7kpMZ69FsyMaqKgiO8fEj8xPVq6rI6nOc0iAxDJ3sItsWeFqalmQW9XY
WksXW5VQYtlPc+6t8yOrFkwhGfHs3HYHfCdXZ/BGzQEWddqEJL1nr1IJ2rZldcn1
gfo7usXzUJN9jIz4NUVPLSZL5tTjBCSsJg5C2Opy/OFlF1n/GVhk7SGT4bL/rFPj
7DV4ZJg7XI7V3LtM2MfINWBfSbuFzgie6kLIOZjWmvrqzY3Q4QvvOXYnPuVDPEKR
VN6FDZQdb7DOX2HJ+V89EDa68CsRdq1IrdI32LEOO9lt+pDO5cRwxqjztNCi8GzT
hw6bsPr7xSRWhmWSYsSYKdauyEFiOh6Cpla1CpnXblq8bA4u69/PJFTWfB+uJMq5
/v3GMI6yp/NhRZI4XnssRVfOeFZGHT04H0Smkb6P8Tg2BV4Bp2x3vqsY7gIlNHfm
VLZRXHE+DVGJPwwnEZmhLHKzQbMdNx3GjaYBzaa5zDMs4DZq7hbMi9n0K+by0Fjj
OdwmVPxaLbhNlkXDh1ukaxRw4pioGcFIroeJHddA1m3lRI/gf0BWOwkMB1tmWUNT
wKY2y/XSVmfR+yCdFwqgr7SwOX+LUj05+UZ7Fo3Ychq/k57oHjVCJj7juWRBpKe0
PyilF/0K3STdPvtJjwkLrIo8OdExNPIMIYRpcUN+hKbevde8mD2PSQZLjulePn/k
W7DUgFPtVGKKB7wsh7olvIv97CaRhW87jMZIO717sA8xQfVYnRX738sg9mxYeI8n
XO0qfP0iykamT8RY1/wTCTvQN8H5lNVKv5jFdQSKSMkQju/Z7sh7YEYFekjAbWev
7vIsPzE4PRp8nVEYQw/cHWgjFHQY4GVcMdjh7Kp8wlh2ktA+JocmiasXX/o4PqJ8
/JmqW4yUrM6i0SuxE6jbkAc+A7YI2NDjUSh0fqRHGjSdMDItNVvJPrKAe8O2KE/8
63kG6R25g4Qdl4P8VKP8mJjoEtHQidMy1MyrBTO7HoKxVwZUJxIdG+vQPBvIa7bc
Ynhz2+GDf3C4IDucI+1q2ahhh/cUWUvcH3Wwwl/pJ4PmiCKs+wwqvVwzXeRcHi05
933ou8XMlKYuCDSP9XaQogu/ZYC8xG6El0lSwAjbk3lrBb45dVgNPRTlIWqhGwAo
cCVgq1k6AJ3bsbvwcdJ7Y/DFHo02ajLK0dMx218Iq+rYswBFm+7qKCG5ESEGwiMP
Z3bVoAtRrfgdt2+XncRGHeijzHI5NvFjDUN7hsgxVYTWswogZMyxgeZMk2ftJ2Jt
TePTUeFgcNAMy2UNoqGaz9UhJlM3dLQOx26X35GFsjMlmVDAr60jsc4Y/+Uu8QnL
21sq2caiqac3G4uGWLjCOTNnosqii8J5aCrHcPHreJislficNNbqYciXIhzbwU8P
8YenhOXem8/YjooJvErEG/zr/ZQpCKlo2VSkuQoPxWnmim80GCynKCyt0cKyr7Co
NSeirm6ImFoREpj87Tx1/uqxsehAM53sBT8vBH7FpPLj8kk5f4V+RIc2iiW3CjfH
OxDG2oCisKvLfoVi8QY+gIG4AtXA4ABzs82S62gMcm8FiJZ5poJSdvb9oYv1w8Ks
HF+BpGyXkBxa7E2xVVWTq7B5HUnTkjCj4uNnJBTydi8OSyH5uYEv1TmWbiIlGwdX
Xy6O/SUUDAK2ich0Z2QG9apslfHMIeJWgHktB4K8FbJHrQ5gDGTJB6VtHXAiVD7y
VIEdGjubHs3mBjtLKefvUqyBoJPv1vImxPpBEqGMRbnRYOXMtPu9YbSZifT6ocDE
ge4xLrKOdTKS4hwKLnqNoRZnRy880hvkPYGaixKy1CqxY7pX3n5WIoErLslBZmdr
b7TkNjpKEaxwqwQn/eKyhA0Is/uZlEKEc2o67xpAeJQ3SY55sXxUC4608f9JRRyn
fUxRSXe//SeO3Wd0K9LhuYaY1WkfBCDclFdW1IHQBGDfhKhenuFiGFTF5poQFXaF
ucxplSC/P4Z7ZbkzSPG+bxUBwv9WE8Y9cgnxlM0NVhi1eEbjb1NxkY9cC3ovtJxz
VTC3Urss5XrYKSgLEC/iR1JSXYLoa1Fd+bK4F7Ux26bYgWom0e23A2k/XBza3rm2
/fna2Oqa2UeCP0wY1VLmIc96YNitxwhNTkcSUQyiO0TuSPHD8Bmzw5P6CeiUudPC
w7HKUeVEIRjWk3di3bVITBmbhAaWYfkSpSlwJawjcTAOj4maHDCjnFhUnuY+rTcQ
6TEI9XcDY6jiEVabPoE98L0fLwTP/VqdJnlSwDb28cZ/6iA2nfrmMKveua6mjP0F
g/clSfM4AlnDuKc51bs5FeXxdjkS5uOindhQq4jpjxxKhVGJkz5rKgKd1woqua6m
YAaJLwFKrHjqK6luqwO9MdC5jVqzjyXQtfcHyC8UWqi7kpeuye2PY185lFB7ODYC
YUlur+CskqJ8Gq2bSOrpCfCxvnldknd48Oj0BckhaO+Y+av8KxEJalEc+Oso8xHe
36Gge6OATfF9WWru9XqcL3h+X+iKr68tkDIaS/masLdTXdfkwcCmdmP8NpBhOe9Y
Tmhu48SWm0o6tRgXNHJH9OZARIBkpKIqP5xAiqGxXwln0Ez40EGWhuaS3JfMm9Hg
F2mfIlsljQYH/EjowHZftTye/NchVEU2a98E+wc5dmA0mBzWWtw9S89gtUSTsTxm
VMPnN9lhleRdPXjn+R8xy2FwniALYLVuXpOxNOcmrwTXcitRdNCoGsNIZO3V/Dm2
CxfczTrm9IojFt5JDXl+dFFPJkQNuEHSuB2WsewNBwuKqcvAPUc58g8MXtl4Uyog
ZXrMBff6xWNA/HmGE5vTEFBwEDS1BLo63EJC9lZg8EF4+TUp7qUf7pqj7Mcbr7jg
Vj5DjemR0LkCBnYTyomx+9bw0Q+n52SWEsIXxd8JYUZ25dmjhrM4tXh3G7UoiBvK
FGKYFdqMxeWsX7NoWxvRWC5v+FhSnYMVkb7/GBfQTLW4bOetMhebOxDotU4OBSuG
NjAgMnEUysT9xty9jZ2taNXZ552ss7QY0KgFjwYJncLUXaetvqsloR5Ms49MFnBh
HpXO1w/cuqya3uBL9HevQZRYRat4iV/7G4VFvhGYtmZpdwbjxcNZWuTirPRrvYxT
BvyxJCQEzhLwJipFTLNxuw1xjbvrz8Em3YhflFG5YYN3fM+Ajk7jj+Q3C+adQiOT
xXaCbL8EK1b3cjNxTHb0Uyqueb94gDgNdWdKNCXrnlZ+jGBJMPb6RMwoBs36RYwT
zqcGv5Ydww8YqMuy1pYHXOVbg55kE1qzFtmqYRoZb+fsOlYB/Vdf/9Jtpcvj9t3O
PhvbSY0pyijkhf1wK9K0jHnTkCACwduoHqtY4G0twN+VCkEr9/oH4WftNbG0KHKV
yjiqNvPOm9/rwVxywLxBYfTNExbtc7Y+X53s97c6wHvBzWNwXW2GaPupYW9kKKzL
lK+KqJxupwZqDCT7TGvt5w1Um7Sx6UOjMFTPSIRLBLv1y+5eTwuJSZSr/83Lu4nI
aBo5+kfC0L5NpBgS56mBdhn639QxdDzboazhBJ1dqCIUufKFFFaunbTYPgLWR8yp
23yM7KezDrFplsCy+pzWUk0pTPbp6ru9Ed8U50BCq8USJRnbwrBCnoWT8hDDwQJh
1Ou5VuPg9w2qh4BXd492uKfMXTuKUiz/B++9moxq79GPJBlfRBmu/a4AOe0+2UE/
yWavK6iEBvDvNURnlUnTrGGqLp48a7Jw+aZakF67QBEO0w9WU9tZ12+1M+nMRYj9
0oFxFSt6dqjdhyjMiCyfvyCBbrwwEtASUbIMkgqtg4W8Cg7w8zIOHNm2ndW65NEd
bROEWlfPqRGJ1tTX+wl5iJ4Q7kW8OTNK6PeGo6b5VjOpOVCZwAgfQBgjL3n/lpG5
3SzVx/mByF2MxR+z2bWTYPpdGqDEiarMV9EMBUA7jxsKunAnBIyNxs5alUQApn0o
yFl/T90xkdfrp1+jh+mMf0yQSC4SQLyLyOWzzQhMOYPm8adfHvUgzgEF/HSsjzFH
W+aWtETr59cW4diuczDatUMLlByvv66bKDVaY+i+4CDVjHeW316dQtRKNnnnem6i
kLCdX6o20DqKDEIZOsEGiv1qclC6JaICYFuD0gJZc8M/pqiPWXpkJwuFuZAovglx
LZS3UOxc31Ef4BR5toZUnjYDtEusvBqheM8sUGCF76mg9O+NV41+DPKb5n2Wy6c6
Hh+31n8mLtwLQC6c5JmNfOcNnbMnuBT2Lmgko1TRhNvyfjF8KSuAOWH+Jry3h2TH
GBpurI9/lZ6kWLJ/5oGnMg2nYg/GkB+c/BvEUoBVpoupIL3d8bZC5TWQG8SuOHYl
gA3JdnvhxngArqEOTpwFjDR7KGKdQ2MnnL3/Xoe9hC8iTPLPPvnfc/NzNlTkHCNX
LOBzG5f/D7z2/1dBRMM0OItwzV57Zdk23RRNA5ZiNcx/WHJHoHcPzf68kqqEMxcj
tzfqQNdBLBXqdqXGuS9XS0KDLMa8tDvearANxO7WmbSAVSbyA9l1jaBq47kT+ytD
Id+55E3wsc9bYSSSglQnuEOPWQHavaMNdXdXrOGFCBARCzkc6WnWQ1UdczKHSnHW
OIjLKG3F9tJNrq0ZqcuDHubfGXLpNT73JqAATeJMGnWJCbMVcJEYsIbNDFvb77Hj
QL3kNudPvsF7Z6eXQR4zs93GGYnjVHN7XHhFyoOd54vo3qNA5/4ovDhReLbn0CN8
p6m8ksccAaAyI6dMe4ipuQ7SQrJjhowxagQ6zheYmGz6+/vcyBXVTRNnwV9sIUyn
EMnhpkT5g3LxNrD04V456s893dYQcFaPBJIks0CBgTENAL1P1XqGM6dLcKLA7obl
jPyLNgaTJI3O9co6HC1bOyQk67ey35CtIe1KymwWxW7D1tRNF+LXeLipIEJRXTNv
eCYH95JPirobZJgE3+lUqACPZsOslNd57lVpMVr94nEWEDlJEJI0dF5J8Re3uZ8K
QdjGx6qtt/fSp3m0wuvM2uw1JOOlT1ZzZxHeKmYBXKzLLDuSXKEV29Cceep6nw5/
UsFpYfgeW30PQxkLfxYOegrAUD3El+O01Kv9Cj24++WhdZZb0DIjhyciGsDG3ct7
yEhjWpjrkAM9/aYdqg2FJO9MpOfuojPuLKK8L2GTvIRpusDu27EuWEti2M/IW+ml
OKfTyIMPibyt6AyLKsD1e8i+UwK8cutfidMYH3FAQi0MfJa2qh2lieaKDGViJqPG
8ABsgx0l6cS7BYSPC61XfeQ+AJp0Swhk4KdXytyaZTQkhhdCXaWxcTr5Qc/ZQx47
hZLndR8YsS8NsS2trOw0cW0dokuKnSqksgZr5ZbsISp+PRInB68bS2dGYSz5Gg3L
ZZ7WYPaFjl2nk3Bu9yw+TzS4bGHwM2m1ZLIlK6LuG7vKYekltbcq8iYSEYHjn6M5
0cFhEB38CXAni992Gu+mc+Lq7LYI90GKOmUg7G6LX6n2iZr7ihseAVS+DCrtAMkh
uC5yP5F6dXBE1KuVVEbFjB88Xu/+yEy1KfKlFj9IICbhTrfjaO0m65GgTEfkoIHR
uXhDHzWpDBG0peApUPm5F12iG5SnUeKGe/wDrBRIOE1YjG5xSrdJtgDwgCJhX/Kk
4hBZ5x6X9V4cVLj27WedowT5smrq9dm1fqTO3K4+pcewk4HZb1xh5y5PDwvmJkhG
oE1kx8E7Q2+R1VfqH6zWI5R7D8XWtnI2hS/hd/y9b6OId9O4IrfN3x4126vc2AN2
gUEUQ5ZVH7IyLDWz0dlrbzhJ6Abs2mIuZIX8clEHn4vew7VcEXbvbYTVndNERuJi
MaqRuD7+hvqdtLTyPD10z8JkULIpsLFb+LYeB4jYGVJpOar6IqU7sbb0P1ZS13+Q
tEhRw9hEO6ZJYT1atqQkTZY5v0VIzT41+4RlwT0ZhDEnv2z5x4mDJdWhSne4LSsN
F31UeIDuul4+SUghjo1W6zaWI8GMMaMVQdvPWF3+o98XHioN2GjmcXMBCQbyHd4O
l4/Nhf/9/p+w2y/S5Y8z9mIHi1MV8Ru6wU+Hsk1q2NxNDnRClSVNzIW5aE3+SQFw
fSn9SC9CM7ZDMTbY14MIFKzIV7gMWhpa6+UDoVlR0vWHWWzp5lJnyjmydhCI7hXE
9ZwFrkko2GpDRuUt6uZd9U0y4kHOxaoGVsB2FnA/jm2Vg3l2Pua/6YDS5Z1t6Z+C
BvupNXUQxnia+jWg+hM8leD3hHLQeLlzjoQUpkEp192kRvs4bmSU39g3TviuO4+h
rw8diVAC9pQ9cZ/jtHaL8DJH214wtOTBeX6WgrqP6ZYnvDYt3ylQx8nmN0CbLXrt
Cg6yyehlOTMZFQBTNy863QFN0FNUna3YxoRZj+dmsugu6A4fb5iyT1cPK6TVMQ+q
Li6plWQjUS0zmmRFkuVCEeZhVydER2+Bd6KGZ2axXmKKIqVKrXVjcjWeU3sO465N
YonJqjOXx3VTfr5v9H2KBMbk7nC/TJ4xCHCYHh2xmrEl/PZ1yNtzjDo+6LqNb/KQ
vgymQWUNXMe6lkgmdP/FSqAdU0JzoXbXDzY3Ujo//iX2cQiVlGbHrt+K+IAT8qp1
r0T63LMfyxlZAJDqKO7K9SM8zPpcBltX2OVe7bngdMd6gHU8s0qhZsPPDsTji+og
S3jvl8q1u3ztfSYgkESISIt1yTlIbzFfOaSXjjLQKYg0KR20dr2KeF4+PdDIl/MA
Azi36zDPPu0PIRJLhW/eFTkWZbozt0RMpLQDLznvYyOv1PBy7+UzQMjVigixTrUh
bJ+p0Zu3xIidsvQznFQ9Yiq2kCQluZ2MNKS3LanAObO6BbXxGdEt1sqwyuaR84Zs
wLtRMYuQfzDXU++1XPsWpU8WH+6SRZRMBwdb6YICAAK7GFPtMzBsx2J5LEjpWNew
7oEpDxPmlVgOIWO0FemzsjftHTjOCrkFqGvSJI5WPk0IpUng/HNyNBuIiRHFGbJr
26menIPTC+8HomSHjwn42PCLBRBALnySkCb9Ecj4BOB0zX+p+kYiQk8CEvHUvLZ4
v/0eSJpLy4EqKh8FHFxgjieGpCd8RHm9guoyCuP0noBhGW/En1Z9BYa/07MtV3ba
ay0BNCwASX0RCxlojLcC9slTK2UOYX1JLiUygB9iVNlUSNIAv6m3KYIk3ZDmaaru
R46XEg2XlJrB2oXGN3VaugKIxlxLrhjpnUjfpZ/dfx5WBUtD1FgIJrXi+3kOIsjI
jjt4qzZnPng+pMkkKtH8tCKP8n7y/5vJSPFQp83ZDcrDkt/Po9ymRcnC48yjCoOh
iz28bgF06XG4gnBDO55AdpC6i1+PWMlL4LFX4Am1eCd7E5OP6lu+aRFLAgThuV99
VruAiDrryAIBdoQxGSyGxLZtlTM9Cn4jbBjVdowCqHTtxjFku5hfbJL/ZWAbgRHa
fg+Yzl9MmIyF/GUT7z+PFohWT0QOGv8o6zTwCAjgH1NveowCfLB87A7akSLwsFyD
NVJArUjTj2Rl9oS3NeWCBqgMZKtAvwR50cJ4CxeQUdzMJJiM1s3bzdh6tzCfVnW4
dMId+ZZLlE/3xRujbVyc9OBpVYZZwGEnJ23e2V/+Edv5nKlvW5od0HAS9n4SV5Cv
tu7hpIs6Jiu12WcKTHmZ6GoqPirF5NE0VGiDu3f57VCUnhB5kBm4+HKEDyaolZM3
Jq5prePWQpFUDkt3NJK/Hnm+ZejpwP1e+Al8U0w+iyn2z+Y//U3Bsih/+VJbThho
lnSG2/+j/imRxKjOFlxYuBTHDS4/eTgwvkpqQCmrdb1S7w93ReXMkoHQ7nFEN7Tu
lwPrJBR+QvUw/Ww9hBXT/nMiYjkx1zG/UnPmpgo4+dmBGjcU1UqYUREcNdzHjr8D
BpnYdMh307NcdjdFotrj2rWIWOUXuVG1eg0qilP6UwsjUKtpdQzM+GMJyjZGMCaM
i/SIA82Ox59jG13TE5V9pCFzOYUUTs3+lsy8c2gx27Imhtb1bAkqjFrADhJCYMWs
LeTGdt8jhtg05eC5xO06ZJeNzYWGssicjlxjR/EsGP7RqiB2gul1HCPU3LhocyPP
JnD4dMVTT/drLxTu+jw8vNlsIOWtk0bQx1+MsUHUeDUXo2TXmCG8902pQ4hR+R2+
ZuGr7DjEyJrnwiNmIyOmq6ccilCAYL9Oy7AOekLOEcYP53yIIHBfbJfd3kb1ssuV
wGKhe6z1e/Qd365WPWgbw18ZRJt+vsFMkDUoy22A8pQTKSxajUXa56HmpoCDOYcK
crg0Jb4oPxuNRpO6W0duXLgLlBXL1u6bjVfTvVrFfPEw5No7UrFCKA+6NFFInbU5
SazR2IbdZXCBhfZF8IZSkZsEQ/BQiizqZMx/4WUjH517VkHuONW2RzTuTe6psPaS
VaBV1i7FIWef+LtMMg/O2ArPerboH28wCxQ1O3zDDCGLhJIFZny6hsZULnFWwRLf
mgY8GLJsBJV3fGRVKr3RzGG66viXsM61fZWjjxELL8Bk7mxogw0o1Y46KdoO/ZwZ
ZRf9raoVnO30p5EBKpdzuCRyuASP7208VYm9TQ/9fiE6n6yvUTMOxyHvL46VMhDd
W+CFAPaspd2WX8vszAKYCGFujrW+nw9vYGraVdi9g3QHvYFq2UXUsj6I4OHQwD1i
8f6cYvhePpS4YDBrnpCHlB2nbgoB9lnBg9u0fZSy3m/zvcllg396GS9TLKsjeNV2
27keJQ2xFY3wV8+7aTJaAn5GJzsnjEFMk3RJoHjijNC20AlelmYmJDrXfAzKHqJU
D6omkccWv0yFOuZVl8kcoSEMnDJooYoPx/GH+4LCw8XjIjpDSrNxfv3eRqAhe+nT
N6AnoMHOS1bf//HuQFL3VRI+nXKYwkp96gDxeNpzY9wfbeW7hgKNbNECjJwfaj2H
GGJEIJ7mLez21mDI0Zprbz0kNm+Z/HkFa76l8gTw3JCuqzFYOFOhldc7eDsakXcZ
VTBDW7r2xAwTWuTANCV/qIphF7F4cT+BE9hFGdc/R6I+nMxWPYZi4nx2GV3b8Nby
Vyr90tSI1ywq2gL+vv6L1w3fpu/xSq0gcFJZPmRc22Kl7pOxygmcYEPIUqf8W4T3
Ytv3+xvKf1GppMkz4N4Dy9msBq/0W0FSNBVLadSBE6UcxDNbOljNFF0QNz0/u558
gOiJvPsVq0MBRRAr7tLRZRfSLITMJLN6xmRXxbV08tjkVkfDVjYSWNkoaowMMjzU
kTJfz0gFw/bLA1pEUhZctz5wrpx8/C9HwmIb/b21ogGI8NxrED9Or9Tw6/U41TLO
tl9PqniV8ejn2juUScXBBquMMfAtssFGCSRbwfTOvdfvZmV280PCf85DeceRMyim
FqFVYsCVUjRPrWzygFGJCrKjCpgqZpDSmBJAufISSJ2xpKxQD6jU+iuCl6YRKU24
mptvUY8V0j2O7Kp4Rg7THGXj3FonHjjUvBU5U1tNfwdsEBEhrnWam7Vz21Qh0KV5
GFNP6/xnPfUzbmSFy+0qi0uo/EkccjfbVXmobi1iv/VA+Awo/3PZKENzSttz6QMw
d5M39CqXjxjrRa7snsVx2vi+3AfOdpRI1WpyPm3Auwu7S438/ojJBZiaXJDOMdCh
xuB7tBl/MZvxM+hRbSs5tu1qsZe1GCBFnvQjJ3KMfovbjcaV8Nu7u0uNMPJ+aME3
BUROMvhnOblhwA3A/2BLNJTnXIhO/N2s3/7REfRooqRuByrhblywpZiSCSNwvQ3i
wxPISjKh7dS4EiizCZafsKrwjr2xgV0bD0Jgo57Hn3YHejUCgnOM6jfJaHLFoE0m
6PD1a0eD9opGKVt6LJDsf8DDEjSVo0I7KOnrbJ63OwVhpIvz2xPSYERYqn7ZZlO4
g7hHJU7abSQ2ivFrpVTVJGnpYzlswWSPUyHy9JNOyFsGL3dCAxVYzcOaX4PbkhzS
wFhLsN2mjku2ypUmQFIY1BA1VQCEtBCbkOSBa98hxPSvmXxuAQuwJzCx5uySHpWW
Y2EftiYGyNc8gtLn7SeaMxUJf5Gce+K5a9ZKHijpSBjV4MW4iQB3wdI8g9l05cXO
BvuHUWyV/Ws/1qaYVO5D6tG+2bJBJrv7TlnwuVjKTU623mkrQ/jovXVBx3psdtrU
NNgeODquj8YfoLN4FIC5ifOo0BMVuM0agvhrOQYZASpD/kNqtFFhBzpkbShZwBtg
XS8SDhcYu47MVqPMYJ6fDkVj7WAccF0g4YMa2K3wgIOwxLU9ceLamDAEv2L/K8si
2kC9GKF3wa6xRgAtajD85xqn6yT8AvfP6lQ3HlMMy3qH3MJkUYeOm1n0V5K8KhnZ
bp5g/hkDVbbzZZcPAUnm/5QgQHR1psKwQFALK3hYWyhxM//Qa14g1q2IP5JP4CQU
ew/GOZMtWAUj5PWMFl9/f3reiRhrb9hk/1eYflO89Kjj7Wm+SEaWc3GmZ9ce+4Ye
qXrYf1sIk7ereCyrNll9NicwCIqo7n5891v2klQ7yi5nfKVNH/tjz1l84FM3CnQ3
NglLog93luNfhXjsGogYc0UHzoKsyBgs3cVTtkpVp7DwE9/hrzNZ9g+HfvUjP4UK
z79NsYM1h5tYZBYBYodSdTHMcpFtDJirwq/0JQmvbdyeFu5ucNiWDBCkp0j/+V9S
t3l0V6kkoO7gStZhu241otZxcxFrW10QLiJek2lcIGLQWHf/LXoO3c79N4M0ZLgi
rIIDTUswTr+s5EgUqkcCKlsvZW8ThnyhsgcMwpx1vZT2n3Xc+ZMYdMKLgs64GvBP
vMezjpKIHk/au803TYTZafs32yAqkdmF1YTBjfR4xFVRWvbuvABVhESO8tsek9xG
mAsQmCVpH7H97gt5MQZTS1uS0gvSigJ3pMU/cMry4HK+wPr31V+eRAQQQRT3ZwyD
PHFsIr+N+TQUDla3K2Nt/40BIEb/5tUEumbQtZgkHM8aKzbXAui1IJxty+V9OlFL
vpS99d4nULkjkd48Cb8owsfKdpZfo2276I0VnVyBOOBApF1k5OFxlz4aZkCOva2j
g/bF+Hj3zEtpDaOz/QY+mwP2CK8V5uiRNMvWyfc1K1hUEsX4XR3P1zxliI7S2+2E
V14u2ugOILMfQC2BbuHesppDbNI7xdUkasLfjR/eR+6j/I+dM3CMHXUWMOvMrh6e
9VbIDtIdrRQ8p/gq0cS1qFNzoyQRW/fl6UO6Eb7j2LSlPfibk8sWBl7IKNz4hMWt
uyRFP6E9qaRffxkPPq6gIY8ujcd5oL5QHMkZmTvt+CnbDHm7Zp/l8SISUhEk5Wzn
xHd/6jeWBb4BE5gNhppPA0YS2h1mYjVQlhHvI4lxDN1DCG7y7wAUDaZ+0WIRdLss
JJXbRJ1FNV09FCRzucgarlWlYUYA12nozKnIU/TUc54fRoDQnl4smXHnvOy/6mHt
AO1ge2y2n2ViwN9nmpIE7bxXK7eBSrWdmTSZM9VbaS/efM/dySaR3+2SL+PvBbkX
t9NKjeDC9JNvTLNNWkYYlAm8ocsgtlqbU+nI+hZsx1wroV7AZuW0p6gbfEsVbtBH
QCDNkygvV3qHHy58YxJLV2SuFI0GZNrZPqv4PDmDZpIuXq7D7WN35uhlCQAEqDF9
vVuu45g3WrcBZYe09hpXOu+1GDGn1a3eqjo3f9MiI8JjoWYsQlkeqzFdq+clBprY
gDCaobVctxOUsln78qiXzlNh61B8xm6mKVmZ/8H7C0J6y5c/PYplGHenFIAfN/fV
ywmIOsC+DVH10i9qW8Wh53KSKjRsfMDSXXXA8B5+J+G28lJ6zi4Gy7f3Twt34zEr
WWcIjS/r/7d+OoEkiRXHhVEsu02VuWHmP2WQQU4xbgtrc2RXJImibkEpNDwth1ap
4l80+jqd+94IpPB+D8qj30EKrOBQ8CLtzNkfmCFR3ys1Nbx5ezm1SnilffQglSEt
OIZfvJI67tnu8fnNXwU1j8Y7SYy8PLUSOFhVh2bcKsPGvlnOCWyIp/fcsFTz4E/C
ykfwOwjLFDLyMmMhWuqzhSymq6iQZQk5sFUGLZAFrG1LuBbRLN5PlDgPWDmu8Pox
/XUaJGMvYnO/Md4v05+PLU3qoKEshoqDRJFeLNYZlEWxsawlMBq5xN4rs9KYirRX
IbDYGV2PRr7DGUZMRjpd4qaAJ4F9jDjt54hxJQ9YW9xG00iecVm0xOGr8zxcqi0L
0avTl7eIra5kEICG4mYKar/zi9MTljDvwJw9VjBTA1Ldi+smNSG2w+rsV9WkzFJw
cVNuyee0GEdR/OnurrG4RIk3rjrCvCo+2DNEwwH8xIIC7MLDR0JxkUvF4S/m3jfp
tIku2eWywgX5Hc/3jzC7G6rlEe+YZ4Us2Z8TjRBjDe6jr1QCW3tzSOTXGNArKlkY
YDMhWPybJN7MFuglb0xef9UY9jrWmucyqUwwfEwEvTMJE5Zi7R+Go2vw0KMRnBts
wrdkcGt4h2ot+YVOsVwdtiLYMcDBfgx5sWaqacIdC7SVTLsekgl5G8QqE10KRU/5
hXagOU/MJrwDjgjFzOQ/HkqQ2df/aK1RbtN+5ESDFah9p4/DTyQkRYeOT+l77r9w
lGf41qz6Ej8OvhwyksKMGTNVBESNR0aUQqHQAiftmDVFNF1DZTWr7+kcKk9565mh
2smfLqU/sthzNvcOTJfoShVyAz3xZTzpAshXbGHf3YkH5WWl0KZSuYBDIgkzjhMV
s1V7EJrzmKjKHlclXwKdbwvqjSgBHiQi8I+fJGiDDSBO5JmJmkHQVo15IqNrsfSO
K7T3EIJqvew2ZV0WfCWYP/pY8aMBg/Asyg9YT0Mqd/QkUc6CD/m1/ZVCJNd7I6X6
msgQgEtxBmnViqN8NWJQEP5+pztN0cZ0n6hmewz9LYURF3m5ib5IgqaZGXpk9E4C
W6NTWm4+w32lNYTU7QXEpwTYKL8zbUE4WCqjYRAZq9CY6oDjYbNhDsHK9izljx/q
NuzqBDHQ2gsLFPoPW7wXBg13T7ssU7R9P37DIRO6JL1fr3QJRmnAtzI8DcAGaOli
bl16NdFOj0OlETpnkGIXLpgQr9PBVwXFlpl0ZoDkBrChI8k/XUbudyB8DnNvwWVg
5A0ngO1ITw1LhX1kZJNErnnIgLg7zomGkUgJZLAmRbvKnspLVWXwotylPTGn0HYl
HzcxTdX32UyRJ1/IJy5fNqvLnS34BHBPAmuFEZ9Eldw6wr6DIjri0JyG0R7bVzfB
1QaLZTnB/nOH3C4rtJs0YDKsHMwMBxuYX0d7QBMz2iF/TB4UBQOj3qjDP4R1nlGD
d+tfkvi4wNsyK/dvcZsv7aw4EmlvAb4GK3bLHjsf6VxluvCvtiHb0ntuCDWyz9rF
u7+vjvchirfbHtDZjWyqlucHdpivSRnW2m6Q7pKVhSkR76pUlgQFmcskdhNA9G4v
7Gv5WX5s0vgt3kv5hotqUNKXh0fDhjWXVlFE04TXLxmP5zz7wBvbnEKYXkSO8org
3WJ0jN3nlkPjSvxX1L/CsP3ZCNlWNJrhd04wRRs67PtD+zxNxYUIsAuR0n1H7ESr
LqiRcT8T5bHnwXGPVq+5tUjxisieBQGrLXU66yBmxm5aJ93Fd/P0rNUejogAlbwF
I8HDQ+kDE/5CZjzYVmd5qT61efGvVHs6Ei2Jyd47iX0tklvlZJa/kYi72kwUMNM8
PAkdlkkVJsmTVYs81nL3J3kX+DkPsiRAip5PKxQdAQVivpZcHmaEg50h82L+RKWo
7kcjZqhY4it3B5NRNYV3cjPN9VLidYHaK54StahrZtslZgNjxtdCYz9k7stn6Vz+
RRxGEHE/REP32WNNiJsQaWuoa+2ndhvKcQesm0QzMoxWoQfYaSgEx4MB7zvhOKGv
coAfZVZuBnxeAZSDdknPjchmTBUpWsS3RCwgyuyE+TI5GI+DoFHrzgxx4a3smq2e
eSEzs8zfdIZQLQAK7c/rj67uFrRZCcxho7iYfW8G29t4Ul57s6kwRIe/oMHEnnT4
JyUM+pom7lchWjFSXiHhSQuxRYJaQSWWFjEs7cxraaUaRoFxDUjl4DWfxBYD51Ig
qthZTMYgZBf/x03/igZlu6BS/ZR0DvHx2HyXZ4CXYdRQhutQpNQJgj7lNHYcy4J2
HHdV0gYRGruqOjZNrhF/Hspo8UFbeRj2QSqAkzR+GFQ2tVwaePKwqKfIfEzFLsyb
f8TNrzBVOIH7M6CWCPHqyX10FV7kAvR5iiWwwaSCFRFZ5cP6erRbVRR0QyThDVNX
PePT3QgiQgLGgKKojkmbFdosVxwmnTcw9fOncqr+/jtSsQnhPayPYA7WVDusWRee
detIXrDAKTMGjE8J2nRFWmk04qPqPWezmOZxaBPZm9Y4xh1t8o01/XQ6VX465fvn
vcUgjnbFqp5qbUqPpflTr3vlSj3WmC5nn12QWFKVfxNzlsgqlcsqQKnTFsIB16+8
mao4qp/8VCrmN1BDenM/VPecQjMT2TRksw0nQjGFY/PT/rO73+eyfaDSANbF5s0t
subFilR+HGTUa02wE3CkRkYXaG+q98JzEVhvLqxcD0mgWsWyx9i1RqBypdi33X7C
N1LoexerY3C3/jvdI+b15wzqyaxH7nylcum98xhpLw3QhR8TD0Yh64mGzJ4ZtVJ8
sp15jIySZ/Lovi+k4X5n3E4IhohTl6IxGqz8JHVFKdQO9MSBiAkuvv5j58aMLMb9
kbKH/RycNOqk29MEyVMcMHBri6mhg8LmZIc211tdnZ2rMWL9B5wStbXc0y3ULo5S
16dZqCf4Sm9SffqrJUUvmebJCo+qmgj88wWaPsOV8nc45AHMUS4A9u7mVPgH3NOj
6r94pp0wSefA2et9P9Q+PmIgys2ozIc9Oeu2tT9uyLRlGmOR7C2NeFMO4GaHhr0f
ovZP+h7m3jh/tP1yOvZ8qeQqdQsVaVk/89YmjNnpXTmrWEOH3R2Sov1ZadUfBQk5
WuvohOr3XQGfvL4HOAqLbJ6atbGWtJdSkXIetk48JC85TJ0CKdjIClDxnh+xy6Xc
7Ow5EYR6gUM1TkqZeqmRNhOwQrQ18CoF/6sEdaPiHWSzj3reunFTqKdSbs/zC7+b
oND8uPHdfv6IS/uQW31+3ayya/9K0mprzFvQIcwBpLgoPhpedWqkJ0ur8IU8GHAW
IIJ/DQ6e9wfui/48F6kRMhf7mw8UhwCm9bsjr4+GVpAvG8h6b/chzToTfE6qyG7i
3BeSpBjnUVLR0D86AG3ENxs21MNjMcKKDfbhDNPGZk/FEJh5oR1LtHDfKo6rKZyr
+r3jcXo9vgiOniNNM3Ut1sHZg4GdEKc0l0LR5YzI9g6sX3zSDy5tBVnub2EfJLf5
6lSAgt1axzRFM4q96V4Vu3WsZWk8nvBS4YebbpChbJhZDahMK26gompV1kGYwlCn
DbNEQQ7sGlWBIKb2zM3uHYvsGLiAgeggW+70FLk2ga6+hswDn0EkkJOmKdzF4zc3
05P1VLJzdJBKnAOS9DB6Pn7tTQXbivifHy8mI0kpgpLTm6x2VRhAa5I2ct7f4iBK
F4D7ZwASNyByuhCabxrCRS0IEdwKaTiMqLS17YwJVmk3W+FbLVRoCffWkaHNLOc7
s4NjN4qNUDvy5fG6UKwa77MYYEDpYrlnfJ2Kd5S2JqsDaAqmuCKC0a7/MKYu6xcr
mZ0Q77stQ7WVU0dLwqhSHmxGOTeslR3Digp+NypL05viFFHYLAG9PxTwH/f1/ddT
ptFCICWJJVkmViuHyGIkxzBvpwH11JjMeWx+kcObaiVEUgZG3d7EIu8nBss/KEdT
mQmRJRkvLemeb5GSpu7017UwxV75gruIAd3Tz/G4Lq7ViOuQgM7b3jI8tDjD9Ros
exf5bkZDnUE34fPP8gFGtj3/COX9I/bCW2jTNlejNx129DmfmJQXbHxxfiPJpup7
PHmnF+hVuDvwjTwdxFO91a14nkf48j9PERnQ+38cO7BMHuaakg4JIFVdLNyuwKom
j4jnL+5V+ffFQD3c9zu+Ibatm2D6yQlIm8fPUHNex9ktBfo4W9TTvQi5GwEdbBTZ
Wg7rVO+RiG0KY/9Dx1J/E8cBMfNBbDa7QJvp9s+s8h6y4oJnsVFVtdBOxI6H8VWL
fb75cwxOVO5ofTxkwahocQBH2AwC8aWbgs0NHzLDiozDhzfhf25FaepDXs8oI6JX
UxcOqN1yla2mvjFIbB9OneOVNXh65eVujTQ06OP0FEYTgruk7hFSaIjxqC0Ne7Ej
IHZVRxv5o7C4nMSK8eV4sdSCYxddfvY2H+JRiW+LkS26jL83VhBxgxyEn6x6A9WH
fcKJaNUcvyGycw+WYeY17M9U7hAQh6sgy3n4esAwlSvGpyYAoAvhen6u9DodI/qX
idsmOu4yvBG9imUuUC8QmUxQrbXTmzxyzj0pabjxZcLU64dNPZqERP6aiBd54dJS
tyGo4CUHBT2wOkU1QCCpJeAr2tmDpaRHwO9j2CM09xqoRMm33vzWswAEwj4NP7xc
g5Oss5bVlu84g6JxnZNEpcfHWlLs50HLjcYfSpkw4SQ2PGL+0y7JZkqZjAdUoQBz
p3L3RfygY/bq9fBZ0wdt4rm/4zyc/L84RzJfGKQRfBTwKF2n2N3Iznen/Ud/rIP/
drJytMg72/LmBu1fMre97CYcrsa35L6hVhk2o2/gRDVyLNsrsPQBZFjfPRU5CiR9
ErFsVE92fEBfL3wHbwv8aEQ6OM+KKWjxM7+P0toq3u6JZ39std1FLzFsGr8/2Fav
a1gAGeh3Xf5V8DS96zka6s0qiO37pbI78So6bu1TliymkDCAeskS3ODD6g2S2JJe
NNFNWgD1u5aXUJyYJXri89vPUMDY13m7taPNJ2bpLihZ3CKsFJVX3MIh7Xn5zRKg
gYUEaJeHK9l2AbpNBKPlTglRzgWei04zUxiGmNAmnuMENz/gi6D+94i6Erv9ecGA
B/wy7ov9+gyDVLnPWUh/XVU1tf57/79L4GdOAtldcS/P+nTqriDHtmuOSsrIMBKF
mi2/1oDRzPFkV3Tqqv7L9tCUtXxYCQHKdpgBSTMJejpTW9aqEMGMob0fZ9f19f9Z
ZvUuPHc3IM8lXaB+u0s4AmdZqt6st7m9/mVpKqg/vWSpN/DnL9YXaeT+XwaaglQ9
KbdWAXWhliYw3MFczHh2rdFXkAimGGscx5P4kDX5As3UCs+6F3htz88e0uQf/Y/Q
OFAzFpv+8inOw/5zGdRWckeB/N5xQ+lwUfpWZ2aKp7dmmDQN2vpJ1DNcTCqTQhua
52VaAUom08A5qWgJrspbatynNJAGKThHDrTcMh6hvN7WYxeoBzqLypheA00a1jDe
XTFONQfGAiaJ86we1Y1OVDoSGjleyRm8WT8OGuldQZ92H/rrhYQ6t2fUDjKhW135
qKD3nX/E0dloj0EsezbzHhS85VA4HLgtxRyEHaMAJ7KE4CxNh6mwyGoc8qlfWYnF
cB1/aCvTdFgorz5/OJIae3YVpOpUst17rbAXZvFD2EUSacibjQNtdkeZx6b9aoov
6SnI8AJi8Ydf2IeBOlEDodrDoVooT0R+XTSZz3FuWSr2Bq519D1EukSoJMpq+W/u
r/PXyISRtiW+MGGcFG7KlUNW44tNf9MjgLw2jZMcnU+KnTCsXFLxQovPknhS4vXK
jy/YdFsrW7Nj+/qIsT7JrOd6XgkVw8WXND8FoWtf7UFLKArSIadA6fX0SpsS5D+W
NNx9mDeR0wYOzod8KkL15IHocs6zNxB62uJ/KojJ8NVKM2m15OA/41VKr0YRBecC
AltPdCj4jVb15fLr7hhuzGPQBVABWIw8Hsk9uf3Oikc+50Xt5vnVaxX2QPHoCO/s
fJxefSuuCclXtRt0BI0BFRcAnSYhD5N5/ievGPJbxK6rhLKirAP+2b1BEbtlw79x
/R4/c1k5VaB4w29hpJXWMtKKcFd22lRdZ1vEgNUKM8oQ9CgwWExM6Gmx0QUX2Hd8
8hP4+sHiE40/cuW65KP5LjULznLOY1isUFSmZFu/SO9wI8aW2fJvQ5FSB1iiJ74K
HxFBiX5MfVC1IbpxVMw43PxxUG4m1i2fhLNtTHKu5ShLIZhWbMw8VlCQFwESq5ay
QsZjX+U9g1E++tpIn0cSVKzAWxe6ESDxuuuo+GmEJ802c7n8LtT5+auZCWeZa9gb
/TWFjPCn3vg5CXYtZBmgdJ2U64ymYxHwTW14gVPOTQCerQLoCr1wC75pBffx/Cb0
kHgISyzkd7ozmMR5blng5AetDa4w3SI0iFXlOQkmQQBTjscDKCE7NOIc/GWKXGwe
CvPBClesQXWFdb+v3Qdv2sycHUUqG/In/OvAKkPI1yiMj9NQPQiUY84QEOtA6/Qx
1lSbEuUIN3UDApjWM1G40b5E1ActAn6jOxmJvAx/B1EPcVp1FdASkEAsDRcxenb3
njqE9W68mo2qP6hsSGXSPSD9lO1lifhAhLTEpPAKQy1HMlX2DaklOR/fXf1VZ+De
AWjCN8mb2SLHxwwAMtnb/2HI4ZnI6W5/tH0wU/BZgA8l58RuCLZh79P/BF/jLOL6
L11xKEieiacKWcparfs5DaTntoVU3NgS0yMnhDKgjYKbqrVTlRZUJ8HvCe9XVFJE
DnmGo5gvwJTC78mm+gZBf6y2bG3V3ATvZbdp43lWaavvQ4Xz64WN2ioCOmrjRO1H
9nzNh12CEqII7XQ0zaNYcjGyX79Id1Y8ThXNrTOYVwjvCOSo4L6dJ/QdK2PD7U6i
78PzE2QYgznCBjDGB9atFHlfANYXhxIek/o3zROjK7Z3v0VMVGUqo3ReLWDf/9zN
saYboPiiEZVVcWgxuhOH1P2Zp3E4GS4IRKvm0rbdYKSJ7UiX49FcNhzpJtlCAK0u
FHjSJ83Ax5Xqc7qoBbOW4Bsyi82grK0gadWpCdIzOyfvHCN3fRRdHIxfZCYd4pdF
g4ru3QSSh17A71lrM5LQ21qB4XoGlKVVHOCfqgz+xfu4I+a2at0RZV1O5ld5w0w7
1A3z5n7OsHkaxpVugiic5lMo6HkEemqCQaDOTeTDPjxwc6P2YJ9cGjL1AoK9O901
azpWQ4I4Uu56v480cV4/I0hgug1bo4Pxf8TE6dI8/iMQP051vO+2KRIHA0Jn5mk2
b4/Tvz+YQig9h6ZQ/jztPG7UOS/VxXsMuyR/FbKK+vn6dc13Yt6qe9gzwQr5KnLY
OJF9nrei5k6m+lLeyezJIFtVGipQvtq9CM9JnSRAS7P9eS0uXW5JEoviRN3rSjqi
mmDi+BaJAHrcccE0W3SbXbFo6yasrb47G6hGZm4nzFShR5CE5aNd12Upzy53KPta
ybs84RbrA0ZVvEgxHIx3uZubUsjiY+C3rzPvP+PRo1CcuRBZnSjNV/br8CHMATXR
cCGAmQD9Vk/L+NpVRqT8aOMr8RefU6lMfTVQZeHbWtpMQPcg1brfjFzGSWA50dff
+lQaSUYxR5/zv4ZE+bjl4cm9WHsVym9htlQYa62soAasZ8kwMTssXgZIhtTIbXl6
bfDz6uv/wGK8sabBpIr5++Mmfb70LaEFscY+uSlpE2ZAlEVeZWevB4Q8+uSeMjVp
CiqKzo2yJlYrgMFDzFaQKrAmNe6rFEZBwvETzcVRWVkkRhmJxL9/9lOyOuebDYm+
Ii0YpPTwMR7Ylla7azbObU6BxtEMiEZPsouTDJRRSLFuVVEsfiFRhoai4XlGacqr
ZZUi+EX5QMR8aTe88YfCrrJfj1kkisy8h41clTq7YOq7yQQlYpRgcpJ2C6iVIXal
3vqfBx4d1mVC4FRwuxXqifygRJefTISqXtn79ZUP8FLYkxHtMA4Ep8izs1VC0s1l
99WTOjIFxN6AZqAnFFjnyonBf/3sLulGv/rqmT3dzynuY6/GCbq0z6aExCOPK7gL
qYkP3lZ5WXsdvrAkCMleLYBroQvbTcciOTZ/e5NYzTBSaDjF5yBOyIcw0/Y8K/85
SMI1O3NM257hi2+/07U6nx/2KHewWQSIP030fHl5KVutoAy/S6q05XfFjePerRkb
ZGdsccLFFtHJUjE+D11704z6qOyOXsgSr9FFMZ9JDWjjNB4jHqH1LMnx2YU8yVJC
0YZ/TRLVb9GJIjruk0dAbW51zYrc6mDVBVQuPjtIOpEKcbOmbsHzpkz+BTyajgUR
+srLtnloyzI6lCkCzRL6pfH+Ubk/5Mvfcl8wrB4wA85Muic8o/fCRZVnL+we4VVV
aSwkTuGiZXebXLqEUQGw9lWQGM5A7dUqwJO8RUrRR9gDbU0+WKGavfdrh8zVlE65
3CTgajfWamU0YfltMZiTDPBNhqgvgyeUH7CDtdZBY853e+yXdijp19EvMAdfgthQ
69uleOymLJaZdTwZu1VEl4c9p3BTunGA3qf3gc5ge1KCrn1tXpdORs9TaK3w1eF8
vQlvUPoNQ38FFPfBXXY+rb2PIINiLP7M1qFfAskfDNKnYUd8ovr507yE//qti8cD
vFm6VcofZzyxA/sBYrjrVve2hzHZQlGNqZCBChXqdfWVvLszrCNkIgeeKSSLAAbr
EMNe09gfe4jTzvcgg0aoJXQ9uVqfD/1opnE+wsD6MHy5Tltv8p+tiaYSsqsTHD24
k2uRJkxaJyGtFDLtTLHKnL8UhdR8TAUarLxaPUgD951vD37UnQTl/d2SmYxLD13F
dx6X5YlKwzry5DG23tsgn8tk+HXBazr5G/rrQWPw+bc8bRmcGzBS0pHqa15v/Ay5
eyAwgqwWwswnl8dIzinoWVqrmZGJCZKC/RUtSWCC8KOujtRgQOV3LvijG6eCUBYq
LR6LEB5zLV48RsQ6RnHlgxDMrJQ0amZvFmb4eHB1OSylDvGyQ06Nh81dQtqhTGm5
nI+r7DbIlmtZOu2QuFfxBqEvCf89pZ7pBIBt3EQUDmCI4RMhz4E4ADNv8BAwE3Be
NHIptAeq1bZkfG86C/bPXHKB2OyvebPeWAnnzX8yorj9kTNflpU91fijEdnqbPgM
bo/n3TLR1hgWWbBFEi4JUVSewWUALUpGWRo6Ad3b5BORbK8mMHYCvI0KQLyRpWF0
b1l1NyoGtQQ6WUX7A78O6N+dvVxSgwoCXarOer/5Fjpd6NWDumv7y+7hQ6kC3Is6
G8omeKAZQ6KfIqHHom+Py5b9KmL12/mVETJoUq52/PpDnBIKJGCYehVXIgEjcaAn
jFQiDoOU9tW6lxezfE7PQt93426XnoSaMi/zWkrI8Pi41sXnVbjovmq/lHVNfr5O
3d52wktGG5NzMBUyKNioHCyF4ESOlF+EEMP/5Y3tzVzOHiA46UOipopicoMtiHvi
ViNBEQlJS175M0ikxTUu3VSkzW0nMeUm0RaGaseUljWmdwoU1OdwFsaSxHmu12+Q
EuJK0HnASFi5qo2ite0mf1vuWS2XWc/F2d3m2jrBPqTV2yphE2kC9OW/WiTcV2TW
f7cUgLE5wFTgU0wGvfWyLQIWUBQSkhQIIt6WjI+KUQl6Dcxnnwi7cSqAgBIvHNzX
xkCdvMZ0KzbAYaTdk0VvUW1303oSUCXFykz2vKLU/C2awdNfeowjpegMezMtBsnc
ta3QaNSXkV1JX6xNliOs17q06RVrQi89U3f05FllGn5vEJa6TZbQ1J7x/yO8CoKs
uUQZwfOAgcFX9xSDhHUZaaSaGCNG/mEhm6g4LCgcAcpQZKcXuRz87YZNKNAfa7Jj
Ew1P1Uw8Un93GoXH4E3FztdvqLz10DYtS2dBJsbXqJi49t8b9LR9ag7QeRW+V9YT
lL5JUvbNRYcrDljvTr1kQsyUain1ZMLHXvnsiRSh3wadx5UfStgrOXg/akaXEjaX
0gYi38GR/4wicxlyaDbf9uo/7Zy0LKoL/8pC2269V1SVq6jGj4rhz1MPRucoO77n
NioZ6lAa64J8n4BAG7OoULUp4zSfFFn8h+CjmhfagsPyAwkbnEyYdzzh4uWgHMdT
r2TD8R0rVoxX1mJ7+VB10BElAo9+gf26yC0QY+9QXm4NeIo7S6HQBR0UbAbTKWti
4+oZXGIG3eZZ3mhlpeX/Zzp9xeKesHTE18ABuXuy5h9igAj1kxW4zM5UOaxzBRMp
2NA5BaVT2PI3yhb5geUSI/iZ85WueLoQEYvQ395QmNNmvuJEHmOo8GR2AeXNCmkQ
Hj7/2TM9ZQ+sXK4ybEuRaeBZ4f2WSmyrrf+lPKSx7BlFJ4Pe+JbmX8gBdmZY2LgV
VT8HkOC6qDEpoOvF+P/nE2Xdx5SSlU1IJGxvdvceMUfyyLI0ZJHNtfsZFeixImWG
/ycI03LXnokbBEUjJSQURYZIGFCcW8QGnXn2gOzSzeSHo6J0nUEGYNIEq/O1qS1e
AUiGLo3xMaffnyRHBYWJ7xg+NOnebO87qAoxsqAidkqyIAXFvkMcTRv3LP7vV6yy
D/gWqIkvb7zm6AP9ydkxQEjmHxI5ffkEL2iQAuWgye1vzFpRpPA+OYH3M2ULsz4t
HArl4qI+ocEHE9V9dlKnIsc5PAxrY+z0Ipw1JyFI4I2VJLRbv0vELAl/mXLBhLH7
EfdvBtHx2bF2xGInVNy65pfFw+OEvmfw2fVaVqcMp68KdfD3e6yaGrU4jNkpvail
Dvmh8K+1VWF3BJjMXbiO5yxsQLMk+OQ29ameQ1G9PAml5cUq2A4935JpQYG7TnIM
GQbEuOlr5qkl+Bu+q20mMhHEB7MGmw72CAzT6m4qWcwkOS0qLlgkqtgLpUKtPuL8
WHgcodkoFjBTxun9IM6XGGN3ab8f0hI+NKD/z49sAdkA9bvPW6o+J0G0VkhRMc1s
AFbx7tlBx0cpWoXpsijQY2nbOnV6U5M48Fyy7eHiqbeAgPclw0ZGv0u6W9FGxNL8
bOg4t9Scv9wRoRAZAFhCLfnKQbRstNk6cLXn/M9xaycDxuYVF3D8OFIUIcBSiylQ
OG1C3d6beckOgDWz/MoA+aY003ed+1pxNRcu8qAmOn3UMkWoH9aa8prH1qMEO/e0
q4bX+H1dKKXei1EvvJKN61l9e1Y4Xa/HI7uj12fGVOGhuOnOi04PaQdg27j/xeXZ
jsUXCgneuP/qs9AZSTruDoDGZaoj7I4GWZtfNcQ7dI/dxz2DpAoHMYVLnsebP2Y+
azInpSu971OMXxhJlryPgmOS4WyCAp+NksdGgjHoDfdXqCelZxbKXlAueXZETpi7
eRC/56g7Z6+oRLhoDJgKWYV4Kj/e+zCPTX+DxTgoodDBmzZ8Y1AATPB352LkVtfH
F4OqcWUEWdQJ3jWiJOzY3cr/DE1I8omfoaMmcyAoZUgwlXubeYRbk6UREhoaUCiR
yeMgIc9LY5qAdpWyVKvc79+2uCBBTwbwWnn0aqY00Eln1JKrJx1beeU4XU7vicbA
agKCznrbczyezzkOjZza0aggaksv2KSC/d9PHMNE9w3cSV2NljROj1QbE1Stb0KZ
VPx9ptsKUmwJY/CFDLN41xjDxfoI15Yb2gErnX9z8Z1N4ZZg0eABgHPEaBrNzVkU
+RSD+0UPy4kEhinamRyHh6OXYrIdzR4scguXMSDpTHMhwzrfFOXCfEkU0wJeHrdj
KklVSZQQzHarWLw4JvKsbRwLZWZPNhvckajsLytjaukPBBrarWau6olrfWjEwkUG
/eqQD5/f5E9eQH/eCbw5Wnzk8lAvoUvDAeUYAp+BlOs9SLXh2uhoxkKk/TCwMCK7
44e2OAI+lIRvsj7oIJawk0mfIJotRQgh+53FVaZ/ms3QuJeUFYF7tp7hJxHkKc6X
jrPWQu1CIoEY/Ftvbv+T3vCkGPd0BlmMB9bh9P95erIZdsQ9MM4QS4V/xBQdQV79
pfeGJAESIwAltM3GBWMhZxsAk4bC1wr0809Afiyt8ZtPPkXrlfN5Oa4C7UPRbGGE
97kMXIgQlq/3ZtlNJ+VMydXdmSdDgHVvW2DRNIpVkJ0kVwFJCP0D52JjEhby/sGc
338Nl4dDDdttB94x0qrWzC8eUMXPryreqF09vKeYGBsbwYXt2DOT/b5ayuJx7R3h
3iSsjzABhqUOs7uErjcRQPj9xBBaAmDp2uXvFbSKA74R/7HbaAvEGznPhzaKGLn4
z+eliA/M+5O4OoB2nE6Tyh9MBHyl4Er7EV2fvlUglr+bcBS1r/Kg+h45NAWqRUcl
SJdhZfKqMbWi5lZuSn3WYGwDcyNRJcQePG91STCtHSWPhQaVjMR6bU8PZIPfQMSr
HFiGJeKtqYO/bjg01llHWrtKk84LOdnwtloDI6o4mWL75V2u7zSkTAUaUe7Dsatu
I5VKICEGOqdcOB9Tk5QGqMPjLG8C+vB70BHUf3wfKmWa95YUFVrLwJFtNqA4im4t
hDRO146LdUd4MuC25eyqL0IU6BbYNtRCSIbVsLBRPffPNMH5dbmyTYgAbTuoVxzn
uqUJcK2ChToDELoGjZEFEPd+cJBvMAcPPjqCm0EDCJZUIeiFcotrNlpBkh1Fdxy/
9SA0Bh2Hm5XKQxnPS2k5zvB/IkTA996z/p5vWV/jduNHErrX18NNh6Uv/rXR+HLq
cr3Z9fMUTMuOFkF33bSv0CUEobH9V4zJtHNy+RCQir696+kF0pLLRLJrTU5yp/WP
z/XMgL/bGGxN0zCwbvzOZU0Z9DLJpfiFvoMX8eezrsY9xdZo7LQ/t+RFY4igL+KG
z0Y9vK6YbZOBNcVRgWEWKwDUqgT8ToZPMoe7cOZnxIZz1g/xAs8yOLP9BX+SKWLL
jka5N0JXL3fcSfW1vmSGM76E6Q2t8ZmSBd9LIQ+XjPfK7epFDOV1Ccs651cLZJ8+
BqDPsXHSR/LQfleq2q2nN+7X2Vkcp82Vsb3ycV4dzGyp+mRAQWCbff86ljbkNQ5k
kE5iE3H3QmFdjbNaZCWziVbgw/W/tMIWJrX4NQQ1P1q/6SsfTWsyGUFszudAOSTU
X9rrGSKMO5VP2ekhphIt8clfJFsGohh37F4P/WDMukXSr8nOJEmn2kAQjxisNt3s
NBxAFaO7o48eL3EYnIK//R0UhkHVoqt7aN1ae9obxQ67qr/cqwd4fTZMoNYLpkSb
pNnTeuGkib+QtBhCEgMhp4zLi4vgO8PGTbQ8X4y/bKZn0lZAeB9CEwfCv4Mt2dIM
Scr9pimGlwd+XTiM931DnWdgqSeJz+RKHYOZkWvZsIACYWFmTFRCSDFGKOToYxoF
mJuRpkOahBizEiTflXX+e78HvOzG2+s2PfRSDUzu+gcDqcKxi1f+oSHf9KiQnkK6
1BxsESVJR9x7xYGeaGSJ6PXRleDgohPKlqa2AKohqb0UjjdGjGiq+w+/rQQb16N3
bq2jMu59Wq2tFCYMEqv40pWYXRFGxx5KyVWCpoB/6eQyRiohpb1LcZOQL0Oect7L
ohurmSWM9lg6Bz9t/FQv32Te5sRqY/CxIVF7ZnlgrEKczh1ndgGNT0CdEPuGPjpc
TR3j4XVogNJdIZx7CoplDj45fg2A1WTsxZBFQ3rkIdWLljM48xL5tBzHezb7STx5
xdRpDoX3TfCHE8jOtq60+cS2r7h1FXz5gy28OAJl/VJRX0YQKSMcqK4eqA4FZEkT
Mi6nyzFi1QdZTXph965tnIPm3LY8VYS1BKmwlKDjCTbFkXz/rM8NUkagxBo8W7u1
graLRjdlnRNpy4pgM3SSmVbR8E20sv4/uJUUssL4vkFR0Dz/6BgUO48D2i/iviyK
0b/mQnLAAexSMy+BZ6gVcXbbmEwCCK4sehptVTnG9bLZTiPpMWyehfaIRa+UNLFe
rgyWYpcptkVdWGVXpgI5vX3zH3SGwsFkvA8JFOBBNRc5e6P/GwgUAxTYb7cU/BT1
ttzdYKsllriFVND15qYyAE4of5ov9zbhGxx5oqsDn2Q+BCSHscaDNSdZ8D0KMXHF
OVdCiwVbuDtNYeQlv5OS9nwtTc95Rr+j+IXZR8uf99GxwxJjjiXapFNZunzL68Hv
V8gQZXaV/rCXCcHFff3sWj3u1PSirGOJahjUO0lQGe9Qb4boiqmEfjAAyw9Ogd6h
Ynm+YysstsbYyUfKhJ5AdRR8ZArAeCZSgW3niWq8bQNSdVaRAKTeu+u/+4Ox14L3
e3eWiW89xL1WExP+iiwtdzQPk8p1kd+uN098jDfcAVB+IBOdIeSfymXaGXgJwdD4
rw3ZP5VTcs84D4xFWSgs3VfLR1UD4idnF+ZG5lihQAfBwmaYy9G53j/aVzZSNl8K
4qIhp6HAmue6fYx/AtcM4MIXHVA+H9M+dy8Iwwi9mkMj8WdY6MCCxWrw1ctYZei7
14uBcOw2ayPJw75OixqlvgV5Ek9kkTfy7FN39Wv+c/HSJjSCqU2Bb0ykdug49YSH
sflCpksq2wsl2HkgU0nvNLfvsuIgw4yt7UM1SXH3+aSxF6Q87fJIS5lMmaU6nBmN
BJ0QEtYobFAkRGp3XNd65wTmZljtoZNY2h9WMHzxAlG8CStsURRnJfLt5XuoHNBD
+NjiJyie1M3cWvFBt7dLF0/TMTW50hHFumh20O4D6V4waMGFJzAeUrQFrkOi2D7S
ravOIo6Ygb2qlQkWVpQfeQtZ0Dr6aP+UWzmf3LvRDIaKYh4KbT7YLzklxuVyBnNW
efT/dxW9FkvfD9ZV7M/vlLTnzlJ1fudDvU5NZzEq77PQDn9k59EWdxUqy2bsL10n
5X8wieRMPa7MMTrunNB/LweYd+2t5YAyrQpWVJSxuOuwv3AA+eW+QbJwLdCb24oN
dk+FJBYdm5Pn//PHNox2Otfn/q1musqYxzngVqJvygQErFNt88d5OCsZDXtgtVAC
h4P05vTZdK4GeOjJM7PNnFl6jRFi4ev7ubzxRBPyEz1kQouSZZu0tVs/8AUfsThK
vygqjHiyZsxPZyP0RgDqDPP0QVAZFAdeydcF/0yHnLqf/3s/ZSdWmyTuHlw3edIh
sMQhadH321dct+kgWxXlUcJkHDQIEDG4RkCv5SsmIKCsk1OlZrM+Fun8ipIMa4xL
sS7oSDPEwN8w871+au4RPKwQE7m9Mwrtdd0NR2N5CsymLh0QUovnuvU+fc2bBMRA
LXsjyWdMFLS1eV1EFygfNelWNIRHQmYLrgQKQfAQ78SHZ2yTROtR3fta8ZDRjx/0
xPpjaviuG1gCTqbLAK/1BkS8ub82Ww4x6UDV+XYu+pbYuaty2M2ye9fVoSebRCDd
/PlOHXS9ZNyhmZoJgaV5sAgNN+UTivXRb4Uiko5HgXIsZwuwTQ7mMJSJv74Sti23
6ptFF8tcznQTqPlVCkMRLzKjItrMCpU2Y5XzrOmltauEjsVVRxY4JWZudhUl4qdR
vC3tch5QUFVC/3kq8TM1z+kfiIxDrk+fZLmUOrfj0bbY8H/fzhpY74RWfhTd10rD
QSELoR022zMbM9JQSdYAxxFHmBjcS9pzdnRjdonMJSKdJvffnUdJyp+oMgHBNlR4
I69Im/wjQEUxCCLAfpSClgTdH0vMbG7cR4Serkm2RJEz05FxlfzPsFpP8g92gjFA
pm/qvWpfTQbTixUY0l0LVBVBC0a0GOPxGGtnVLA+m8fMVf3bCDLy5hpXpqoqqs4U
e33GY56KkprEBmYGO6MM1rCUyKRTnLaPBfD4t8BtH17V7Gu7ha7kWH6ugTc3lsKw
E8HWA5g/qucPQOUfDBIqZZN8tc5VkibaTmTzc/XThPZwZRqG2xhOj1of8xfAPaEg
4yEYU2SlyaTjI1ZN3nVFxw8pN9xiF+AmP3S9YeurLHnCjyGwmVVKrxDQTQLTvp7n
JzfN0Tz2QTAzPhv+Dkpz2/qO0I7HK4Zhcb3blPU1WGot1sabs1E7jMlTkNp+mpbx
3lhqKkG/J6AcHU/58TNtQtBDCqBLMsWJT0BjwjojIBhHUPgBVuyqZXOuleDWjbOx
5b1gUctmj+nlqJCeymAhQ81R1TfZ3dWE794hHAI6DRPG6N3WjRAD54mxO1eg4SSK
5Gf1Q0PQnSmhv/hHyNXj2VTSBp/vDcbNs0mCblK3hNjWVnkRS6IMDgwKF+w9nzFq
+N28GRqtEh4vSHon31glaIzOlw/Z5cNuXEjJrcxM6QvBBvR+jwbM9GlV6d0Jdc4n
XFwKDvbYsy7cLtrZ/ylPzy3Tmd555wZJGAMXcHzR3iTmX71F2LXa27gOKeVxUKob
hZrMhxVY86ZbUP37dg/OgklLAJWvQhSn44Fh2jMO0YsRnlzeJOV5o/eCSR+6byVN
K65YWBS8NrXXEc5+L0FXPaolG7vQkL6KGCAQqz8C6E88jzP/fvTfTesisytipJZa
uahskHhSDnMU7RFOyIKhB1ucok7o3uEXR+X8MfGkxNXpuaa7b+Y3AeW08/uhIiV1
vDMT6Flzs0QtYs0f4gUDnoyOXnpB2p+GS6VpCdc2OdjmoQklkFc9aMXRS3VkBZ2w
UipplaEMsAwL0l/f4GtUx9WsxESnFybMrb2D9GFJbC8hKQhX6U5Yx3fmwoZAaUTu
0JJSGqaxhJZEViewq9OStyjPEBuYgGNM+ZK/HI0tyylxDlJTaXVV/cP/nztfmPeX
CgRmgP7AOXuurrlZWZhPqJiXY1mKmrgroGrPCf7tfGxewiT/+pSgig5B91o542Lb
UAyAK8ZUdL+RbpGzH04jOYW5ZL4cE78FsrcsXpUyZ0VNdKWzW6TM155c0QaypTQs
eVQoKG+lthNkiJ/Zjgfb2uYPFiVhqGRe47oTeTc5wpZU1awrjOTWPa4z05Gv2Eta
uFPLu9Q210XXWfdm6OCPUJ2kZubXWbcQmUjNKA7aENuhS3Y7tdIiiTYnY+/gQCHv
3XmE6Y0oUdpLtNWY9y2xYpx0rPTnsY+//5LlxdJ695EXd/lbP2mVVzQ3vi35Bi9Z
3Gj6BRJpP6SKuBKnwCWxHWn441R7vBSl5MTuluvyZBtikmFyaAvLb7SGF4ZfZi49
QSAZVl2rSRUwSN3vfo/2fsYEad1UJJcfc00swt+u0ATZIk5he+Ftu9R8DlNlVRRm
3+40PQDHwPt5Ug8KGGvOqFGaLvYIu73qEZRIXqemAo3bviqHA9wGy+mZ9FKPelOA
BcqocHS6K1cULVw39cgQwvI370MndYy28yrcBYz4n8wwS97ObI1GZ2qCQHnUJqcH
i/t6o8GTSO3K7/oup6d3gu4O/zwpzi/C6pnCG0nGSpTXVVjt7bdOJ0ROHtdtAc0r
U/7LIqafLkJHM6g8PSLpKhYeqsirqvIZ10BbnWfhQHLPSpzRLSOQnmPV60SQp3Z0
bfOjLoHpWjQeRKk94xOfZfLVT9VGO35aIdJtsmiMjO+qZ0YLqDofIG1wTu+Fewfc
LDgngjwLxl9kCC9RDQ809hnH7S0vOa2UIAz2CgHdqcC9NHclBQ203lI3T7qbBASa
qIz4AMQXZIehuTVI2Qy6DjbsD6sfsZNAOKWIBChzRSYXMWC/pluIAoM+O5s3+AVS
crdOAtmvsebgCe3VahGDWNM9mzIrT7M4MAE81a/E7UllnEBZx6BZzW9VUXfpV3Z8
PbVYiDJzZro6BfgH3IEoPkgKQkPlFcKeorzS7n69z7DQt2+fd3AEsk7JbxJRidrs
H/3An5Rcyo0ZnNDiJYzcqzYkrK95qIsvZV4WooKw2dkMpS/yofAiGcVvO03vhNU8
ssNKdeYJL5aVhlKEdGlkAPl5jnv4Pn4ZSnHQAqXuBArwbMHJMzAJElvq/T23ot1v
VEA4dlv/Uk+JqvpgmvqQUGAyQ/NJdX+IhR0kXiPSyrSwnK74EsSxjmySUdOC3kEu
eSS6O/RVz0d5J64z5mTGPzfsIBVDNFrvaYd6qG3zvfEWyOAi5l5slDSRbRUpFxA8
kt9Cp5gSpU3JtNG5w2yxxjgJrS9Vw+fqZv+M/2KjxlpfU4myn1qz3q5ujwBJsQFj
zk6J6JpvAQkQdPkKkM1okQGH91FZHyujkflYkyOpBeH+zox2pdvmXmaiDE70E36h
bpsVXqjPDKgmyywMnF13oq/W1TcMwGmtpEIbKEYvG32V2Mn/9d9dAulbwR3f5DQL
a/AZIISrBMVLTw6M7XFzQ6KUTzLSz8CX8YzLcbf2azDkKQGTkyPu7e3kEnDq+fov
NCrdb5aQmZkN3VnauwpGI2OO76xExpTliBRT6nrgWdDWIllo+oL9D5M/7zqS4MNs
f0hrrqPEFh15c2evMH0RfUOpEG4epRNDGUGMT/I6uvsTFEWQWub/xsNn1JwNmiRW
e3ASVgRhtKl/MXTWxl2+oLxfz+TDXy3dJLAvu1yFWwKz//i0s19mjteknBkTfNWJ
lbe7VVAvf4AXOU9QopKzqp3e0VhKaIwH0GPH6hewB6SytKJr6pwKHZXQpD0knY/W
st5F7NXzhBUWzNJa1EWO+hgsNgqqlsLy6wsZ7bOzDzbFZKQ8IoJ4APhH2KTvPL24
+klgGvK8+VR0vO37zMOChQxbYYwG7NGdT/B3dimx5o6wvwDo6syQn0rexZPFdG4z
789xrK+FqQwuiPyOE53zK1p5LE/F15IXbm9K+egEAtWlYSBRXotNEzjfFwA46Tbq
T0kooWcCGTq4fPYm6E8Z4xCUITU+4Pmcz+efCfrS3xIgkfHM+a7Wy4CgxIl8mkXB
zEgKNZfG6UN2CDSG73Oz4Bn1QNaiWFTzFaYyNfju5QoTyXVE2IoRqzNrM0Q4ZlDS
Yds20nCWBqS0bJf2k1eqDIjluQNM1S2WIoxfUI8vlX9Jt4YG6USyIn427nclFzP3
0TXMEhnjyQIfVSp49K1hl965rxj6u5yVuL2+xA/SZa8xQQH8ocW+UZlDOnI7T2Ea
YG2l54cB8tKhmp4OZcvtqmFzcvDBcyvuFAAfSZTKgaWszzjjUstPzcgwVhU7TfHj
dHkttxckXCf45FeTxPCOItyV0Q8TE5WGbC0wV3AjZhi381wKQGjHzviFkJjY4nhJ
Z/tONTBMFV92tqtv8gV3scAHGwnXLxlVLkjPpRwjIKPZCHoFmaxwkvostpcnwbSR
r5TspRWgikBzxOEqcOHdUqy5THJLXqXtVvKIhEB0EhWt1sCTMCHVA5BrYTO5QFcQ
ZbEwiU6Yo+3uOzlDjTpeNtYZF13ICJqA22vnrh3GGmGDKySSlIGdhpyZWwaiiOXX
4w6rjpt72FPkH+t/NiNoA1hY7cxEt+EAwuY4coVqHTYZ2kbh0j1z4mnvisLtniCn
dzkmumtxgpcdyGSwjz8cVgPg6VxugOEk1ICFlEgXKDZjZv3Fa3VN50oCJI43mJhi
3PjwWwDGqdmj+reutjJFglYUsf++HoatXJw4Xbxk9zT8NIJDzqVNJxdnFUsykJL+
ufVaTUifaFhJgF9H4ezhCgngNe7NQqc2v5GYJ37vno26RlP+Y3cPPitlwgtQvN5Q
28r466buSo6BfZlEPWBLba5WSezW6wfTNB/WvavfhGqn2zYG029DF29SCEzjP3dr
KbJE7QD7J1kmxFcdvjft1m5ilQPFjyKYg/GIMG7s0gWBoQSoPVpdDbgQI9GJIe9u
8A8hhroPuiJZpjinLY5it8UxAsEoX8d/o1+LjAG6jyU49AVnCzichJbzsflDd0Od
xRCVaCL+J6TmmtmwszVzW8zDwBIXLPAFPVAGUjt58i2b+Wgr0ZjpYHzrfQ9uVACI
lSw9EtXpdyYedtc6q7W6NaATGiYai2iz6ps3nh80JapHAzcdf2Yy7x49lPRc1xVD
UY2uGxOpZSPShndCHo+yXa5OrCOYfyDjgm9mX+jdx9rPhWxJKONVCneQbc1Q5h6H
p9nrSiSt7cS8+4ru3c53ihBs1yPucT61kcDud3m5OcSqDoBxRGuDfAa3dAinbbN/
N5KX36HDwcwO/8O6onq9ms07DxCOx1q3l/QhmwwNuC6F/bKBgdF4KJL9oxBt2miG
hOeDFVSCDtQ7NOyLyharcu+/5Y+RSSdVDIhRkhIwfTvZFvhiQGZOX+/qwkwHbIn0
zXk3vyinyf228kOzk2BIFr52x4CS4rlAQZBXC3/hzDFov4+M2fQkPzDrQjMFnPHs
Gdn0qKJV9iju4pTuJZJMoy1J11fuKJU7k9D+7T+xHxQQrKZEzkp1H+eo9EV2gwhX
8XkfQh+WNhnyy8uxRD7zMXeURXmBvcTXyatbBSuuBQGp6Jkkp3ZIIdz3tNm/o8ax
QYhnYYWpCasvhkuZ8SKzEcXaLP7TVoW26Q4nv/IKKzHeBWqZOyXZxFCYvUxvsq1Y
1pUcBJMBlXRilO3dRehHOvQBDhSuP9Nf0jaVZxi53IR4PkEpgPnIsiJwr5TV1Qo9
sVVPoa7lom9rjtiMkkVViehrMpijeEd3fYqqUDSIFjXvJGYPDeofj4EL1Gd2zDmy
IBcR2l3/oFvkjtuqCXuH93dtKPK0ASE74MoONIIXWnGiOc2vKFtpGh7fd66fWRfT
UEjh1/5ur1rTc7gxGUnvL1zGsbUvo0uemZerRIZkw0b3vOmWHoNo9gQATv5uzirK
l/MwK2+VZwwaO0FW3FODHzyqFMjNRtuGt4bsQka25rUrZanqRjtNVSzcP0jZzrrZ
1SDn3T4MBXigsxM+qlYMNGvrVnk9RZdAjoN8qzMy6n2Eo+I82f5Mz8h29KnHMjs0
3uscekS116clqZAKyRAip4TolmReKyI+vYyxFt/V0BRcPJWFECFYSGCrl/LmDlWb
1iPRbWi3F1VEuri901VF9ZuO5QDb5gbPVjvQ3BZER0cTGt64dLndPXjO/kJBssR3
ak3dJ3is5NgPXifKR7ucpwvjjxRC/gh65AHRTvf2G750sbyYHUPPFnOP2exOYHUA
5b0t98eU6yAQVQMEpyHq+N8oiPpFTwatNjVH+v906QfAnwhRDLm3PCetAU5sA9P8
e7EpnxEEJZJgd1pXiEQHv9yoZGkw1XKdi/fDc+VsDYkH2osrFu9WqbA6s16lgBsI
M35rv65po7h7PkDReaBzdZVDkHw6aMbBJ6fJIu+AWCTLTOYjXzjCzX8Jb4TwEKOB
MdhphJzw+NyJMAA+WxJ+03ElpzTPqRcaBX+EoIDGd4cpHt1fz1iJETIp5v6I5HKI
9guTeRVtaZXXxscOznZ7x0uoN4I+/bKuD5pIlmUiR1aH5D+pf3EaEz8dYzAEUPs7
yQGm3ya2Yi6rOIJ/meMM+rvjIfzWcquIMvJZmWVhmwIt//UmvEbH3FiX4lxQyP1b
wMcU3iDqQsPXwpMt12ErulErsnNR1canbz1iUu4Agf4l2I3kx8NcAte8wrtdJttg
DLeAf61QVcK1NXaZeUQksGZiK46n+Y/gjXmov+yg06nxaueGZA8xeyKBP6qvDedV
gSzUv6HsHBMVSf2EHnQH767UgcGNLhFhreomB4vferjI5Db4uHnfcBDj1mrL5TcJ
4J8V97NtgBjNF8z2uoT4pqtNo1umtzPWJGkmjSVflgrlsJ6hx27y2fYjPldKdl7g
FWmf7eA5NYqUTt3abp0+Hqb2J6myRQcpIYEOTVl0+OevCFyMUAOfRMHtrnALTNGB
yU2xhiOyUcyg60kLKp+gWPeG1+QBeerG6or4ZHfKHEo3hONxWWOWU8jeL98if35H
MCmneJkH0cK7/GbXob32VR4mrAjdX/IRqxLTv43pzG1LiZxivK7Xt/ib9AnP0e58
q5yMPTj+e12WkvInuc4HhW/5qR0QcdXp5hOjZFv3zvggLIK3p5UvhRaLXlx+WqKU
juKMycWyGujtKh7wD5ZjsF5Y37Z6T/LILfNj2DLNIXBK35vsLGU0v+HMIw6wALUe
PbU9/CuJZnrDxXjk1FeVRTFZEMCnL/W2fpZSSHHi0OIwyd3gwTf2e3xrnLC07o04
C7SFlVxfa4AnroKKUxUGzwHo9u7wO3Lwjc5y6ke9PuX7PbConwt+WzRP4isPbN2B
pTbofmt0WwF2a+YkUKvKxD5VRSuCHyMl8bJOtyqfb7S7GAa8l+1F1qKsAf8tDTMN
ZnIR5FFkfNygo28M0oiWQMryiCgxlbP5qU8sMR9PD8lyZ0w2HyWuV1fPWBOdEZcb
EqewjniHjjFO1EDymufsbhBgqGWme2vF19wAdhTkYJQ1VuT1TBDL0fCfKnpSENmL
GHD18FwWmeppl0FTckX2IgQafVuvUn6FjYztKpkQandcrMlysOtR5B6XBTiDrEME
3Ty5lYNLPoqFGdy0+/XJih0RkII+JlUBPPRBrp+exwqDwhbyGEEugs+vO1gwBDxT
idisMyYKMQoTjPV7Crfooc3W5A+v36OhEMu7obNz8aC3G9/TC/8HW1BI79e2uqSn
DFibnmAj0M9xva8V1uAoNLnxKZgYiMeAasD9CEARNim1w2yAaVwIHLmsGaaNKnTX
15sSgjvwZcHHx3e2v0PO/Acg28Q63JjLRVTzXZyTUKSkG9SJhG1/EzKRXzviBzeA
1+4Yem8nzpIt/0GwGcqkzmpRtBs7Fh8rIDOs3cW+7hZ5iYykaRq70ll+JE7waM5t
cmYYBt6WJrazg1E5IYAzzX4Fq1ESHW1NAzgCV6TaUqGej5QliXpU6/EV2Uh//aPa
1ydbtsAxru4ZsrxyQSYu8fySDq/jrUkzlaSXWFVdOBHMfmBNT7SgQ7Q2Z86nO89I
xx+dyHw171g5EmAVXdWrzO95BoKPA5C+5m+ndzKiDHfBkAZeTFp4baBHXj0/nUlt
T9N5+AQ4uZ+faL262WeN+6RT241Izym8Lh2hyZ3u1gTAXPreOxGYSaFDtwSCi3KT
K3SgtBaxlFHEbvw9WIAXRJqiP0DtveybjaJIgNa7NmdzQ3vr3pMtnPuDaZuBhKxf
RGD9bkezSR7eDH79+k1F2aH63W8Jy2UQ+L49BQptitlgoPvhu/UQ3eVE6oUKepEo
Tt7VIsBjVhGIcR3BypE5lrU3nPD072phJUP2gpJOaCSmBj1owlkKmjY1FjFCP2Dz
7RgRjy7FLhJ4VUfOqmaV8iGZRfzF1DJ+TfaRmyBT5K2HE1pBJPO4k7gVgrXFGZBn
5wU0m54BEwKgTwh7KoEzM28yw1MZ55ZVuqdD/FaxNPDiNp75JPecO55Pn2yGVvzy
A2F0IXZPLVLfbH7hagtEiDBIP4/kDUgLMQujGyk4V+BNBSpZqs2I5l8sps+YV9vN
sMxZ+06hFXAmSgxdrGiRAPq+Z1/JaT0s5JYNCSqMbwLJnNxEGwJXr85i3MUkH1Fq
WLOeu2nowQx0diUteabV+gpHxYhbPbkKBy0JKP+E/Uz7fDC9BuAJgJZAQoeB3bzg
J+xTVpRy9APiaTnYFkXisOE3lld9aJ9Mvwwoab6B9oyvJlWIk2FZq5vKjXRLOZVX
LYDVdnjwC50/2S/7uXtEsQy8dkBrK/xesSyKFaRCO8wvXFgTkIvH66yyOBbyDU6M
kLNbz5+AzYSpsOIuAy/AR8XsHyNg82sSF2RaQs8Qu71fIF2pspighXtCNT2I2Ih3
mAn559FDI4pjYKpocnDEFo/npIJneA0EF02xNnnXAiaay+TWWr+5EuIf2tfRfa7+
kzr63rlaFlQFZPGoNdSx/m0l3jkIbCaaf5TF8l8dJ3g0wctIWL/Aj4txLU6NumoT
J/9BY2XjZ5KSpAIEtMkjILkOd/O4aDOvMACRFFUOfc+gsdF+oTt8ZqTub6QQP0Ls
nNENinrVS0RAB/N5RR5p5foYqJXG14GScPADZ563e/O79IwOiHDmryX6hhvR+WQI
6/0uLJd4/rizygPujsOIXTDvzs0VyXYuVBVK8xPWEKLFwT6gSrrLDuzcyd6JuuIj
Nn7Nzko9llymVU7bU12mRtnF9/I0/O/tnNUnB70auMpNO6pKDy/OZ968/MdLfO9l
NY7V+MP8iDKzWgy5cX/6kvQqyvA0NJHjJUPVm8tJ4BEdfPP15mN9Lm2Wb3JqgdgS
1g7HIfmpGOO9S8Y0vJQClQ4DkLT2kE3Z8UyZufzgzcrkXJOJ2rDQFrgl7v31LRJe
Hc1PdTxYD6VPZipbIlqNAyWCKH9Mw+Q/WuRAWJnEvaJhXKQ9hLzyP0Su0UnBE9Aq
xf8TrXtbAj/4PKPBNXCIA5KCs6wa5PT1Xnmv9/uUniKp7Z74XgLu9zyXuKYPEzzt
ZNeUPeslKXY1Q/e9rjM3I88Ae0tWn4H0X2zylDHfYFaRs0UFnrXT4TidH713JjSF
chu/q0NReN64ToN1nzfQowWuBezNOGTkvOwJzNKIcX3QvN+ofbwBM7xn7B6KAHoZ
raBCZc+GWomHB08R8j1/QVr4cFkjKJef19WShx2jdpTgb/VjNphx6w1vYJTLAbC5
AgjTGRhPwOkLT4FywnlSvc+fR8uRrovKKZUnGWj3JQNfRgFqRdXt2hS2KGIroWNR
itquPECm7ZbbcmQHvxLhHK9Vnv+5Zi1/7YOSnUAPRiffwmWLLmwh4xBGIxDzGvE1
pi8K9aQRNTAxiN1YwDgSVjPQioFk9GR1sQooSR2XSak41SfXJVnjg9Uhkr0v2zQa
uwPVmZ8gWNbprEgPvaTXX5lK5RmX2q271Pn04IQVM5A0u3ic8ifyeuS5/S9LsimN
MQzKmTHZHvPEK5uubKd8ckuEDfncZBAOB0rO4h4386VgNoRuC03P1qYNr9ShHY07
TnDnBD9deebJAAIeg38vnup54lN9aVJKe2wx0kGkgZDqBb+K62KuneJlpQSouzod
548JFfKuY/pX743B+gF6e/O05vulf8romF7toWVmBH0mGwcsv7RfhwiroYoUfZjg
ENZVXN2mPgdGLYiHhmVUVfwqpwCq4q9SOpzTnn6Avssc+m09vInN+EiS1s496lcD
Ikr3qRB22qoBhEmbFf6cAp4LpsaoRPhkipp6abGOSF4GuM2wMRNai2OIFVRDUA+Q
an1JNp10ONLTXwLWmQcQ909jrykuGkbXOnA/5GgF6MoLi9PaaY3KfJINLsXW2zea
E/ZXVqWqVK6MNQNd8dLBUvZzldZKPmrct+D2aKe6wsraeHwsoOYIyP4Jg6vL1Cis
P/uxTbw7JRFk9BNeqFS5h7x7Y7uMkoLk8XKiINHnl9ztGyVzcAuKUeWn0eF0pfqF
SEVq2lpj0PJkR0aM0hxRf454ZOzm+P+sljgzFbiN4xIVLICLWYvSzhcXryZzWkPv
sQQky6+fSV8TuOULlHemVqMZxsQmeXPb25giZukhKND4VKpXi1Q+gNgOxI7b2ev2
4xepvBxDvG77hw6G1ceiKu8zzQUoq7U1rfZ6d+LhHQc3iI/7oy2MuVnJnRLKtOMf
t/xbsJB/n2mc6b9HvN+dh67gLXpiEQSymQRhy3QQ89j+FUXq+3ZlodFHY2MBVlnc
fzfQziJ+WoYleUqfpHqhWJflaOimJZOrWDviUBos5nzk9fCcXk1pBLaGLS119xJi
7zXHvj9kjeADYfg0iCQIrOesdH4zaXn6ClWTNRsZBxEwmmnL1nUeXi3KlOklQPz+
P3Fh5jxZ2HHzGGfw0tbjmjm5rmn2EkdK5B6J4gI96+oxf6DHNsU51yUOEdCZMQmQ
3VQ5fvYC/3sAwoUHzbrgLGvFbMHfu0iM8PgCCCx+9czGK3L9VZKNfxHPMCPkEOLe
MIEJriBUgX0fDBCMJ2sRcz2GjMu/9AwM/Q9Dnub6OQR38SYoNPNIXxdOyjq/smKO
EBM02EvH+cRhmv78QxQHPsY3qEUn3eq9VcaSVIBKU2d4w4i7OEAdYFN0Wuwj9LDX
ACMBG1kF2lML1aKTdsfAaKgRERmAj1CndPFIwpVtN08mY7tlgdpl/+huLD60NEpv
U7BpceW3e6aB4ijbwJpxNgfFlN/IMU1VofmugDEVd1Cc33KAXUU9uGj8tQendynf
1f+5eD17QQSj2+/iADC2YcJyYCFRZ1DbO0wKAuvn9+Y=
`pragma protect end_protected
