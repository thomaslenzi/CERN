// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SxNbLZFw+/AsiJQp21/tcNjkbtGvPSrqRjWG520FhXxot+98UyCVUmt3JPns0DGv
ctbg8YfPiIf9tmqgKsmc9JW5LJnkMqTrtahH43N04I/5B8G3sT523HF0F+MHQ3IC
xWizcZLaqsH1Ic3mrPexDjcd5nlqef46d0o1eXDkqbs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13776)
fV6+MbTuRHYKuM2p6An0cChr/50YrYjWjBQvZGPWzNiH0dNFKdkWeBdRCRc5t9aI
EW3LxnuHfoI0T1Ak+atZzWFjWPaZjNqpBHQwrzl7uVSD27Z3D5oRJ8Pm+NFJSAg0
jPFefZWkmvjvta/NMIEqP8A0WxgoHFxUrww7Gix5mpjBjH6G/Kt8Ebo+EMmDUtOq
blDQjDrvd3mWrIaXsf2bGqTi3YLIHZyktCYnPPwgUNqj3+9qWfb9PLAIczViXljg
2fvl2R+ki09vNa9BmifKvDXMXNvTCz9JuaHS2xqAllu3cvA16RF7CrGDhtd4bvJ9
MsedA7UN1d7JTbcjpZiqNHXfcUVcprlnB9/C8k8YiOIga9rb0Imn1gZ7JweV7GYC
Vy+YqMHme0A11shIycTUCVfHg8yG1SWq7ItZQSJvz92cmqEsFZVyS+/9I3RTm7cj
0xdNG/hUS0n5XHfDUjp4fLdIbYyT+/cfirmPmdtX3FWxQTJPFDJYqo5owt1ax7n+
gIrFhfaHWLPFHh0FezHl15Wrz+RIVFkFpQFHKICtXRm57es2L0cxbFrhrXkygQuf
cgkNliBozy5j6BCN7e83PKNeDjSY7GZHUCe9UHVyKrV7rHFdkp4nQXxl+4nA5H/3
eNSqVZvWp8d0XemOh3TbXg13HB6XLhO7owrJjflB8rgtMntpgju3bA61rxImzfRy
O6NTRmGjzfHZnkCA4VRcgyjAWagbZMSjpMsKiEc7Ao+LN5iWnG8DX/YxcEPoJNNV
aZga3L3szCZzf1eEFdtXDoqPrayeLWyWmVPD6A61f2prNYs8nCdjGZYXNLO2Yc3A
/g3Go3YoOmzw4X9gehv9JQIG+h33eKMTsyK8tjOIGQnsXNSyk6atRoSqxae4GgJ0
rpJxm88dU1XFuO85Bv57PJHvSL06j32w+Aa1lu5xwa7L3sN3pIb0W5Pza3fMcoIJ
MgLHMHRI27HC9JAUSwf2EovCF5QoESNjSs+R2JwT3+IztkQxRyfu0xwiOWs1Le0q
Z/FE6QWu+Shmby7AcWnOAaqbZ8yO5TI3+VPYecUeFgL7GOKioRTKotrDM18MWSWC
9PGQCveZUYcewsK30oAUB1+bxWdOrF1OljkcbFk24a7YMWUSi1wvongB5b2kZL4N
odTa5lM7HBGq3lYzbnzb4yj5FoJ1OEmyVl25fVym1w5AgvlI9f4AEAI7atGIanPD
tAYBmY3bN1G7Ox+ZmAGtq8ZOL2jJKhbSpZKNS6jHXp+viGvl72Kk11oZQLMkd5JU
aiqTAOITZlZHIhzKZt38Huwc7p1YdmHtnowJoIPnWD0kVQf9oCeBxcA/HDh915yU
MHuOUEiwmJ2KEFGYlg0X9R5jjKiaWXCAJoIiivTEmHQdsYQXdMaSdmbjizzZ6GBl
ev4eN3R3aXA2UYL4SUmWBnWsjZfT4sZxT4JUwMsFrJYH3WKtBS7Ocn7lH0UvIhoe
V/HXT48+7t4npVlsrYjtbme55O+7kSrKrnf7E5heDKCJKLJurtQA2dIfitznVhak
wZNdk55ZHvUJuNFJjRcY1q3KcL+5M3rc40ZwonzIocYigsZAFGsE5PkN56EmiuMx
L/SJky+E9uwL66Tcl7pvCQ9bRsjdzEhozftPakUseFiGfZZ9uMehEJ/Ee5SO6ob6
RGFBNQph2GW+GslG5W3HvwDdX1lpqyGuKYi0QG6I6yvEidrHCGZ2iBSuW5GuQr/m
w9ALy7StoGTSyyHj2rGUXI9VMPZahkXttScE1+sNvevdG8oe95rpr6GX7ThlFWiM
ABAj85js8oSYr4b/TSVw/MweC39uEgPFw7aZLTFeI0V+ybJYRATgo06tpZbHZdHU
7OtO+NG083YX1yF2Y3ZZTyuBo1tFstug7IRPlB4fjHCdsasAKRYPRGMUMTq84LeW
DEIqKnlEWxdiWt9GuqZHLGGAmtOGZOZmpNOQTdi+yxHQsgUwxStMZMVpitlFiz3V
AHxb0wY4Egg5c4QdBmyH9KOkiDL50s+LiZvxTOjX26zqOwUB06V6HA0uDBvSwHOv
hBVX9ANdz+85EDKexqjxTvroGksqkV9ut11CBdrQRIpPqz5QhwF2LcZAkEJmCg+n
lC/M6sLDNDkSktLo1goNiz34pT7SG9+RBuZH0SY1V3AbeM3Ol4/pwvnd4WrsmqXd
QVw/r4bx4F/VvgZs2StMV6puWUD+OwttVGhd/GWOIZPoIXY9LEXcHZbDW0Pi+TJc
8562OwGThDNtq3M4jgwrzSH3iMn214xFSIJNiax3AdHWtxB5htlEDw4q3lq33Ydg
1f0oWgiyadl3Mkze8/EzxgU4KS5AAb1s3o+VmIzU7hk4ELMe/aq2ogJ1hlLG97WZ
nGpXewH5GAU6meFbRgJ/+7h2eu+EAH6u/CvjDbhm2iSL5p5rhmGbUWxc+M4hliFb
1yUDtSfZ4DaMIeUZPaaHGDO11vytOJF0CorbUEdSeOzVkQcdpFcTCDNgiopZVwdE
OQ8ElmhukeSFdJ7E5DVkrHgttp4cIkXr0baB32iiL/ahESq7KX9YW9Zi92PMOcK8
DeAEBT6Mr9/qQA0GUGp0MHKiarIZHK1G/9a7krQRsldxIqO3L/lULfAzb/EJ0QwZ
m6y/9YFIic87F7iRb6Fe9NBdN6B/I992jU2EZU7tBkKqg4o6caM8mHLb1LrEHEvT
rOxva8B5RII4nZRD4qOYMvR02xMK3r38xy3VsR/Z08dq1jDMzlh9j+4mAIW627qt
r6GzRMDXvZryH6BxC+lwckLCu9dqx0SlpeBM+5KAQArDgCWjSzoE52nZLOY04zRK
WdA6vj9JPSYtca/7bk3sY2CgsXbxHz3XScmy1W+ZLJ80dTiWV8yfkQ0zhZU4vsx5
u5pUFQoDvpcC/z0I3p+QDsIGxv3nUulpGZEGJx+BhBfDbGCAk+0OWzB3u9XWosOM
D7BAIon1uLNIJbQzOj3x2l1vnUp8sgjsxy7RU5rgR+vA7nzSg/w969bCGiEewqTn
u2ObSmb/lX+mA7uIVQcl9/YQQSaYwuduDI/SDm5hXXL0ZQ84q7+r80o2Z6vMtkbN
bK7mdkeSHoZKJKXiMjl4Q9RXdFKVC92x6jTeG+urhxGe98Cj0VZFVze/U8yw0zM/
puy/GVh228HrgapdZApu96uuN5yl1TABAG8Whvgb+LKWUJsAo4T2uE/cwvdqURiB
lPkjN8NnJ0+OeLSbtgQ6aFDAuVWlRk1vMb8l6LmRSQf/TnmVd/h5U+uvPagJ01Yq
82tPI00PgubDPa0AmcrjAURxsoykt0Xi1sgHCLQTlHxqIe83LqQXY9BXMtTdjR8X
q2BXFKKH6jlGVMteGK98ZV9/oK9Modn4r/1Slv4c3zMGoJla+yJOQnwYmn7aqD1L
xgMDnOixqSaMv1/+LUARF6zsjUMWk3aZosCCwi/MqQ3EEN71T0rzbSj4CkDvVozC
8r86tOGzrSs/Tgy7jMv0uMh6stl6ZPvviJ0nmYl3XqxvOUsCf6Q4yuVUseriGcV8
J2RrOatuHDsTcy4Z3fkJ593SJXRn9kD/mqe5Ratapi/veJ8f5tOzNyy62NRAu8E1
ZIl016gIgXkVSHPqYReXKm7iyrnf7FBfDA9qfqjJxaojdDWSCP68bdScmrNelc6/
Q/u4Lgo+0c8856QAIAEk5z1WqnSsk18ES85RKI/o13C/jDUlsf8GIgcKU1dLuTOp
O0BH11fdfczI7/WQ3M5uXKJm8JnDeDI8LV5JaPrSxnuQTWdNVhliRCHlEKbiu/R5
1ucShty1M8pf3KLiorPqNKH7SgkCXYWx/R1YG6vD7CNtgZOme5Mt2QYjIblyE14N
6PUF4xE1wtG25zYk3OmZrwb4aD9Aq8EaVOKmvoT1LqQhyuoaEQ0v22A3nZ2JisP8
YmUI9+80HireYNkCn38J9RZFq6TdwhPYEl47y8FL+1KsW+JSuJBf6CDrdblx62Vj
HYi6vS+u2UKbwtZQ43dBhwU6ytbmtT7476dr8XS4xr/M5TpdelxGRZ48eyUhMwzw
yte6UAZ6PR5OSkbFukU6nu0nq/Hcqaj+LW5p2Wn4SEaNXOkOaq66c995rUAea2FP
nqYUbc0KERoSc73XpsME4yVl1TSVOVhFpfXcD5WqfZ/wtwX2ZSFbU6YlqxVP7SYX
rvQ8+ESODsks9CkZ9+l+4Hr9wLLNpw7g08GHVqtW740BYoIEKacQyMqj69Ktp9La
FY1dg8ICf19+SeB6Ko0Y66YNYfi9eqBD0uARfskEm6kkpv1imeYJjLJpZiY2tP9d
9FsmlRHtrpLn+4j6UBcojOzHbvnQzDLEBm0YdU1fvgxtuU7d9O8/2jdLOG4lcQ1f
Utl2sRDIkrN7tXDgvbLXlX7VL7aFXufNi3cTOCMA5dTHDy8aOpMx0COdFnD71V1D
kkZSnIh+g56klHBWmWrBSDj+1Oq8gE8AEnR5KsRaUtZGnJYnNNRje+JZS/N13lYH
rDEXyCesqWmHdj7zwD7uBoLmIZSDozL9fwl4/PAsd/WoIYE/0gBGCCCIuFeZ2oqm
tDhPCJYWJZQOQoNMwmnY4PK4QGewSP9qfPfXroUt4/XlPwcPro/0CoCCz63Z1FiK
ONFIUap4PPmUahSfZxFDLy8xdOwyIM4D00sBVakXvdZDTwJfsbTWXmyElagdj2Xr
hhVD4dSCDJoxAF+P22jSajZTTqLPgAXMmBabQDQOqXqb8/nkEarZuFp9zNDp94Fr
PvGNGeRmKfGF8X47y4j5XCziRPYzmior9Ngi9GWxjUc8rh7S+lBfa9B8BnzN1zUS
rJpZfJMguNcvs6naVgNE7RJt8U1BlzzChfgqtvp6pm+HCTqDR8s4r1I5vXQJ3oKT
2yI99Yx1zMA9Gb7+6oFCop33Am67pGV7nRSF5yVvqUBXAqks06+pjYYPwNPgHqB+
qFPno0pFP57Axhg6JdVmhpTTr5Vu+MoKDNKwtoi6b9YGSZyX4kEKjv+V+PbAsjyq
BV6yKuDSKBSgXDP5w/GABP+I61Nw8HvXk1dB6rYQc/q2w4k7FeCP1FCvqnaaVcaY
6f5o1pZja2/E2iKrj0vvt6Rw2XUlWRe40WM1wWBw30id1xJ36PZH0LtUIaGZI+PM
RIxq6+dJIRw2mgprsmzZ9PA/50gHgKPVPGln8uLOID9BdJYva9Wkbu03rEltTM3C
lAdEp6BPXIFUPWbYCw+8mJ37SNJ63ndH9cEJwrwv2ZFpbF2aEdLAorfTn6PyTvM5
xd9uMVqfCiJ1PApEZweeAOI/+HT5O751HX2pnFBKt1ffArJTrDk6wEw1h8+NoMBM
fia2VYf+8VqIco0kClZbSGePGGJivvF00gG2bkVX9ZtjVF7oeQh+GZNSBdWyV2Be
DFEW8wyutqaA+Bb5zT0drYNL3s/wkpfPMDMm6rbPKIh7c4ZtwiiwGjj/esKDmTnG
/E5c89R+dgFp7xdfkv4JkQj3LjpRudslPX3hhGqjGzWaW/zSqlt2ipDDrQehLI6U
7oduzeMksESo8G7sB6RDVFaQR2XlUmfB/nWaeDHQxktU/8TX8xW/Zf1BJ6Dwa+Qq
7P2FTz3/Gnfj855tkyYoutrEBs5W2EtumIKmiYZzCGSk1J1f8SiWMyjjGSYqalDE
/hXvn/c3OUmf49iVW77LKptBaEBZs0Kk5zlWPtJiHTVcYoBUT/SQcQpBU57gKClX
h4zKHcL2DyEH+V96/7VQClDfzntM6p7K+gfyVhJ81DVtXl62E2DsRs73CaqH00W0
ca+j5FWNAdDgm4JEzw6EP+cATERHXqb0PmuEKnt8kqafOFaOcxfOJBGIB7P/W5hc
qegk/nWBg9J3YMDvSlSh2GE8qVPZ6jPKCSPp99tmwMHajOR2FO7BEbFpdLpOCkit
djbAgLD6yQoI3ki0zxX2qB0PDSyxovtOIstU/D/mopUomFyYNh8RYU5YeWrsOqX6
IiDqpLfMt1FxeQUJjtLNuzB509XNoshXiSNsQBhBptwoq11vF/Fr8iAkIhE5mh+A
IVp9ta1N2bQ++LG+0nCf3epZ9Kz9XlpsWHnJ0aTkXltM3A2Q3/bBRIQ8VX/7t+Ei
JBTN2UPVSI5Vl59+/sOiPNsDlCEHm1yCUzOxO1Kr0x06RWjloILa9NHJ7e7wCMQ+
qTqdQz3a258vafNoMpG9QcBFlIA2T2xPHnqdBc0kC+u8wo8OGB2lfDKGGi+thS6n
NJ8zF8+LzBm8yKwhAMpZCdJXaDy3LmqGfYaeAbSjDj8FqVevRtVoiIlX1AMNWyjT
sU6b4uy5TCTpXquJgqHfQvPEmU7wBTZhrxH/IVTPtqYjXavOeOvRfMzaY2unj0d+
bLuGGewOvkvN4gDucOLo8sAbhJ9AwaN90jhnx1pz4jMNPBqpcMnCL7YwKhCmPLZC
R3lYb/IlnOXP/qLxyuj1W5uhw/pEMg9IeCEMtViIHEBbjHI4DuAVAoj9bbvW0CpB
GVlU/3AgvmkiiI863mxOE64qNAqux/moYV8XZTnthmn+9KkN4BniuTNaqbavt6dZ
YXFjcAFBcktSszLAfQ7V/T7vCO6ZNcId9/AoIEIQkJm28/ZwrdcfdTbjdG2rV2Gq
JPu3g5JHQ5TQ9llostrsFGVhm3sMUP1Lp4aGsAQ+A3M8iGOuz0fpIFM/ybi2WcyQ
M7w904MeayrHccaK/vIHTmzXX8/t34ZOZnUiOvpyN7msnplQX3Q4dT6OmQpcg3Yo
kaoKuR/UxmV/4sBdg08At4jaYl0aCG1iw2YL5fcz2WeDO/I5O+z0OdW3VfgnqszE
rd5jO/QottkMYO4fCYKGiELstDcLUfrKoz2Ou4r4kvKe1N+qun6xpbt12S7wIudJ
L3m6nqo1KPglg+Ve16fCV+4hOiy2SeNReywJTVjxqm8sgggeXT2IhFnJr7oShOPM
JwOFPGiosk9GQnErq8UvAsampWRINp6aN0wyGAZevP3kiPSFlV5lh8zljJmz99kx
wAXRKj9fdEjFb6aBokJ/5qwxxCw9+pH9NYti1l899qqYEfEiaNNIlWeKL8jzvNg4
0YcQV7rT0x9XVHT1k/b/IG1gdLVa8DdbdihugGVizKDqcAMthxRnLfZ6FCl9HdXh
T/1iSPl6GhZR67uiI/qeulA7u77Fyncxq1MMW/pxcHqpUOWRcigcl/FzpGF+/TPL
vt8WMqmwUyxOnZXsUqjvsquG8Y6WLvzGEk+AwzbvLqxVuq8Je6ryMTxk2aF3rTgy
ma+b3NJfzrblsR7RinzWFtrIMltpS38ig4ROs5Nv67zFHe5N4k6WTmK3U3xqmh+i
nB4mnuOrpptk74POrFxROZQknGofqaQKx0/QzPsODgfEm6XBsiGhEMEZlXAtVwLh
6Kh8OxvGl5mMimtemC3vhJS6+qIT4JQCQZbDBGbHanmS/CSdFsvzv9HnMX+xe5sL
C2uocH8VjA91IiiSWwthMzicMSG9oNr+CuunZk7QuAv2lYkjePMe9b5zTkeX69SH
4ZnwTdDev7u4TOD0zt41HxUCWNd7lzMjMZzo2BdRPZtOJ/2PDIcH2DdpaqlVhUmt
gv9ZZB1a7CwBNbA/w/Og0H/cxJo8I7S4KsF+2re+2UsmIzKy4Uzx71WeHj1mClPc
33mahCDzra+H5IlSpSqzusoH0cLuLyKFbBZH30Pmb5qmCVMSPJYCy6Q/bY/mh2Wu
qWUAibcM4A0mzLXFZUIBxKgksJmiU3MPdhAub+u8/jpqN98cuegIaCfxKqnaR1cu
GUNJoKlEqx/aI1G2hhFo+gUSkLIbuI0G/7kfo7COxOgZv2mK87rPghyfkzFgT1+M
ngK5ekQJKa5pvvUUl1d5J5pRdrRDgRQ9e4+ZTyxCmwqnqKGtr02Mgoah7qylrXwY
/g79cERE7DDgr0UblRRzHfh5rfMXh9llxShkRiLU9jXq4yrOzXCeC5bYNaVKuH9S
jhEYw1koTR8JnBkiWHMqBIoZ6rMLDUnJpd7rzTS/9tHNefDahtXA0P2Bpkx6xnhD
znpkqWs6OCA9AXhjVmmbmNyGnIlc2ZyhxpG8J3w9z4JbTsZmEoN9XTKtaOoFJGy6
vvUSSsWaSY+pnG4oJSU+Sxh5DB4e57Ib3N4u/C/8y7nb1s/jI2RmTVmhghoCk7VN
fZG8Ki4WahPD/wxrdM3UvTS5Yw7vCbbG1SCH2KZ/LoJ8lQJf7+mPtApC12cY6WZg
AXbqSE1nBfX9Kegx+ewfYr6SsAMHgyclR+ETdzAVNBY/B+3ZdsWgyDfTEaMuAZxz
ous50ygYcHz5Fbpk+TpM/aIrM1a6VjxiES4AtAVm87mzvE7VHA6A28sUuqw3FIyz
W0CEqREHZMQzf0yHkzElsFKlnWcpKPGoslUv3mr5I5I0RUqiyiIs74/wX6WAYmvG
EHOPcg0bIKtzFhDYovz8k+D8PN3k90Na6LF7Cqk53qKSotaniFbvMH7X0u9hX9It
5McY1QY4wDcNUu7563bFFU5uuiO0oW0v5EZHhnFEGL4RBtc+1FFaebQ4RsehV7//
KVik9e0YtypNjYhpF2yT+cXyX4q/R68kM96eGE4UaO+Aelk7rohDHli2QxC0MJPN
sbf3SvOOjfCptr0Ffl5G4n46SIGpEG3nmD3CherzwFn70kqDHNgU6YuLJ4s65rg5
wnusn7aufTv7FRPKtBJVu7MwI4UBYk3dcVhrLgMoaWxVTxkWt1qqf6vCEFmAnBzf
g/c2JHwSUMqb153dgNi0/pilSTqGGUs50kWrHLzE8DA41pdCFTm97QtU8MpWvx8r
zUJt0udVkLXRG0kPXr5Jqo1qvxU7seMWzJwZKRq1dsoCH88qNCNoX6IOTRkdaSUT
mVs0DS8voWl+rIB/IzkRqNOEmr4Nw3XyCaGAVJdVzJ0LASLCha5lKa2/07DRLU0g
zKFBhsyTfNQ9bzaeNyVzBTOaOwiPutGyb1V2cDzWXjZKY7AZyOwCFEMRenUjm8kl
ApXE/4ncTGTxNNuhsPc1HfPqbjIOmqA+8cuQPQzbKHycX0lHlQlNRzijGKK2WLK8
JmIlveeZTn1d69MHbMkhM5+JttIrCzG1hD6P8rRKklvr/0oLxxawjavzYs5Dbe3o
KtZ78MNODhm3A4Dwms6Xt306zy8nWO7y/Oxa4Y5eZ6/B7tfiAKkcO5/Ajvv1go90
bnwE3R+ktkMUk6q2KnfhdpCHPzpoakAGIWTdeGbsKvj6W3DGLQlaLGHn2ZD9+QJ6
PsIKKowdGO6T896EmZyMx/rb9DdhusonUOMKOXrnMU7htlBC42VvdPkVqQ/clwHu
AuKsa0NX9dA67DOy5myajJcLAlyszlZ1FW/p3NDuJRxFfpDJXB2FYz8tYrHH3DNn
WtSW33Wsc7oWtH6n5n7CIjWmfSIN1vS0S8JMF1H1Zfb76sea426I65N78b+BJeKE
AsedN7+JKAdceEBVuYcnTrvqRdnf/rlU91yv3R6oyn6/riM73cLuEToVPuWIzOWu
6RV0OO79yOlN+ciWpG/RmSzOgKxAN4Euz1TZAlB1efCKN8kdJjteP81v3Y83w5wu
Mqat7t8Z2Fvy0yN3CbjfgKL5A0yP5mSVQ8yrOKLV+5nUplhoif5ycrY+ZHe22PHw
+6z5BDbvumoIhi2KXLQLhX/k+zOGGOjElPAKYLGfXItZZw5DOCBHlGht2r9Tlb6h
bNbDIV+GsV3yLkVHLaSMvl17C2iNbktaOBVgcvtVh7SeN0NzC/pxeMIKqef56DeF
M3P3kJ1DxHUIT9kZC7xinJDMBbMZGxE+rm6BUOpMtZOoMsYlPnnuAffxbWgBNC0h
c7xhToJqGar3WGrshm4J8IFqF8REHyxgEO0am76EdgqQ1fLSlCy4Azc5zgcALcDL
GmG9cRAp94iPqGhHgpE8MVDk+ojKnntbAcuCFzeLb+wEfGczUlhHm/MszWPQRqFx
Zvxo4VAE9Ujfux0zMQ+awML8pe9TkcQYsf1ECzqF4U6z+AymrjzHqu4dvOPS3iYY
jz5nMk2mgBDreW2J/DjB5lthfBlaCWOrmd82mYHmZe67p1MJ8xKm137RRuDMslxg
fWMcAWvlsbb1ygy1NnIEuFJ2osWogMEUGF5D1w0t8jXc2yMmZDsTtIjLJHvGf9FE
rWR0phe+YnMFotOnUkIHyNCs4MCUkHU1KVqRgCGjWHhUDSt9NOZom3MK1Upd+AV2
kl5ZMR+H/dZsyN1kYaPJid8SRwf2rHmFes1+s/+n7GE6XLQzBa6zLNLsPNK5y0MT
dNrOxBJZHtHs0ehAsgkn5IzdBi0REkOd80t8mG36rye3hez3a0awsTYkTCxITwCG
DlzvJMy5s/CPCg3y/cuTJQ8OhZRBsvxCLEf1FDhuf0j/Xce+mo3FvBfgXT4hjYsq
v7ZryvUc4twT6Pi1DW3IWuRpDsXDv3eQJkO4WMIJHz+EZ/q5fWcBe5Twgqmw4C0O
boAtX4dfnM8sEDyxzewPp8OUVzA6V6D8q5lx0gC96EPB04yOfwMGohHl8w0jZGO2
aOt5ZstwqvPUwKr31Jcsfnd+4rgkQUhyne1olp0ZqA5/EYYQ3zSBNlrVV4z2m2Cu
a3LNqVciDmO6vX+GF1986zadjSX2sARB6q2qbhVsVWEBUOLxMZmKW+v4ut1z/WmL
Gm7eDLHhKAEkR/Jd2QJgENNAEi1+dJVk2oPjeGwpDoszru9L0HnwWnD2uHqADfd+
m9oNKKcznwmgc8t13vbGNfJx/LrJLd64anCjlCZif9AISQo9bc/malc0o6QaDlQN
9sinkMc0RtroQ4Vr4kDO+vKIAMBOaVS/c4XIPFXJdxXGzuGnikwuo3BM8BZOPyiY
67dcxMeReujgw2kkKKE7Egjm72icxXX77PkCV3Kn9qUZL/IR00ydnAudAmp4nwRQ
fP6lowVNi7EBTcdO4P+dEm0+PBwr0TQooYmMnltkkUnHdkGXRqBjgezdj8aRZ8g4
BnGJuHP1me29DKpNpiCkYae86OIKqFwAhCo9jDmrx/B8CTMW60Px1/Eyeu3iGYj6
CRkTylu18kY+CeYK/B3Srd0MlAF4TuGZ+wcvAUSLWnk3cDezxD2WYSQ3ZiXzZCc/
AZFsc8ggSRA+TxSyDPR4gTsUeW110hLvKIv64yHnMrx07C1C+Ec/CsVYroZjUDJA
Ve1vuQBxfNA/wQEslB1L9eQafUjFu9gXkx0Moqvpa+k0BKvqUtTxBWlP+rwj2GIe
FfxJl+HfKyAFEhAyfEoEU1UJq5AKAj5kG/Cadb98LCzhe5ejjmglUKHAFPeM7IMH
CZy3qgQLS4ylSDvSFfomkMSNQL73eY/ajfO79ynrTrb6tyeTiJ/ZkaThnsmymOXm
lXCNpRtQZL9cWjyz0geHqHYUKStruVtrvU42QvHTmzpQkwQKDXoPJI5OnylA8bOW
aBegNJksFom5tlxo4JAjOnYOyfTRj4ua52Qz1TK0t9XUe8EJABN4Lcvpr7WsLMXP
8HgdyvsOEPPcutkn5t/S2qe6dQmeplF2cAO1uPKpC45dvzQJlGppro4K82LPnK4w
cjVPPmRtPymySvnjwho4wmUBWfRk/AGMRj1EE1RryLY7Ead5IlxBq6J1Y6x1Kla5
uG+0wFih/fQZORbMdnz0TkRlJjFNkG8pRkTtghZW/lTB9CHv612y9cRaSmoWq2Q8
Y3PYJp+bTPzLmPMtF3SUFiVav6T1Ng7gDwhAx5lbvBndkwl4HZc+hK6zWK6P9teS
IjTuSXW73KTyFGUY5O8AsHHLsCIEmLDXpJMf0D3b/zzRsXLF3RGCDYxy06RMxupT
0Ow1kZRZakTVlVAH0RhuaIy1Xa4xUYXYGnm1AlAZIDrDpHm3tvHLHwsHgL+fuQDV
TW0QC57taL+6mX26PvcM/r5MWdFGAMTaDVnSsQrhiCWpHLod9GStrWhqjJ1JmaEV
kEH/CDWc4KQDWMAEESv4EhoBIiR/9htu2HfOY2rOh3BawYgtWJRLirZK+ScyE/L9
JmO4Pp0MEubBOCUt5eKl2RrGIG+j5+TeeLwZl0Ntb476Tt/WTgl8YNf3FSPmVAKS
FrbEGcVnYbbmLDij/KWD6yqpwRS7E7BkE8XrTQut/CNDy3aGLHYNjRkz4CEWvYtu
DZH/5BdhYpmQwZjXqZyhwZM168v/bCy7HU7531p4EaaJ6EokrbE5mH7igZBsZEJN
ZQGeV5wa1xTzBO7xiJriKapPW42D7BvoaEhlNhO4NTHhPoGsT7R0bBrqXB5URVSL
pearW3IZq9fJevTaEyhX2yKu6d88hbXr8swlGDe1/SLBQb5YOBL5H8oKg1Xgxveu
GObtzmI4l/h1UNzXYwVLgGSavq1lwb9AEYoqKNpoCBB5K6cnK5izbwRjx4E4GrxU
W/IXh0X7E/yUMto/LjHL3z9D9cFvaqB0BKj470EHBtGzUvudl+9nCK/mQU68wW1M
W1WiTmBrn8Hdaqv9a2y0alJ2w3AiQAHUnRt8SdPPVzsxQn/Ups1qKw/Y3Y3Liqjw
EkM1zDTwvhtcEKCbvbsOHXxJCZg62Q6bb53/AVP514mRhmfH1CqvmXasgwUvIhOs
bq7KSE3+R7WPdU0hU3SeSWXuXXkKC/fxH1ouZPnhjx8T5ouYzxeZCOqrBnYkCOh7
GB4iEMwjV/oHTwE+h1kHxcP0H+Mk4JoUyTMljCcRzSU0N4tmipqgMfrCtYeR/KmM
n8bpMOhmG5Kl0HBcgA+xL9Z/ngGYCPki0EeeVcOHa2yHOVwqd5TfCD2aBNudUEs5
+1Du021Q4SMV06596m8UL2E5qkBM9OB5VcJWPr/zvUuCx/mfx7gbP+rBrZJsNBwm
0JAoTYD254k4jssyJiMiJbLZZuxP1AEnMTfzk/IM4W8CxvqU+TFfTqQ6BrFLTpOX
SN6LHr7IzaWfW3TU2x72/pu5HMMKm49Yx1r3Bl+dSZgzUhy+R8BZ4R3FbskWWOxc
b2J108TqCGDfn1lccynvWgx/QynbBv9jzel0r+TfTtE9Ok474vOtti7LjjlDp1yE
G9q+5/t2I0YwAtPS5hm3EnwzOF/ZtX97j82oRmFWgLS2cSBjrM4KDOqzVq39/ef0
608l6VSzZiRbsmBXlzbWJRj0/VpU9nDaWvYFSrBctgFNPX7ZicApBaiH2QRdipSW
IODUlRLXSBp14Vs60/b4eBzfnj8v2eSBffOPQA9INsqdbdM6jfGyZLqtN2KTyZFm
XY50BX8QY74QmlZzg1Evr0G53WyY3uHQfrCt4mt5Zwxn49dcENTp22xCYmeGo6W2
HExah+YyIwGoAxpHDu3Crw8D1tDwwvTco7qP9R7bMyE4tF0i5Z9b6EkFgrXndqi6
Cc1ZrrGjl7JNYAmXl8LlsyfLwGDBKQ3dOtUg2ZYHY5u31YZJdkr574YjicHyMODZ
xdj/KQ3pujHHjNR+D8o+xEm7E+BtRB3RhOj478cs8aVfZqG5VrWjMuH/UZIGRPFb
bXZU90W+5sP0dfOBrREbw4B3ms3OA9WVSp1Xse8+ffZW/bhwrKRfxMWtfQkjmjzf
1KlgWhNT8S8/e2m9yafcVImHnksANSD6t0FVquO8TnrbSi4DMpB4ICnUvBV+39lo
8hneoo9iABPnt73AvVHEcaQqnOB3/ZkACjXUXCG2c6Si6wUAnQS3i13PpFKc46KK
vioUmZ+U2HnPiF49L1sYzhIu8Pdea2BvMhHI7QHE2RlORLRwiUhlpEXgae1cWFSY
26JPU+Am5xEtIV06T5HUxDy96DQHdv4HKksWpXa0N3CzXDYoi7x/3HhUbrk4t2l5
TIq2DfWOuYcGiH9j/ohn6Q2DMQ97DQDR40R4xE2wqJFqnoKLhBHUT6FJPSix4ecg
1V+iFYfudJnKXhvFrtJUjaENEhZn8WakB33vGCFyC90w8xeIkUAED47+S++xedmm
YVXua96t+b7KcLL3APN/aRyuVOsUr0b9Gt5Kiwp/038sUhNWe4C+JccnEkCWluAd
m81bnuAR0ba6zEeFRAUCjjQRr2PmKzanxY92oLgOKE+VoIgEmpRqiq2/d3BxuR40
ydyL3E41rZSlZ4ZTAUasGz4a3+CQr6Wj7l0ux0zK2FOfwF9/KSGnz0tXOoYvAYPx
PM7x8K1HyOHtkw7tTHdKW7qwqr7OrY6ojCSnVniwTzn1lxmAnBvrIpJPc6CAIu+9
pmAW5qxzATQBtvu5BAzcM1R4a5EJOBJ4aU72471RKkXAgRYhPKZJCSX5++NSTtyI
DNJXKiePCSjnovUU33cJzTrp5FgMqlWN+QhawHLjYPqLbBd5OP/tw7YESEUv5ucf
WKLsCwVEKd5Ip+Bftx5kVRNEoCP2/8ZJ9bNoYg9IE0I/X6l5Aem9vc12Bdl1YkL/
G2JTN5R0N7qUzmqRdNLZzGnwkUNdHDNokoyLj73YfRrQknfYqkX3cvw6XRR4qbHg
owtyBe+rjEFnumarFjJ/FY2yWWjbFDZMkFUHwxq+YCoh3z7D8MVSWbMRIZb8q7Z6
9gCySH/sQu9WmfSHdfdWjIAywAZgW+4dP/1PKAQxVaQrW80D6UINRlQTELLT4V4r
dB3/Vr538zXDIRP8YESmPVrdQ1nir8rVonzLb8kUVCwV7XE7BYHUGeFhHu8HsAdh
3CJDosYhxnHT02B01lQvv6zv32w1jEqtDoDwKMOLqwxs7pfITTw4t1/Q41F7TXEA
1HuCQkyQ6jH92PSNXdz9q9JKKI2osIoJKfScUGDhVhnbd3JOiB1p9vgNvkR25QsI
wh7WwQwf3jMktn3BLL/zfETbGwvrh9kHK7TsjUzaE9iW+aMSBDFKgjTLR5zoCF//
lP3+PSN5kfT+1JT1QgrD4Ed5u5omnomz2WHF74zTYCGr28hTSwRl4lcZ+PPi775w
n69hyAk3Eb2OJz7DDeaP92eERjtvJYiERSe0S4MXE6wUIg3S8PXjADhUbZnbfnD9
QW/hGbDbBKrvIGiDojktGgW3lpII+TQjeWr3rhP9SS+WA1tvcL/WueAv46oIT/YT
IVlZVHoCxPXb4+hzxucNc064NxN7mPCjNfHQbb+Npl9B8PwG/yZWm2Xt+J2xyiDO
KfqfjruTY9fvU5OUn/wXtyOZVL/vR0vzya+Flrld//twUhvHQ8lDIgZD9ylbdb32
06Bvl5sRNQDlybn95qRXcsFhy1H16ZMLcMQZlCJ0vz9BV6sjNltE7YccNW9Ma0oA
nUNnoqqmTIwwOl6vLI5bWnXuoXI4HFtiW4E6pcZJtqQEbRCLcyghp+Zm/0+OSaB2
geT9EODJ5BKDasgPrd3XuDx6nwMQfF2uAQwzAimGYKiNehsI8DZtedCxJeon3SzM
Pjy+u3KNJTnqCjLz/TcJjj9H+1GpetztKxLFWqZKdaYSWC+PcngrjMixRdPBKYjV
Q82IfCm8djczB7x2DdzCZm38J9ojb7Iqv7IpWE7EyEVbNJq473M1hQAAgPA+jzhA
ShGlJBGQY6ieDQZ21JDfV2aTnVDIWIU0F37jBEtcsGLBeftcA4wsvEEGtcOhY+YF
91yPrRxyB7O4g1GFit2jIXK5qfrIx6jFdyxYf3Jn4g2l6heximFCZscASRuO3gTu
d1UHr1nKs0MaMTxxhSuHW6F2/WTB/VJX0Ez5XHcqASa5gCIWbDf5pHKB8tRN/ZzV
J0TQE5MO29Q5C4NkYk87AR15SLSgKDHj8GhQU8Vrm4zs5D8xr8RTlIUlxCKMRufz
ryWadY1jkQlvopQR0hLYS9KOAlo3XpgPmsME0kLw51KvacfQt0k+vvc5SHDZXLVM
yQlTvT9nQQkMPLGk7xZWbUROuzFQugO0Y6O6/PmoQJOAXeLAxvMHlQKGme/6laK2
/pvrQODJhtM+8Iu4fGXRNP/4yGQR84ZgUI4lT1KXlMI4apPFtAoRQBUMmu5ul2ol
dAQs2OseANlv1TV6xOk6x17+iw6yvUjV4gONiWePwplNKTHEEgrKglKINQufjgSN
UfNG6veMT6eRHF+YOk1dxIPtEFbUcR/n1XiwGO7T8F29FfylsKoe65zg3Airvj1l
zmK542OsbXEFyPy16foIRl1Pa5dtZTiN04xY4S/Qbk2ac97PZHlEHcEtJQI4z5GV
fqD+hPDWunMOkZP5akwoVwdZUQwT4RvSU2tQkUACM/cHgJ6oEau7PtgqAs5cFGQ7
xv6CNvlgr43W90eU0GwcSPM1gQJUN21XqgOdcobkm0UydKTjivr1rIzUB1Qe+e5b
IN37YvjbC1mzcplQJq49PP+w1I02gjbTa6C3AND5QWOlffwXRawi9phywbsjVKoV
2mczqAnnpe0jABQ1zUuNPHwe5uWhntSqizNQ7umHzD70o441/36ngOBRJmXhHyR8
6UQb72/1d1pXa00TssQYsiyyyEUrObuVpBWHJQIwJN0wgqSLmpf8p1HJU8qncpAB
dkzgMgANDIzmt284EO58cy4/WnKnuuyaGvDxaUX9XGR18g5nOtmdLz8W5usX28M9
qFrMXxtECxlW5fFXzrjf4Lg42utQTeR1qPcUdcRis/u0AlC08FMl6Au4lGZEVGQ8
95iRhrgH+TnzEEjmtSSZqw/SDimY8n06thkdjBcPsE/Dj6nT8WNyu/V7P+IU3sc8
8yuwuprr29SS9QCsHRyfal5UBapjzbUTPLj1s4R03bS7/bQXamH9qwnoVECJc/AJ
a7Z6xTXGOGQ592f8fA4933DRU8yJFEpRS7Csv4HTu7wiZzgFF/6cZMGAVKmde99E
f7KqEV8+I2rvTuInE6Ce3ogUrH7DpGaKgQM8JMO7VsVJ0VPq40sCLhKQm3Dsgrr+
cjr2qJlkgFCO8KCKFXO2wRn/gOOOO9DT++SxfGkSimoznMryE7FgbvSMlRDYuF5K
Ni0y7BkAEiciiKE7jnDLI6XDufhi1Y+apEXO/GgMyxpkQxO18UGbiEEr/yq6HLKG
tm+vqYGpjP1/0LNrdbAcuQE8/OympF982UN5dP97rn9dathn6olSiJcX+eumW1DW
tc163OdtqWvlPNAOEVz4TuMgW3uebslTnFM1ADhSztkoDUk25NWyTwr7dlUFqt2z
NMtCSFwnlX32BFcoBmFfZJKJ1igR8+h3WGpVfjHA3PD9lwzT62Mz7UL6lLcyruNT
hvrrD5HWvQRCnIZS+5ncS3bkwtqkHbOP5xnkdqFOHB4csnintw2c73MlR10vrFQ4
Z8CS9sxQaIx0IVr2hee0IwERhIi1H3xKAfdGvc3KhyWnCvfScEQK1VjAIgh/Brx4
hXHn/6osRTnUNJ6ZKR7kT7S4wyX+b6o8LbvU+Dg0FFLR33Ok6h7mD5MHfbkEhT6m
QytO9uAuz19sH+r7XlTC7d0bK2Gif+uQaYkWvFL0/Bd1xRVYg2I7n/hIKf/ED727
3WSRcrSr0VPz1NZSTU14YR7aaXKG48Taq2cpTYuA6A298vEQ5XNlpl1ihaPKCwe+
O/wz27w5/5f32lCYVCKxaKcNFZbKuHsrtXNjSlY9cxZ46IFHhfiw8d3Q+ilgbC4e
JCrH7soU7YPXpHJ+G2g3hQtpwfm3i21m0xXEBjqetyhPs6hjE6DqN9ioIa1EIqkg
9xyHemHSKxRDZnSsYkH/o2PHTkMlpIU6yb6lMAvxJLl+qfUjsqUgZ8Ug2LGwT9ep
JmRjI0T5l/05XVGnuwCj0FafWR8s0txFw8UwSjO48mQXz+mECtz/w3YDxjptN66Z
/pbRIGAXDY0Vau8zdHHI849uDqF/oZdC4Ny7dVxCa+MocJs/XJTea+MiVqaLQsBa
qosN1qzWMg6rKfCP5Jj72WAdqRr1iGIqTQ+JtSc4/8Kztt0V9jqR2cxbwMat9Fwv
0QQ9FxRLCo5KDSQiQNAINkqIn0ZyZ4c90v2+C1uNw5UbgYKbzaOlSpVdSF07MKzF
FavzAMaqMG1k4edR1s7Kr3749kseyJi+GCK4zyI5Bx0pl9DIcc1kO5nYl1apNAvx
KCyUQMRT5KSlH+bhpJejOyWU5Q8Gy+k5lKWdPxIXxY1/6Ljqiyw0ImIxXsoBqseI
3RTf39R8B0xtUu3ZWaj6nVa7rthZLIptE+k1HfaqJ5vUN+uwnVzateMPJ9uyEG4k
egNEK5q8I1eFTAhg9zEHWJemJTVlgf4rZwPrFqRhl4vy4qzjBSoIkxQalO2/7Yu2
R8zbr2PghRQQb3ObX3SzcbSWMfhEou9pnCZ/3cKqwRDFvOi9TbfH+byCXsx06tJI
jjN1HfJp6uZbim/vthghprMXPCu+iARrvB5woEkhyhwNWqP4fdgS4Sush2vGf6i1
OPEqgMKwCpFO06zWFxM6gHl7NTEkgZ5kEQHyqvAwc1kRLfO/5iV2q36d9Yb0RfUi
WmX2qZ38C3rtJMOy6zeXAuIuX0d9e9LgSI0umpsFBvP3z/E8YBV/r9YyeTw7IiWz
`pragma protect end_protected
