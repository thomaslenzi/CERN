// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RAZftgB5cMDMuJo/flC+tIoV5DDtrin6jfWVHoNC2GMTbnSAVUE8P+Qvk6wbKIRN
VZbMlIFrAy/LLlkKqnTq/AfGaSeKp797C3/Y1+foGYt+mC9diU6IG5BYG8WsQ/U8
vV4B6ToRy7PqQxrPywgZy69xRzMCpoM5hVYtU+Hxnnk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4400)
iaEs5qbe8fJHTe0j+pZtpPQE/1SKPvBIDcYMhxogBQA5/oTZ3yWMFTLHHLihiG8f
+/l6PlyoWoe02gmL7Sd3+yEy/SqOcBq/E2vXWoDnzgxDvEgl2+c+R4L1Zsak4wfV
dlLNQfbPz9VsBPPNgLGkxifNdHp8NiyxNMjbJvEyqYh+qAC8EyeN2IZBfXqci1OE
iuCEbr4GH3KHNhJj5rDi1qkc/iHJYTqjUPZis29grBWrC7I6P+VyzYkp8pNS9rmv
jpPOdxb53gn3yYaL5/P93TzuOo7qET/STKalV+y7zSNMMCevMXfsad0mrqh6U1ye
q4prQiS2THtQs10ABHrieYl+X9ymNxzFx0DUX0kt9GeJOvDiRs21TGH836BeD437
0S+fddugFFvZB+ePkJffPeB9/xgXRxbitHTrF5azTxmyIQPZAGFTDolaidNmCEd9
TbV6cKzPss796Nud4WYCsHEqMdvlqUPjREHnIw7mcB3qbr1ALvXx5zArDKz6IsT1
sN3CTB1sAxM5GwETLYAgGOT1SM9ku1HGEBZp7JtBtiV4u2RQ0X21JMx9T0L489Fz
CjvtCuvUVss4RYfatFF13DpNRvrdxRuGGB/Wq+YdEJ5xdpmgTMwfnezSSX3BnJen
HYStKY1P3fyH6hPDYfXuBBwseYvQzGBNMIIoOVdxaidEKiKMuew97u3qvB0347A9
O22zLoqfmwSSfYuyqtr5w/orJUVlK7mlvPH3uX3u5sSdUTk5h6swdDLVLm/e6SkE
L0T+bXjl8UISC626zGgEfdN1ulxd2OKHdVelev0OWZTObdYtPfMA2zIYQxAPY/py
cH/i5mSEUXUwMd5+Q3j3UdhpMAHNDVcV0SY7Vcy0jmSBotwYAWO47oBZUO12tOCT
m+wOK9gOgzsZPh7cumdGUeo3Ks5PPfHtDYl/CKLRrkyL1jINYS8ylDmdjcpvS6P3
aRKNNJNyJzfAFoYAA04K3ibavl1Cc8PlBxfByQ2kBV0PNKkPpUFAJCOu3tYTeIoz
lWqI4TKED7w4i7oHGD+WnIzjfqBMKQVaeANXMQeWbPRBAhejLmvOg136XkLXMHq4
Yk1YIpjs3AsR0Bb9ISh19+DVN4F/Vgg6YO9jEXwu5RULF+PsMsXtmqRK82Kk7HTZ
aCI1iophYr08N+MU/JLnN53ihrgA/IrE1RcFUpBF7EozxJd7SAEUkyHv3xW+qWO/
SF9SWsV1T+8A9NhVlx+Rz24TkeCwCp1d3vBt65Y2sxa4+pxxUV+O/NTy4fvxqz2z
DVLsKihbg9fVVGNOe6zM6ED/XxEVyvSQLVS6TJhsku4Cg7WisO7RZehGgOc+d3FF
ZCNLPoWeylib8ZsJp+ndjTnAjhPe9XULjWoyTtorVnKxh6qpi52q2QO3yrR9mTx9
kmMlmTzEbu0Q3RZ+NT3lcMiL4ZNRzw8bkv+S/6n02mUtQk6C9sVQsplrtGI3TD4z
TyVtOHeWB1sEokKOm/Ez6lP04I6m6WZz4WwfBHEIg3pZ6oXEseJLCg0iuuXIQfkk
jtreGyAeK7m+24NlorKa/AnUKPrU8xcO+gYdNPjEAG+62TbBIwsmVQZZjYCUrsrt
Ba7Non/Z6GBjGXRc9dC6wmRcKG1lN/tpzm3v4j0k6Ycz4vj5dwsXNkwAjRhGUJE2
lfehmBArF6saLbrWrgVLntkrvAi5fI0spLXCteZiK+R2guKTSjfr2QHKGHpcfflb
SCIpUp9bOZAEZ/qUjXQGc6yuRU7c0uWxJH2UB+6bT1rlj7kV7P4Pugl07wgi5YTK
L7NY/kMqnOh1aOHZRfG5NQdBdO3R09EWDWdRmQo4vv0RB2CWjqmTYewyeTSHR7a7
9GKeK1HmkOoxrJWvft7PWBB00Tqz1dUNzoY3WGYD3juH1yJ/4waemazZLT9MKkga
Xxe+Skmc+cpCCn5sE+P3NU+vHiyMSN0YfGFkDzth3949JIXZzG84rbnuEGKf6R2Z
V964aUhiJoO61TipPccF3mIYtEdT5/uE1FGwhQT8JNRkkio1YGlLALX+Le8cj6M2
QZ5KngLHCqxDQ/Cgi+quAjcjyo5rxuZzJ4JGBkyd4/XkTVeQJTtQMXrWwYnwbf5w
+pA2/FJoNJ0MbsU3V12VUbo9O85TdiXIExW677SbmOzSQXjNO4lvJ4UO02KQ4M8o
R2EoYiz84qc8PwYBxcKTU/0jRtqWKu8+B761+ygxuq6nUc2uJMw0cDQGRoyD//ZX
TdPT195KgeSJp8Kp5YguAPy0zAp/AuFH5iJbXHd5KxNpEDNfLY1kI+vf1lypuL8m
/HVExWrbX+sayTiHC4te5uNuB2t4EMkBAJMW6ckMsJmvaJNTnOdLilI4d/S1kHxy
3ipzq2g7OmRcq4kbzADNHuDjoqeEijWcKGo/rovtiZxEjOlG4+Sgil6zkSOhBiT6
eE/oUGQPFBUfffYEoM7QTL+XfazIymW9HsdtjBCaULkkjzRNYY+m8Tgsl6CANxzg
I9S1q4rwBxEtmT3So70TmHZqttE4MeBJjtwVFpEGWmJdSHHyp765siPbWqxWb2bE
RnvbQcx4F6bgR/njo3XqDZ2/VBLvt38farFWk/HG2tQHYvmIiI0D+lgJIU2f/m3d
jrVKZlYqfS83z2wJTzeaqGrzGdaNre3mivH22crw1RbAh35Vs2Cp7IPrr8LfhXwf
unEQDinFHsXVGtLnEYdYO0s0Uw2yJZAO+9hI5o9hbOc1+5g1muWT5WBZY9sQQyWw
z4t+SwuuTN7I1BG7828m7AEIuNsA0WkQcDieVBEEmXQABjeuH1Jm2Rux6Ja5e9ND
5aq4EQ/ry60nDOupJpJGxiveXcBjcyyZfuVmDoN6Frcaz+urm0Y7r8YS57fLnv3h
DleJU3ov4BPRALFabDGYO+hcdrnAE4HeScql0D379SpVlC+AIjnFjhxB8AuUx+FV
oBCMkfuze4KPn/+IhmGcWczeyLz3giFV2prlO5A0X3/fe6UY7EqvxDpQhKiFklyE
iLw+lyJGccklOMvn0yorH5fsSpGbDf6aWnJfVfT70kdKJulxKwD2ItBlPeMpCDZW
dyaWXZZYJlDQNKcW1EzGsPd55FWehzBCduTyaOgJ1akYhHYL3Na6cB1o27oYSvus
C3ROd0RlEChJACZ3SKRvmmolEy3JhUg67rJVrDlrRxe9Gz7sky3K/mjv3L8zqpkr
6G03xJFG2uIYKQId1U6CPG4patSZyCHNhk9TWDa3/g8lfd+KAW5hoP0Z0G4v+0ak
5AUVy3XlnNM3mhkzh3hNt1aPoBmCj75+NiCQfS1ZCSxdOCZlAdAiS7fZNs/U2UO+
L/1g64FIBmH4u9+kaybKucJItJaKqvBgNAgj62pE0/QTzmrZ7VKjcCAubslohTfB
awc2acohTSHuMYkz2QdLkOGx6JsHHchecITJMBLObyFhn6S8yAvYk7DX38ed4rJp
xz38s6z7o8uc5vFDAsKDzvvMhJEdPYbg3MywIHiCppMpxlRjyea53BCQaUJ4iVHE
CdU2I3zoAVZFVDDN1hFTu61wJ0AqHwUmxeIBhMis/NVbKmNwCNYXfpQ4cvAvS7qx
lPnrCGfUQYP0q1byHiROlzCm6IaXeTP8tZa0y+N+VawDvvcCvc81hy+2FwqlG/Ce
ahuIN7HWAQpQuXyVmf1eic4SMc6aKfpVtuC/TdpidAvW65330zHKlW4HMfMNp4Qd
wAZilfsIwbSthuKMVjQP+bBn3FNVIUirdraR0A+7LqQrAo3pmnuSbz+4M6A5W6Ba
ZCeLjcP+6SP9zLISDaZ04TwajCm86IbHPfA7LKeOsRS0k20g+MKfGQTO5k5kYzhk
Bg6qNcOuA8lNBkwBnP9AKl3b0E1DzH8p2rgkMMXZOyeE2o5ZicdnhacTJvzcN0Oh
tyhVZryd7I/26djW04qLfHUt072JENecSyaVEzA4LVA7X5PkzfKJHUcxDxEZUOnH
sOGE9HDzundSxsjB2/hcJKrarLiOObbOwciW/TmVAzXaiYJPhmw/UI7/QnYbPXcZ
Vecu6aqAPYyOyjhy5OoAJuzX7zX0k/wenWTUioK34+N3lASQQ3ODmm14CcvROQJz
isF3zObMYQeghSSj3JjWkgsCl60xa8J55AxMIeRACKYvMOvKRDKpLbY5vIb910TV
obLZcFAAzmsbpsVZwJuIcNlP8s21PCs7BZS4bbmFxaN8XzMqWQIyxgYdy/EkXy0b
6t9V64aqpC2E5qTtLpEG+GRg5yG1H/AjoOKjbpjz988ygRTILfUAVaiWHWpthePg
+HGt80lpspiK9zi5F3a5Vhl/6GnmiJF3chmZmBdwmKC2F8bnyTClU82fc9vFs/ht
YBWQ3EyRzlMvTDA/wUZfuH+vgOqXiRZ3VN9tKj6/EyCRmB+fYloukZHbwH3csRAQ
GNU4eLzZIiLugxedB4g13Qva2grjUOa6/ZwbzTIkU5tqGsyomlmTwozQjmQBF2eY
xKVj16Fnu2wATdHL3a4OMs4rS8GB4lbCUY/u/qZCZSU3VDl/HJ9n9+Nhxir94tYX
9BxEOSILv0Iud5A3tQ5W5WQNsE7EWrxlIRS6eeDY5AG7sl4shnIxK8oMjHCQqSZd
ghu6Z9a3zZw9U+zjrKSgcrWd9VzcoASxnmXAfoM+LBAW3raMe6GM5gqRThql1zKv
oka0ah8UPRZW0LFDoCT+wew/ghiM9agl6i6xi1NQTcSDLjWmbeWLPUDIcKdO7oDc
0W5JAkugrH/TVl5MJSMOiBESGF/mfKiGm8nM+QGInRfl6uKKCzpbnOl5e4nOBWo2
TboD01HtfJ4Vfua6Uz9pcCFrT7fbFY0F9jOnX3wlsyDL2lJL+3c6QkN20lpnfmYP
9K7yUYzEj0TLk/BXL16lP3fNMu8lg75gVcjYxAQG3jWwYb4ZSTxpvJK7AdEMDkYD
wL2vQ0wJjYHZVP+10hG58aphFEoIkl+EfXr2aUlXvCSODJULSRiW7veVn1xdFZoC
YllIS7CrV6aJg64Tv1Mbe1qfTlbxXs9Epnta5VbFqPZtkkBbjlPwq81vt4YANy50
vF1CN3vbOawh3TRtRMPk1EtcC07FbCkco1lisGX7206zG4VRYQalVE0FCDuAZ4YX
ShbunjQX7Cqy90+JpnwTtYm+gFdeVyPAy/pnvMHJOd/z3IjiCB+TF4uI+BiXfPkR
tbPVYuSAutpuY2zUOAfTlpGFHpVZT8ftTT/5l8n+IkUktc3FUnW95CMyEbwqDP08
cKWzxNYjXwz4x7v5inlXLRXLFyY6bge3PCG/ABighsX8Isl8T88ocpfL6jXs4+/L
ZNnIJ3rLIaxD+12Rtlha07Re67enwsRpqxSXVyWuc3rOlLTPymRJbmC9dytq5iF0
6yTFq5oZHBBQBNfjUEI5XJWCKD8sLfgkJGTTfuTlRimFL2X41hxZ1QAUiV7RZJU/
UgHp8ozBV02zhyClNcl+/aQ1FfVmEI8Iwsmg6EB8haJHdOmuYJFc6WlDgWtNBcGz
KTj1bvT7arO+nTrR/P+I7FB+VM+Vlb0CMxqQ9gF9Wni/ORq0IbE5XP/ySQ8jDyMk
FOFVKEhp2viQShi2g2hhsjXiGpH8nn2dSDbw3mzoaPLZmWLGORiHKgp6EONKI3/A
EA9BYjCwNeTlYM/g9jCDWKwsC6WW3mqL6uOR1OPWq8tIsckdXtx7qlRTlDE9Bbkl
b6ebrn0mZW447x5v4lfsIdcxXL3shfNQ7VrEnUWlXJAdrw3i0eaB38lgC0YASNRs
YFfl4DGor1bKADmTnpNyLdDMuBb2vAH2199iAGZI10nVkQLQe3ryKvE/rzizK9/m
8F3jPGVCb5qJmipiZsAYP2hvswoVFHfZLQ5zT8mxX9g=
`pragma protect end_protected
