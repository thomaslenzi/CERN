// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NDfY0KqLP284QO9bhnELb7V//Sdmb8mSSSb5/LJV8cFshxoyzylvrJgTrU0KHqdr
EoVSGm7uLpYtwIy3PpswgoNBWpUmEVBnNkgffxqRjaxQIJFXO8QOJC+B8xBw3XdX
YAOLgpHn+2qrnzmLjDrwSQzc1Xaz2YMu7Z8sz4aK/Og=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10240)
zLT+MvnW1rgYOhk8elgk8fELu6E2yrJ7HlchlOXJ7q16YSV3EY4jss7zT5+Kwztd
eh1TQTA0s6LLYiKIr/+3z1VCJQRFrtI8mjRNyE5ca35OGgMfLTA2ujMpg5bBlEPV
zRgeOv+lSZVmuggI375EkGN6qCCQen2habpD7eEr4OW/JT+GgQJOv+F9Q37lppNH
UmGix2T51XRIsVKPumEfRPeaXz7cw9V7EAoKQWiccRtL79X5N6uROg9qH9a0PnuO
/oYn4L/vS5xQgVs0lky+gbeFwdAhL8BVG7OiM4oBVr4C+ArNRLL0gsAQsnRBrgus
nc+hWz3+VWQY5MYuxK1R3R3MLN5ywhqrR8We+2d1n6svr6oK8VFXZJnnqT2KQMDh
WjyYMdXOtu07o/lNEDu0ZRY0Pkv8OtQh4MYW0XPn4wtvxUixyqlRCU+kXQYnhcag
pjZ/pbXOeyIFwgcLZYU6asqKg2JaW2PF7WyMR4QIun2NXM5kvehCNwzje4Cq6Q8q
ZoMVLAahvquS509SrVMv0I7z2zqVyGfblKkl18XNbG7Z9jgjE4XZ6jzALmAORjSn
82KKlSz/jXbn0GMJyhRU/SbL1/c1pIaPgwKjXwyqP+8ZRADquZliZ3x976DNrRk9
xsMQMajEnkOPuHZGfdpAmL7sTPI74K3gqRsxiwYfCr49aSEIrRZqh7g9ANhLAa9u
saqzg1yu7xsPV7TE8tEnSywZ18koqJzrRHzZmnCzv/ETyqZc/z9WaOIa2XgcTec4
5ZhWPCwdzdGOPYPFzDBG8QepTcxW0++4mOq07LAbiuEr10jp6ezhY9xw/fxyaxcz
8bexfPnjlXLdYcRGZS4a6grSFTSJKghYaqCSB1WCtThnrNjI4p9le5pCs6Zo14gh
mgDtlVNzWHchBy+d4MK9oDakyr3GshzWv9x79uqETSfapebYQk65nyxziFm6wojc
Ot9PNEXgBZbUgjoJcNqVP1V5NzuQzC30OCdtxgMnKL2DXfTesR+SLhC3T/HPf++X
dcWwQrjkGIvsGynfocz1jmYiWMUykiC783baMYqkntIXkE0i3hqtSS3pDSquTLG+
WsfTrFHOVc8UjKfag3770S+adDoHVgwOV53AxfhzXiK3iRvex9jBv46Qgc20+JUv
zBgReVc6+bbQ5DcqsSMUYm2XJtXPAdRGFf8JQCbiKOt7Tuw03XZ4mkFSiQ6gtEEW
JPqv4YBNxsZvMZllOy1/Gi+iwtbOKDQPY6MM4T8nvRqauJMlnfcFWXwwV4sQP/Wn
uuthF0qLhpoAS3nBqQXVQr2qX1TG7IpSsnedXf4BYs+JXq0ndYp2UVNVoGE2deUi
GZvEINmRsf7ItD1DK1c/jQtoCi3DEAIYOCsDCPM4wsyllNuLunudhMinh3QlqSfO
o9Ye7kJUw2sHNh7pyDBAvZF4J75bx83i8M2wtRWkC2p1agHkbHdLQcTrTlFc7eHP
O2ULsQ6Xuv2Tx+YMGccKF2eln4y/LdrlQctLKoeVUdmA+UPzokGATd3cU6r/wmnJ
r5GpPPVk+Fm1r5mC5yi54L15/zAS18FVMg+6v21dZNLQRqg4x/QGFI+YOkf90bKZ
15b786BODFCV0uimBEvo/0Yc9mUNtxnJMai/KnqaIkM/fa2lU6iEyqP1+OHMxr/E
Xj3Snma1ELY+ekdHM4Dya5ROckzdrMPGWVdDVCxK8c+8zhWo3UgUz6juIdseGhvP
cCt5K+nb7nATf0Bp64sXqRm7hk8vuWFTkTHbKnU+C52DtVS8fSg9+eRBVf03nwZQ
oWyf2d1tM536qrt08OR9+aUGiG8wNK7vCy6GZY6jNmzC/dTZYrzP90wgN41HsXnL
WChNM/SdMPperLc8ZEeb/+G8NiIbS6TFyibviA52n+34CRW6kFuL2KV8fALrRxI9
3nlcQcJtl4t4J2gjnlaC4souIweIcdCF/jkbRg47xXrs9yHO+kO1wh3nMsxOW4FP
hP1FNNLdZ7iUSreLWRc+FUdeGRfpGurtsgfaD6c2R3/wsQAp8tKi9pLnJfiER5vt
gqkXCedmmz3jNxk9V+bLWMyw+1rKKrI92NX5xX6x3lDck1CbOTdCEDPY9AGVDGIq
Wy0XQSt1sCjYlAigsuGqJc3HJlf1+PCKL2aA/Gc9E08s7/e44ly8sU0KxR/49p9y
tvlIxFMhD0TOcaWBzO0rxTywak1BXf1JEMFmCRdGij7ep3nb+JGaXiQ7DfhowVea
Xz5BhWyVFGpQvoHoKzr4V+InivjFZaDJqckBMieZsvsJHV8S+GZqoYPGi9OEjJF3
saKniVQuP8VE9rqcmeZjoMxYhDLP8qPJydmtPehHNi17QVFfvMygzxmKFOZwIAcK
ngqcx8BJFP4kQ0g/AHT5uom8HOajGTTctFK1BEuwOfJ7XJ4SrHR90NfvSo64J7ml
gSZhWhklhY/3Q+hr3zu7aQGyV8Xst/MvQrZO9Um7MZ+ZY/l/2/3kxHpYKykePB4u
zDhx4geVtBPV1xZoo7AZrEuWGEQmubmgcSKhUrPp1yEW3eKRnSoADQj/REPcCEYl
M11uR1/FQklTfhfhWIM89KfMDvW0L0iMiybIbHhFfsP0DA9ETbHnRpIYCrftl2pd
fk1Cn4dGDdYXKBzkAUWCw3Q+C9VlWINPlbGPk+dsfsbM2HMTaM1Md06CNCkbYIs5
XjIV9XTWXRgO2moo5X9AqkFSUtPJ9D8zUbudY4aPrZDMhVWR2xypbQaJqLdLvdl/
G0tYFZgQ28DuHdOM1IVGrGRXlu7wA71l5/zLWWEEuQ85eHTYiM0Hw/6yvyJlOVuZ
wQVWjCxryEJx6FkyAc6JQNRtwQJ56WERVMHGHaKHXQC4nVuOU4+GuMi0bTtzqttO
4bmoVbmw2sZeLo2YoMNiPNq0bRg/bU2kVqe6RqDPSMM/dmeWNv4qUGPbj0PpaJ2L
T5DZk1XRB2XQu02K4tuakGkjReijCx7eQRFk73dMiqPIQrvJdmaTcqZ3lyfMB3AK
rDsKV5Znmv78Q6Ve+6e5C4CHRTVLBRRrQ2o9Brk7eIEnWf3jRYUN6l5CbeBX8YAr
52XtTYFBsL6+vaFkZ+H3Tz3YbRQ9wtle2oIn5l7TEFL6ZV+UPPms8ZIXCB+ZyQuP
IrDra5FGBoHUuBoMNmIhxrs7V4I6vG9qzc0iCaCw6btdER3bGHp1KtNmFlfaz/Ob
y1DFSrPVE5uae7BC6MrUoUDaKPz8bPRs2hjHBBy+c44v7hmmORDb4e8sA+Tlaewc
AGT1hrdd/T8IE2z7p3VeeSHlE95DP1n/7/mVlyp7zwaHeyMLr/2WQ9XFXn/PgIx8
sFC7niFOT4EPMZEGGA0iW9gbEaTzshPq/RDtudKx0kTiGJ4B3k4F/xS5dYDsxwWu
bNhx85jgW7B1JZQqn33A4TZqm1RSpt8lUT5cNDYH1o7x9iI+AnuUshkNU6hizR04
WH2h+B0Al0ZNOZDo/hDiFY8XQOa9UnppDNKkfPCA6r+pcR1Eui2d/BFHWC70Dhc4
3j6lQsitT/vHidEZYEFdelSC4sD1u+S1gWSZy84869/4Lrf3/IOq+X6/WhgyvXoN
rHguKWXggWOtzg9OrWhHJOz/g+1+frLHp+eKoCCGU0j6vW9cQ0PdFij92qCrUypJ
GQyIM6onc95Af1c2UfCFxE6PFB9G496y2m2ig9kT9srC/jBDA/R8xRXfroRACkWc
DI86ZtuHzX+xFMMBDMgicjI6PJKR5KUkYeSctwbz+OB6Rreh7RZ/LQw6r5LHIWG1
WCeOJEH8q/eGM8QHc+4xVHtPscRAQkCGwdqgsQzWHxC9DNp7oscbullmeUkW4nA+
V7qZLr3pzOpaIqGKWv0L9PUf8w6cB47D9wl7OiQyOI0T0ZCxNnx5rIwQcUuf8RHn
0xh/mZF2eoI6sNYub7XJ+NZmUfcp17dg8llvuM1i+5/uqlxsdytZM0/ed4msLHox
6KZXKMpRaCnJALSC1GcfrA/T9DfSCViWMmZBPxo/xRJITS5Ql6gUWmn+etkY7iUS
xsHCmEL6qxoNcZW9v7N6SqoTBNAqhW+chkR7tii04Jr2dg1Y8GvcOpWrB4Xmb1MH
oLDRVagCzBJPlgS8mLt9tDEs2M09n+/WNjsGbUvUtcy7DpMQAbqzsvVFD4hTWf+g
3i+8aiBPQEkk51rgoag/dqSE4aagixUtfUbhddgnxIi6eXaar8JrpEtSQaMM7R1T
XB5KdeXJsj0BNFxDuf1tvaVfh5523yuN7VgvSkE6rO5dzbWValnqEiLKYGGtvCYm
x8E29cr6aUHGaakRD5Qe94DzS0Niq276oYmG4SxLRdJKMIzsONTonUvwaVSmzpO/
nk36hwF6SgDkd5/Wr4hut1Mf+da9nMEOzauN8dqsQJ7p1+RyB9xoJbbNCkpB3NE4
nCptU2S63LUE/wZXJjIlODJjyqyfFHIzMkcDfcB0+iOSYsbWxfoo59Bfns9mfcqc
EJ5ANKKNNwZWgcSleMEnSUYkpP2aC6JM2Ax55CO1imkWOpq5zp5A8k+f0j46pBgG
6seDyRvuxhOubzJoTte4V4+lxr//gcbnauMl6h5sN0O7dsuA+Nf4rJ+fm8Y1NNNj
GQyRcszfPRIEP5F2nvj+YuwQ8EvzSLWr74Iqk7Q5BWzxIc5YsRl6FDItLn/YTujb
H+xWn/kPCSuoWGy4axqINfTWxpbbi+p5+g24R177GyLL8Wbps4WigSV0HzGM65PF
DpvVr+AS1juFm53ZHEGFwA4h6AKiB07xowqcUr9NODGV91Hgznh0e9PoWDuUajxP
2plkuLGCQpYoaTYNFYPtudE3Vx5ynrNWng31kJVcCLmyAbo2B3y4OiEP5V1CUgdm
0TQRLHH8MTq7I2qlwqB4L9FSHwvsFQsM7ffw5EuYLXu+tt3EqGa8ARBQVuXk6dJ1
Rn7rlre4iutLs51pg6lvE6Mq+STBwm7s3T1gdyVQxUTjg3mTj86RmNqqATSGZeH0
OkgGQU+oeqL03HVbTxBx7zLhn4lAzN8mnehi8iyZHlCpZRbNOe5dISZ+aocND1PS
Bw81nAvXZf0vMt4pALv/P75qCHq4zdYJgRxGbOh1JC/bGNTM9qeSwpMZ9KOHi4Ao
YNfho1O+W+hJOmtZ2wdWgI5NihvhaAEApKqaBcNtbzzdyA1w+Sudh/Ton8KOgwZL
WhqZx9YXVuEZrs4KB90ENOGuQFuJJKCnC9yx9uNjQDu90w0mzDrTB67KlhtJE+D7
MaBUj6fwelqM3EQ7rsgdwLeRmO/0ffMi8oRvfW7SKFovHiivSkEj+PiysdZTmAj8
7y2g+OW87B8rmeEE3OcHEXdkb3DEtffARrWd9Vp0yWvD+nQ7i1nt6eL+5xH2VTG2
nCB3MXG7qpNF3u2+tgLDBP4A9/q7neEe9LfUVhol3q7nRZd6WvvyFDbpic6xNt9b
Y9cMEM7dWzMCVSTTMV52RphS65ugLAUNc/+pbCrmt3ZJpjakvXPfQCyIYuQnh6UM
4e+grLCyEA4AQESwWveMMkCRIYAUBYxO2ddEBH+j4AaqaylgGkscvJHjbjs3QsEN
v8P6BzpoiYB9Djm+ylwh4CiWC1D1O9kpWoNZNl5jEWzRjR70QL0HBi2QPkVtDiWw
/gAIzNVn4/54gr9fYwV0qEin56FgdYE62M9nK/OOjwJ4Cykehb0FpPVyNIaCH9Cq
cujV6Romorr1y63tr1cl4cG1C0nza+WtY+4+5Xy1SVcjD8bS3vZ6RmUP1xLglnXt
6SiLe1xBl9tnfMwY5ULoi5ikN+ertFpltVYAcq3LdyTiWu3qYNOhUjwCbCgvNQno
C8zuet6CAabt206BTaDg+10m3rGWlSvdaib8CaMeMLTZaVV9ImN4mwFVgKZ3ZAAH
WEmyrP4xwsKVjZNvtDbVg3ge3iiVtdSeVSYXQXhHxYbBUSPKfYGu6e1xL/XwRvmJ
4wu2Hoom+a70aLvK+1vKKveiZxxyA4MLgTuczdbfwtOvg1eKLR3+fkjDgMNjyiZV
djVQnVGgSbZcmXDzBhr8+ASfXHkQHsbSe1CUZxpMnbSdDWOgnUe5HRsNygrQfm3b
TFQdsT6mukU8O8Bu+UxZpuc704zaM24mwMztV5M9zCvsA3knxgtQAFLXpN6IKHbY
Dq5LxqZ6Lh+jixgT9FPTX7FBiZZbaEWhBPaXhELqiZFpremHn4QrPSEwEMGUdxsD
jxOmygPPrPlOeAu5a9bbDVYSHmcpB09XhZp1Cl/39tOxyWtTPFyr1soO4DSqKISF
QZcK3xiARsqH/ym8zHKkHZZ4ioNsesVdYsv8XRKOh0aqmXz9SmtElGA/lNIqGXka
q2TIVi6eQ8qakIu5TIM8720gV9mXIOoUYLhKzqjyse9cG8qBRcHu1rRPaRFtyyKQ
kJxJEHdFSgyJ4lghh1+Xw+ZIJunwCAQC/MKhICs5g5ppO35OLN7tGjkf+A3gnrQK
OWvH4z1Bd9Lf57i8t7+9aLOfi5J+81fEAuf3jsIdgs3mCesqxM8hc9XHHYKSS2NG
68ExpM22GxL/vg0+gwBmjg4kMMRbSyTXQIayo7UCTsJTqvrIwbKQ7YJtfzcg7BaA
6EwR9eMcfL+QXZRrFCIxdOy2fv1NVyngLvEAR2umUc38zRRyOYZVEmVWLzZvb5Ts
5RixybZfaTuTbOnhYDCZNDmlZBu4BA5Vz+Lr2d7vFuvTcfE+qjlwXxdj96a3yLIR
d98rjsgPloQtr4Zi/clultiLjVbbNEy+uwdAxK3n8uqxp0uInAJ3Hdezy8FR+g/m
C5NkPcROh55KfrnepoHhNktGb8unaY2Qb14vAFrCv/MBffAJ2pEG893JpoNC09EB
QD06CCZ39SINJTNIlHVqPEYoLLupQgCHHBk5fFGtNBAAOtkkatiDc8xFHwdEDVxR
F3ODtbsJ2Yec8zPallarH8GhIgIBcz3AZqNAB7ouCQyqA4TB2ItLos/xtTkApul9
SHLH7jjKnQkM/Ou+sgXGFCUctAjFpxRf5mhzi24OIsvIH+Q97j38vi9IaKsI9mSe
KFIYZASeEcxfj8g+NMSORv4UBRI6FUhFUBzOKjBPq32aYj9i+hC1OdZh3CUPxmn7
I3C0QVs6tB/8UUZ/8GP+nxhHr1pyWpk+wjvAZSGi6dSV5VXye5r83qnkYXl1iBV0
w2L+Cj3lGpyL6WfvtMsbwAhIMS86jPaCIUgd1kKjlo745Z+H43zaH9juYX2TQpGC
rhmLExcXdHtV8z3sB6ND9YffQDAC2VIjuhC47GfXwzOfIHB7vk29x7JRIWIwP8fj
8RA23dVbwY8XCkFVdg/p8Fqk4u2JOqEWAtdKgtTSINbtsuNznAxcixOk5EiJi+gk
h/eyyaL78rivSyJ8u2GzEmKeRN279M9v6wSsyX977Oq9c0d4wxYkRvRVO+RK0ALq
vK5lTw6q3kzH6nJh5gvfC3VvGZC38Al6r80Fw4GSfv5mMqiv50iqBbKjWkSrfmkZ
3yyc+jSAsOD0JIH82jWiqM1cPNWtcCszbEGr38zy4gPrfHMECQB8PSprGmOfKjyI
KproldWuJexEgdW1ToRVAmvgArvzgk+E8BvNhraUctqAlBpZBx22eEPS27njgBSF
dJnHo7cxXlmyUr4mK5dz72hfzFer+wmZNQrcfYvYKIvex/eVGu51hBId8sg2fZU3
y28e1lL7Fr4M1S6O4+nh+A92rst25kJSPWNcdbo4ObBCx3+Zp3WuGUE94NZyUoUe
Tg77YBTLFk9Sty31opxfLWutELafv2FMl+Som2wwWg2gTIOWT+I0TpcmJQWTLRx5
JHMcSY7C5tNmoxIbT5p3cuXUoT8qYJ9UWnYHE3aYU7Gt9G2q9zGq4flhuHwjTHDr
TZLtRCfkv/vpWwQy14/6XEelJp8PvJ1yeqy6m7Jti9z0JYiAMGmwd2YXSbb4fNl6
OoaHjMpOPcA90FSSGv2VmK24CJwsLhgph+QL5TbxP74PZ7w4V0h+OucFgGB0Bx6F
3OuOtJO2FB9OOlm9PZRps2xrIt8c3k3JUmSl22BbdxKLN0Q/t/YoC1E2aTfiWYxQ
AS7rj13+OqBqwIT326zqlg6C8+E2jxS6b9pzYWsKWmZNhMi8OoPFEynnHsWwQJ87
Ma3yowrD0/Y/jl8X86xDF8oUncKGT6RmHSWOqqejuEKk4fW5goqKovxA765Z8PlE
vUo0eSekQrrHHs/o7PKnfwqjbIfm75+cuSqrHYFW3THKQQdO98KrnS8EV30nmFUk
nGpmzGz5wiEI1yOAn034A4vws82WSDZQiaJvxWnpivh4Yq8AHzOtoUgfeLqKBS0M
cGrmtU0UpiUwttxPtVc1uKr+DCKUm/6qdayJ8NZtivINoVo8Kd0/Q8+kW62LD7Sd
54d9xKsvoywrNVFp7+XGqhVp+pBj+4VnVcGWjaOGtYscIE5+djziL4e5oxkTFq/L
EuzRwi1kIrkzmH9MRkogtTcYOaHFT+2OVuc+6cQwc4yDSiBZg524Ud9Ys93HB+s1
+GMEOELZNwI0Bex9Ut9xlBfgT4wGsTZp3Or+kzOzGNpand9+uU4q3+7icrf+YMay
UV7k/liRNVjXJEZHIqS0JX618vyZhdqSF1fMmCn+aneunqnS7KSOysgC1k1ECgoy
8gcgQ5Z4+lRCwj0zRefxxXHbADdTcuAV9adcFozu9UmNBRQOVDwFuSW7lVtKroGb
jCacNcmQ41dR/Mdu3/Uk2admDj4y8JG8cbGsKWKfZ/Nc/Sv4yWBerhAZMdqpUvhD
qpR1FZGM1oCKfRtKGq1x7HH72bE4w8ULBc6avX4dr8kHEY0Y+RJ5pdN2saQBZvNW
L8fz6FZRJ39AUwqlmrl76rwMsmXLTxfFhZ+hPi68/sGMr18/2AQ9/nZf+Aj5UnWU
ORRlCoIlSfwVPACEqODY97LjywaERUqTtSKLpQbMw88BWMBE93tN+X24WD9C8FDf
0rhvDAQpBkJw53obPqOAgHSnGoOf1vck+wohWrm2AqHhZ3lhbX1MtbblnS1Zscv2
PRkiS5K3wY03sBWE5dC1xa3IZWZ3hGws0LLGgXILAQMHDPeJ7whgnz9sZ2D/APxH
VahU/UK22GbNiKBTynPdak+UN7oiaSUuPn7UzubxrD5zShpxj+h9/0ca233vJ26K
7SKUw00INyq0+jGA5RSoMUFmhSW3sd7RwkRzq8JmrSyu+UntzIOcT8u11DoBu2X3
Kn/7YG7eeVrE0ZbNwYv4qeqvITvkQXycdDuy/Op7OptVIsEC4et7TQjcMzhpfj11
jL1eL9pOsRlRgKw9ieZDDRgFT6zoNpqms5I1p6EwmUpSl+x1+SdUMqTG/B6Aehv0
XSW9Ji08pbgbtONLidHXTMB5IMpKVEX5D1qHG6PteOOvBPUWc+fKboKW2KbPMtCJ
umI+jr7DPMb2zmu2lzt2P+a8DhszHuJD96mFfVzET3IvZXV5YP3VXIb4/LoyI0Ae
0KfgkjsfUI/wK+bD/hNaGxvWxDZVYCq5yJ7opp1lhs7aPT4W0ubSHwjAiIKlnEX+
PC49b7/L8Lr4d2cvSQeaazJ3w94gqDpl2lPamrkybv1PBrOHouOWzr0Ym6UiH9Gu
8H8zzRQTV+lBFZfyS1GfF9vKYHJuqMmFUDnbljOu8OXy+Vzv9R2UBhPfbSTTZvxh
0pXlqpyX6NLSSgFmd/5G/JdKe1FgyL82IkV40SIOsv0EsGIrt77ltN95PThI1YBj
ZVimKPUM3kPJWYDugkU61gHYr+tN1wYxezDaK0wOk3y1Q7z3INmD10L5dk/Am6wY
0HdO4i7OUL3P51QaXGj36NiWlcdjk0I7Rx3+r6VPuYA0D5a1a9z7aRMb9HjCPpoG
usIjYS+9/5TEYlXYLkv5FbxVynagEp1cZFWmUVD1daSA+/GoJnwC1IXGvBkErklz
hByD307Cmk7jH4VgTyLq1QXF4p8nSKMal1tBSZjDD74cdDK//UpkalreeSbRgB9j
49l71LrGwkkv7a/VcpAk0mTInQZHFkfl7FHvWC6tHcyWKsHsqgcv1jtWrKxG9sYW
eIlS2eXNQgzVRPaaIPWNesqrJIzuiTNaMi8dD1FpEZXNhbkmxy6/5RIRTwjU98tU
19EXGrRs9xLxXst/eYraHYQXGhHwjrwXlTRQuoTpbAaKrz99zcDiNuuUAyY3wJYU
1V/fn5MoNV+v6mMPby6y6qAp4IMhCTWiMfS2snEYOR4XFEesV+tMacc4lMUeIZvW
WBLvA+pbCFFUXtI3GwENTEwHyUE/ghTvTsBtnV+bb4uvd1fYEnJXUBeF8lu0wUqH
+JbuwO50+Bvs3kOFdyysVRDRtA24I1bJYoCqNRCaz1r5V4P2Ai5OMb0lye+RjLot
ZItjZjNtewWtbOwiE7VFq43Xh6uOQxT1i5qdjLDRYjApbTWKN7J1Eb1coyZFAmqD
Lo5YbUWZXVI8Lt5aZtYguaRyLLp5O3RcjApHKUVYBjARxe3Yg0vCH+nP8v/RwO1X
vcf7kRBJa4JaQUygbt/ojY48Km9F5PjuI1/4s5O8NkDMOCpHFxvzXhzeXfPM8gB9
ptiHnblo3CcolTayCO6JZbeKKnpbklDD6GG/mEpCDyG6qqbuFJl85ZY/r9zDg4kV
TVqfoGmq/CRiIzYIv/p61l7ABFihSU9Fq7b98ulbduOjz+SaeB4wWQReVJwI0bnK
8jZcdsupW13i9Ga0FthrSVGHGZNKvmrmdi+yfhj+hC8X6QPu8i+mg5nwSYMKsNnY
O8rsQ+UHGyahgt5IFoY3R2iy0lMV5Gr9lg8mk8ktHVZS19kbUu8EvEz/xANKI7Ru
oHwQV2OASS2d0NZfOkpjhTKvT31w38RJ3QCc6o61179MCf6tUn5Is2Tz5VFaIWIr
YTHQEcgvQWyRZ3TGKYdGzhOwF/UFIbQRZOE1RZMXbfE6V3ZCHS0HtwXu843HH5o/
Na+SUXW2lntE4F7caqJ7y11vlzfjSZ/4nk2x8fS3GEUS/L5wK1p/0reGZuFzt6iO
C2bhquENnSMSeoZe3SBxK+RYsnE7tdmTayyvv12xtLhyP52lVc4kfIA8Ottq8hLC
0aeAkCAu1OgdZLl37kEP9NkTETIBH837YSv8TCLZPh13oiqa5NzNKB3Bk6rRGm3N
fYUjZ6LejM38sN+BONwFQU1FeFN2mKMWK48G4z5aFNuAiy2Xx5L/kM2IiO3dp0Kb
Uisu0Ad7jxrS6BVLM4B+x4XFECI2sS5Xu1fqs7L6d4SfesoTXXUHRz8aCEfd1zn7
28keBVLVk4BfDzSIwLVRZjw0LEkr1I0ynWME8ML293c7k1NPzYGyHm7hiEmrwRJx
tYBUpE5Ig/Z02csz/X7Zo/D/yKplo4pdcwB6Y1LNBI5BTsjVns2s2QyPAhsHU64F
1ib588lDbi3NKRzTDHbUMBUi+MlM1/MXBMOXuUvCbIPWKJZFoe8+C5ZttIJ4hvqK
+yKC1bL0NlS8mNeoktRMpzxGls7TO8VQ5+vUgTP1/CyKCbT7/ckIunXDG+LVAvsc
cYXQKWEvdKwO64p8+3O4WN8iW3hKrfL81w7doYfLaxLSi4Gfe8mUW1ovL+b0UUyK
ozrpCnvyhYA2eQnPZrWp/dIGP28hV+EjxDLHF48qD+l1DYobLYIKqq4bvhkn5rDK
rupWmG7zfdpm+tjz3O28zolgJ0tEWXBIzoXddSBw/yt62tMIjoIfShB/48Bn5ETf
O8BgK2nEDK4b7JlCKQEdnNYqPHDg4wpwU34UWWjrRFORLG/ZZG9MG8TtlwKtZ97t
rsZ/5lQEkOvNzhEpV9BOk5Hkitd1dyRMdd0WB087m/azrMwYLgBDiertNkNCF3E/
mXNR7v7qFN5NMWovXL5ItEKPX2xMIPFsf9aRYbW2tQcFl4++lct8RWP3F5Z8uU6e
4/J5blfVS7dvKIKToUbLwpwDfxPR5luXZ6QckKT9r+6+OP1k0YvGZSfAAx8UArUj
t2r0R0ir9ekrNS2LTwqVQyO/Sv7piJfpJ28q8MZEWPDie0mOrqWHt1ImZOTgwwgB
JS81M1R9nuZSNyTO/rvu9sE/xqw5xrMq60314lAr9OzX1toJOC+OHZX1N6qg9vpq
kKY6UEsk6vvQygwNqGgMX8MTlFG3GNN5bs74sXsiQKfEH2GUHZpsis2mMfx3cwE5
QlHoDIV6tqnqatGqgS2RJdLJfUhIDmJaoe9jghZP9DhBsl370O6x0/+CWCaVvC+f
O+n/vkWY/VO+H/Wf1KBGvIVmO5pFkODWNy0k8t2Sr+a6zlmGDXefrvaUxWVE0gmh
6028ALIRKSrkHxgUM2S6W7jr13/hoRKgk5VinuWg6tFIclEKza+FvkVEUqmngjkI
C3GiAfdYb7IYIZIJCbvtsU2HhCgQVTkkSrNRZPoCUn8vWsrNep2K6xvJiyN6PLNs
sxsXy8RLAf7oyPk4rYdXmfIo9+/HsHHslJvp3Kjdl6xFLLdDuvoY9NQOTjSL62tn
4FFyPwcEcoakUDQdmzOpAkG0/cwARoXAQ7aBHKMDrs2iwDsUTJHifjA6HBE1P4BC
tByw04c8wzJf3+BTWqWh1a6QFQ/EQxLBdcX+XiDwZqIz7xqBn3sI8ZI2fiqugsJ6
+PA6vj9UFq+O+9Z7uIa2AlYxIXzuO858+0cDEeNX6SBA/T5AbwhhDixapeF5fDPO
JIMt+5jo4lOxAxMEAmsC2Md+BswTZ/+mRVEXceV58q1w9nv5ykTtCmyvBG/XABXR
hZT4s5zlv2wmGE13U3COdbMvOY4XCKZA4fepK4Sv0pA3YTtBTzJnroQAxroZdrF6
99wdLwYKBBPstj9NO0n1r/PExPwjz46i8NsHebILyJA1F2UOORryx1lDYHBqxYek
s947LeP6rrZ5NZq6Um12npps/q0+h8Z8k3iA3CJTkbWsgkXSKK8xuA+C3egSrAir
thrROMa3QTRD2C9cs6V4Ge7IhT4sY9Q/aoAZKRyU8trAt63Dd9gXAlr62vPwQVpT
eHnsgA8ljbeeqNEbrJ/OMwmf/f/UPRP1tmhYw185HGIEJOqQvlsJSr7KR2bIHJp+
sF2TC+RkvIXp1TlVuJPZT9FXaoKZVZRyS7Cal2T6p6iANIG4le+pUJbUgQho/ZyR
XtlxaFA6OAmUr+af0x3NgMa02FJc04Im3QUozCWqSGZCqDBKZBRRrdPOVlBY0u8x
0XCYJwSYvlX7nFhGSuxOKg6e9QV11rW3PBZNg/nDtsWKxWBixAfba+zA3gOWWZQF
0ZbKkuwfhR4nUHwnXd2lxItrt231A0YXC5cHVGaWrutIMzVvyAJqH8ZqmWxQE8bv
BHpYaH5L5WtpUkWM2+6MKd9jtFfoztyBNWFfKc88D+em9mu3aIugQeQYwyUYoRnh
qZV7J53JbSjcvbRcSjfvMRqVIuDfzhDeCH2mcQn5za7hKv7bbrHPR/QYYQuXSc4o
tCXlDxK7L46+3LGdw1WUT9fbHSoQd7H//R1zVUgZO2CHuh4GGDWOnOEkGY02h3sy
4UwpCYcndsoWjUrcCbMwOr3ahlLjjlNdSE37uHlLShA2xutknOe8ppyeacP/OOyB
r9Jk1wx884S3d2HSixcxlA1wEWaaj7YblPi2LwvxmI4etO4aFwlHWWI77YYMT4ai
JzWnyrOZRnX1HhxxhAz9kg==
`pragma protect end_protected
