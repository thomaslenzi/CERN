library ieee;
use ieee.std_logic_1164.all;

entity adc is
end adc;

-- ADS1015

architecture behavioral of adc is

begin


end behavioral;

