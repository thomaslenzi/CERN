// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WEocctn16CWsJrH8Yje0IgO359HziaUiiBmnWrdWT91aKz+slYPAS5VKSYSK5vx8
gJDfeNhFCHfD6TCb6AsGVaiPhnJD1qzs8iBodOpj1XEuM2C7sHXeHqdQSzKPBeow
/ANn5+ohllnTQtALconpMnFw3ClN/m0iHzSzAB29iqg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 105120)
gKT3LMKoKmurqtv9ykhDpMKvpiL+EXVZC1EJH+5UDcrZodo1ZsARoiCnLr+x/4of
9vMywWCuSrJ84Dk+we7a+ktapxcAxbhvLgeyTDW1Xb+XBwy0GJneOyLy1hh76zAx
lcaK4cZh4TPn/0WI831P/uBlxSwA61rVup5gs6RWq83oKINtcmFPUvZ1TOGnU8Hg
MqmZPJMg2UJjyo5OMryt1XPIB6tAG97KyrcNrw/cF1V8oDK7ZjheES/pdaBTuWOQ
P9KmxbRpPyUwZf5CokWybJJ2KKq5jjg8dSpfyhaiJiJnyjMWAXhpaGlMESdBsPzI
Ec3PhBckI5myTi1FSEjkDk64p+Z7zf1hjXEQvQ1ZCHD02Vut/OTuIhQl/yfXCfn3
WbrufNUBt2Mt2JKQVIt+s10nZmoMx58j8ofxtrTGJBdOEz5LhssgQvt59cxeu8Sr
K7/z8jizf0M0VyW92GRb5H3cCjrA9RFwuq/sOkR0undLNVvOrwJikx9PrHJ3+Oa7
hRd2bANaUtrJtRxOFKvrjYRN9DA6Fn5486l+yWBSrdtCV6mH/wndv2ln7bq+ooY/
0Eusdg9h1+UNQPbh2W/KuX5LiX9YJE6dNWNKTFp2pu6Jr298ObxnmYFSepv5igD2
TGf74ARqhCNICQu/ZP9+5MlnFbGpCCc6WueLPno3bXIKOeqSS6HyjUZA+rNT1eJL
eyAXCkwNRoCR7OT59xcfX/ZlwFM9nfKU8lb3YRPRTEdXg12XmaLVBLCYo/rQwPwc
MP/UOronpUeeJz1+mCY6kyfkPV7Ve6+Pn+E3eirWYT3kWejH/8SWwOlr/H12G3Yi
Bwhq3cS7zgBdMEeVmeOHVZWpxP2vWiktx7i4rW9hYngzYyJzaehoucCDTNVkUJgw
0HK8dmEqT04RqC48qlCk3k+BRraFoY+gcxd1YSouIRn/7PY/GtaSVMHAUuyXIXou
zRP+Q8zyHp1D5UNGW2hFbDiM2V691bZxY7aC32PlhsffaV6wiP49gTtSTmfFfzAl
fAX5JWd6SreDFJePZP/IcU6D12gT5B4lJnkDJ/ZEJ6uDXy+W7SnUAO19erQRpX0N
PDKouXuBvFQJ0w/2rAiCDLyPOTfWEyJofDnzbdkKCZ64OMP7UvtH3WnOeF0OZ1L0
/v+NMlV+bB3KJW8KmftRN+wWz0fNPIHjY02WXyD/bHXenxJd6wKmL9J/J/zd0lYL
xH1CBY+qPgSy8fa12OsbNBA5G9DEyJHjSQ32XbSHSE82sQ8JNZomAYVbl2J869+T
/smD2lfMFBfQro6ZqylRaCZ/2FsMOnCvUVMAFXS5yO/VZu1CloBEzTXn6LH6Avda
WwEoSjmuFR+8Uuw9JiGeFcmkCKW+O5Tc/VnXy/qhTWN6MlXWTxNmOT2PDQGA4/6w
2ziV8K9U5VYyP3bUD65o0snJGwxjcbnfPaYXtRzAIz4TaO0oNTh8+CeMDKWcdshk
I6V+GFpmvpvgfVXen4Jv62xNKwQuPTriKBLnNKLq2FFCpC5VZkLdo0J7CHeaEHgg
4G3T5tXWPxdzbDuC4+olOJFFeUEz7ktrjfGzuWJqTWR3JJxClrQO6xlPo34CF+DX
escHEtA6BkmWjvvmnD3haQk1bIj/u95ekuRbyOp7qXsrDdckMxUSfvXQ2Qtwc2xH
9jYX3mLGCI3l+BHiZ5eFoypORAFCvPDlAq95YtjdpzQW0xXRITDJaPr+QZsQRLg9
/1+KgL+Fe12IwfWO0VDrIYSYFC0jU1MpWxeYhYV6J4eM5+4k6GyWpsi2Ogxz3gVT
G9jU1y4zQtE215mPxk1SqMaoxvwF4Ltbkt7EWeIukhHCUSYKN2GSwu/p2cc2SPc0
HjHR/TmPmj8YiXgL2wcAYHNQnsiUfHUkGbs86faxOdEzSGrubWl15WwSMRiHQxlP
pOlTCrbaCpVozX2UaE0dxg+Lqljvjjgavc/FpeVYzbU2GM7+MdCo5+uODTKqq3x3
EO5A6yy/3vBkSdgTWEFCP7hcoN/DP2pcYi1Zlank7PB4n+0prQ20lQPDuMjX27eB
Jm9ajpX/ohfVHXcpHVuBnKmuF06QfFjmKpR1T/usei/XbRMSkCwiRrW27Ud0isMa
Fz7GiFSQQu8eoIYITSRrLZjc8NOWL1M3lI6f1tXBdLaAZ8OYf1jzxeR1vawNrFm2
OOEKn+ra+vP8oGAevM6DnTQmfRY5pppBMgjyD+/exQZ4ZC5RY8Ftje13sJrCiEwH
iQ2CHDWTmJZm1JIJuz9SjuA99vpFGt+kMfiY4kZUg3iNagjkn0/DuPSYbh+1qMBp
FOi/rQwb8PhfEIKgCY3DwxwHHRaSHdce49ihZO6WzqKzHcr8XMMgfvVbp/60fjfK
1r0zkC9FZ+K5srvHPmyE/M0QUNkZhiCCqZTWn3iztKjscuUsHz0tsLtCMFbuJ1r6
szjyaeIqDE+syRsAeL3xoSCLyALR+haqa8TGOgrgVawiCA5FbTiPaBe2WiPLpAQW
Kr/a82td0/ZKRkqN/CO+wSDg9vCC5cSp/Xzcbuq2M+jv4Q5u+oJj9vfnvCjdSx0S
eZF4aC0zGFE90tgVw3dzoG8xuDoHdJzScJunLYTqKXjYACq9gPDuPZG6YWoypmoE
mRU0HLz+MHXFjzsdBLY1vjOLQ8ifsmvNlYAvk6Pkys7XpDZz0usFSt2+HREInNZG
L7CQcT2QjtYfnUGbcqy/zRr1lZlXhAgaIN03qvbzmuU3rcYyVQ3HzNnDxzYUn/S1
z98odAkYoXrBji68s8aDfrz+LvWZTNcyESpnE/IHp2SujfiTNvSdxEWztdjutlao
b8cFRA/fTduVeXuPLon+/zUUePWd4isj+hb9j6ID3hpZtunYYi93ntVp8CMB78M2
9bA0KXckS5o+ydUSaVXB50SuBbeRwwI1CdqCT9CfbQjsAtQtsJIwWsT9fPp0sGKX
gcba8vGKM2S0uu0eWKIc/uiptMXRb2HMYbnoIAGbBcFeD/wSwpKSSzeEHIfyJF2G
to/DYUinGv/9EvmEL12M1pSayn5gd9jHj44yY+LkFMlLbe79UuJ38jQSW4IHOJia
I94EQxvTWDBvo9DgH4MFO/XKPiM12iJSXcK5TKugOSOZKlnRFWFPSu7ecSSQHrkE
8DxKgXXJXEvT1J+mQKQEYaixx+kmLAw9tQbOCyVf++OK5tonamibsBqgFUI4fDDA
TpLJzfYfwllLVFANYY1EFRfvnqU6jorFdZB0WVA03cNSHzyYAcX/sM0c3JIs6aUg
jUDa4hN19xxeUbnmUw3x6eUORKABC2rkgDGNTodh0wo/3OIbUaQ6p1YXM0D98g6i
AOTkxaN20yNJUVl4aSfHSMfZGfuBBQRf/raC9yCIlTmqki3uQif6MT7pQ8uT7OAy
CvQz3vlwQrWsyYRi+7Zyej7l5jxSp2MSJb6vtB1QrZKdw85Uez/gdggCALjIGIq7
V+eHaeTO/g/p6qU7OVfXza1DCOyS9ip5jvHq6D34s13U0QgULW0MCQJW/WgL01eR
gE4w5wEwTtg9ruJ+wFXVVJ7j3za6Af+ayjSB1fLjueG4ldyB/YY1yc9GiJ/GjYtl
OJJCeCqJHij/uBbPdQUlUWk+wznrQa2+z4CeviQ1ExSbM7ZlqrU9V1phQm8Ml6Yl
pyybm9coP1mBgKLwVzQ9BN82Icy6S7DAmv/XT+3FSHYM1bRsQnqbGrK4vTaohX/6
lk8rbzIDRFUttmTcuhwgjXt7Na1fHZDpMviJLt4tbYl32N53unHbKLVF90/55fcL
0p6zyVgkmAblIM/ce1oKobBwH+2JowuIxS6GAsGM+qL0HjO8lBFTWohnGELs2jqi
Ejfg6/7yJz0sCgnSU58WyIsetu+AD4zc+89TC4GBlkkm4jct77Pbh2SasV7udanU
7KP5jQXCcc8yLNagZ/edGjdce7mpC+ATW9yI0/bo338jwsVgif7mqslGjpiBL1Xj
IVk/73OWkMReVivjcjb204+q4X3NGKXVUzaq9XZkrzgUuOxK1RsDa2iubTdrcN5D
z/JCfP4N383jtJeWY49nZ1lV7dNPp7jHRirm8LFAXYbUQexwLB12oX8w3PRm2uXD
yLU9pEGEvgwcQzJWGvLxycag+DH5ERf8DcoI45Y7IVwbFV9xAr/DZUL1NwD8t0Eu
G+hJbFzCW3VHKdzNwIBlT8tqDd3tKtY60WXqyDyMEpMXpxmIZBKUvHT9HKwA6f8h
Wpztt682Oq+Qb2eq7kVvGL5kJRE2fNdVhJLGJXR94s/497AbjZktAQCMU6XXKaJL
62VOQx/9sLPd8NyFn0SIpkXCKzb5ulg/cBjretZ/57kRkA8W8pzTb9xsrS4c1/xk
6AWcuhuUkZWh0C1+Vp6kc8qZuOaaMK/fR1UUo/jBz0PaNcqrBhkrxeMUMRq1PBZ7
kG/BS45B6lcBJI3mW30N8z6cK1oMwZaG3EmF8w+3TcDJhnIhfx8QB5hfqeiw301x
CguEj46UGLHH8hlt+DKwZfuJ3aC0OMIaW9MJGLbyjfNLlBWtf6vNpthsBnWwcMET
/wGizs7t8Iz05UfxSz5+SLdTTkoQFbl1o+GEKj6J3bS9fxOPuDlfPn7SZOgeXRqJ
CoTHM/PYm5UF3lnsAayUPIj+plTJMdf9sDBQK8hyCu9JaxUEkrajjtybVRhTJKQQ
3R2HObBdLqEZE7yI7+TJNNCaU1LEdCWHpzm/hXr8z4g2qoh6KgsyYHF5hX63hPD3
/MjQIbLhHHlrkleWMcnN66yBuIDjltd6nqDLPSEya4kbfhe/f8sJJ4QDO5R0xh6l
ggL8IwcGEgCFDKN5ZppA5G1KY6qi3NNecYNk2vU06cnIYB24WdFedq5WoePVshbD
LOGIMhfvL1tRUySxMNEPNlYtGfKmnAsXcRqnZZlCPlrrqoTiyIYJ2GugXPKm9bOr
4k51BWeGnhi4wS9lAlKXl5Qt+GO+EtulPsMpa7kwacRDrsfJ8bZG/LKj7H1ovsWP
6+x3UkbpL1flssDOl4BOSO8xKWtmqi76Svb1pQarm0pOLqHPtzJOfnt65XtCRbqM
EGfqDu74T5NFuuAFVOj4YESiVtIuGP47KP5/b//WPI35v2GrC1T9bhOkJ3PRAzac
YeL2CSNLgo9chZnZTZ4Y6vehyeYCW/s5GNnKjo8PU+2SIxG9KkMp3Y1NcP6X+bwA
QkfXgh3TEcm5j+x9jMFuiPHkT1cviJE2ZisI1Vi7bprcKcLcieA2qRBfw0dGWMmT
KzxOVzviIEfm/RmyH8a4VoZ23VCeiGtMNB0XnYjwWgIFHqL30zSEDd2s/k1HZmoD
kjMy1Fo2vAwl1f1M2+LXM2XLho/2Xpg30LMmlCvyPNWaWZYnqcAH05Y23rDQz2BR
1NSAT24gF3M18GsVTL+w4OaJlbtrBbmj5M8rE8xHwYmb159EHyQb0zY8kpFsDANR
YLO6aq0b2nG5HxLDI8IQuUTHrhVe+UAAXq0YfP9oWSgESOgD1Jb2Jh6fs3563R3+
mo0g13ryFf/xRvx5H+jawgzKgpHpLb9nsCIz29NhW8riGktS3lOjW7poBzSjnS1G
XbhSsDNv/qA9v2iBXRVQMPrIfpo6rMeY61Qm8bbjbtf2ItgWFUZxZKUrAK/Nnj5+
rtCWPvcw8/b8AjG88qJfGMRJen/Nn4Z0+lgg0CFJsOz93sT0HBFYa6uzvsCqbpn4
yfD8ogHshVr0fNCPTGF4sJZMfC3yfY8DO2z5H1f5rFXs6VoJ4zD60KIjoHCzN4jS
bk5TYgoewdaxncxF0Eoh78skQREQabTkhnxdIWzLf+231B7MmidygQ+q7khZaqV1
afbdUgcTfH1HwFebPK0PfSIKrPLtmfxygYLFrYGGW+8/N2tsDmFAPy/md1lW1wUo
8QUCbZQAwMXZpBfHG8N8kzOXQL4M8rFDSwhcdK3A59ShyVz1xZUEvbPggqzaM9AE
rMw3VRrxM6vv/BjWtutGYYJMJCobkBOWDiBeQPhQGTlLGO4laCk0GehnQTxQLV1L
Pz1B8wYph5foGAsm3BbznlqsVWu1raIFWKla2JKG1OYgM0Xo6xZjqX7u6z0CRo+p
K8Z+i5isAD8fflNjEZkLIqMYkd1LNiWbga9jsuwU6sV60BGnh6LJYAXFA/avI2Xn
jyEDk9JWLZaqFZQVwalYS6XTwUN1Z+ugKfmHsfVeanFa0EwGyZyole0NdUb48bMW
6wvvNPG/B7EyoXgCOYWRpFGgom1edXMptkQSL8F9vNhU86YM46YFGBfm0aogqu9U
MB++34xMriogtHRcv5WLGLq1vt/gFA07J7/yC/Gb+Tzmofdpazm2Vynw6mFt0hvQ
jNYcDLo7nz1q9S7wcGobkzLzSe3ht96eu3tr/wO2KbdS55ZWI1xUi+MC6F27Tnxq
WjZNfrw9EHKvPGeebJhMOD97lla5+z38q9OSAqaluoSZdm8PNYyCcmcF9pvU2cT9
5l2xQD1sEjPDbr9rjvkbZkTInhEwXt0rrLwM4vQHX/v+5zru5CXOkICPApUHGaix
c7H/Q2OaduUIi0mcq2rfsnlWwcxnMu244qtrQfOVUoZBmieJM2fE1BcMxaRe2fO8
DcBGcRzTFD8MMDZ3l5BxQhl8Zqi5bMjGS4hG/gB8tQ48KUqFXNyH+GqplfS6H0NA
ax1dHZLrAvIGGmttuQI/W6kmYQ+SjGS7jZKHhXBk3EDBGZbYdx+nHmUK9mRU0ozl
OVyNR5sA8Rs6ngLoWFeOTPH0xIalchRDXK117DYVVeRWjimlSoUUDd1IP4QkiO0f
GOlYx+vUJrqYwZKlgyZkzhVrRq72LcW3cx6OqCF+bElshAQJRnhIANQ0f4tU+us4
xd3XyQFUEn1+SWO09td1BZ3wU4NsBC+lXNQY1jgzR4GXd6V7uotNOPRy+gOhD7T6
31uI3ipS6U6FiiCNQBEsBw3myFLQ7zhnojljYdpaNpLXzPZl6530+X/aw7h/Yflg
5fSSv8HW9ez6MxfqKeq03lR4OCsGPm0fo87HG/Q3rMOfTd7SYyjmL+OOyGVeeSGo
l5Cr3LJKzL6tYaYpTBosngbFUe902T8WRpUt3pizJgT4FvU1XGqgK+Qq2X02727s
4vxLGRrxzrrVkgmq6PSOMa4m0ahSrz/4bEArEJLyegNxOOJNy1tnoM4vU4ZyzPcY
iSfISPeEivIbujubQ04Yb5SyP1QB/0Fc8iDxalqlc62exiiVbcDyHDkgfb6fN9V/
iUbbnuH7G4je+tqFB1K+lJjYTpjva7mzNHe4+bI5i6z2WVGjm7wRMf6y0cdVIRbT
QNXvbkN2oPfyBn80P/hCwlugNEp+nRhFiG3SzAWDnSOF11c7C10r9qpLPolZi/IZ
Hjjmfhh4TLKP5yOGEcVyuNGtiMRpPkecu0A0vUDWwGDh2ky8/0AMK2ay4q7X5bTf
v17WWCHi8KYwJq10pRNXfl/BrFuMoPFt6X2edGZyz5r2KRi7Z7IWIp500MDoaKCq
G/gDSwBreP+o+NLygJMSjJJcM0RybAqxrWAHZq20UOfYX9vRNbf39kdepwrPsJOv
U8+bxPr8nqlOnPtDlX7U68rGnigKWnhWjM83opzcco7gyJse0OUOJSUHDQOpo1/r
zOc6EGfKcuTmaOax30Tg5LeJDsG4aKkN+rd9crh+7l9Taxt8ZNa8y3gqpO9v4SOn
LHtFjDdNAZO/L6Nu4QUC6JbcnC46NZ/bkmMI8PbH6uuNXAyA8YBjsWRKXqWop+PH
EX2UFiWTKnGPiepBE23/RnEofbCatnpmWAvyIx3hkCn1KR2w0cTwjWfOTlVoVHdA
Sgd61YpFOk4bpR6xwQNayYgpqU4ANtjrjAEBj/eUPH4VjdkIWX0RdO8djfONxdI3
1BVFf3ylNfJRLdNwblbpV388dK8wGD4j0bcJfv/vkbHOc8ISiciRMDFKWnKsttbp
DtH0QoTSTEP8MBQyL7Vsx7C6W8cPLe485DnHCIX2Fiu8wWc/TftvCLAvjXziADqI
5NPaor+XeUk+menyVhoQjknRvfyIozH4+ZcSNLI5e/bf8l7+4VioNj7PmQzYl6/5
DjT8rixNgoxehXGYClB9bEHxHNc5DjB/6C+YoOyZgmISgwfdDf3PvD3D8HzUwyBF
pMm6tSUGnPNnKKB/5oBG5eMH6n5x/DYvcmaB/alGvdv9B/0YV43oofTDx4xfHV+k
6ED3p79scFLP3Jrkb01D7rDS9Wqw4y7vLS+aqTTr1a42tUowRHs2WBuYCE/dl0iM
/njIsUsnenZp5hhH77xInJsdjbJuc2D3NP+c6NhZDW1STJy2JKbvYnWZrCxqykmt
5plaJERSbqaKkDiYmpOGamJo4hfVI/UHjo2lXnokB8Irr2j5HUx2+l7tVbtSBwem
5KCMCUoJYS5wC76bfuD9x+HKlxhjhAWDnchIRiVEanhCuFk/gpP99d6uqsiH0RdA
dp3pMMlaF6yvGoZY6MQssuZOyzkVaGqLrqejuMKWBUGk75iXmI4IuNmjSL2z5Irg
fKhEpMRiZj79IefIEnj/HcnI5GMY+deemKQe5PLNe3tIUQm+B+8527J3YrcM+5dE
Dq/POablUerQ8xTR4k1/nXazwDOjzLlkN39A5TIwgZ4MBvxnlxtf6/czc9sQVbdS
TqkCMDXp9obhGo8zSMQZ/YB/7Aj16yyg9cKi9bqk1LD0g76QrHHZjwYWu7RNjEDl
ZDAV5YUduIA4k9cBqxhNAI4u2GxdzNz8xmC3ELZu/rpiy3xa57CNP/zewrTCfTY5
gPRzkYyEp+T9YW3wOBhPxSzgodzJ963tCWugDFAckC9yAh5XNW6LHTgqAlyaB3kP
+xZ1vXvFQwzgjWVqBSUG+3ZZ4L0Y75DCt0Qrh01QT/sCFha9NXPZpJlc+oV1+Xsr
8DnsRvBH3Ygw3Nca5f6yn7U/EbcnC+XKd2qOfscocftCM5xMGxud0/aRJdB/tJoT
/xUStJSQvESyf5M9n9XV1oYsioMWbfNWKM06kTzMjDuDZXpwNii1DtvpJbYKiFIq
zGk6KmCvFpvozJhvVumdRHjJKbmyBiYUYWHUV9ZoQ22YrvivU+wY6NdGl6Cf+SCW
QHdZzrtsd45I0krnxhXytwg9eHH/Dc3KorVAEnTqMWj/LtD+VLwecBg6Qirz6/S8
LR8NrwOStwAM0EUoAoWrVan8zSFzb6PpOuLUv97W6imQLIvFljBaW2MAJytQAhNf
buixZL+UzDzShK4QYvir6K0X6ZidRQ5CSNQwqUVjgfk9L7LUWRny9c1gvRl/eIoe
l4K/MOloDz9hjx13JOTYQoAA3vrBY0ASZ5/XK37vn0TpdqJFQ0/cqgZEfL50dTvq
+bZncDR/w59kCqg4vfj20nVfFKI+EQ2IORt3AOrCCrx1SOnIkEMyv/5Tp5hJP/gY
mAmjkeZsLC5dETlxMe4/xU8f5sKjUd09e6z2JtVUar8xukjWFBjhQfeJn3XSoe0c
SgAgyKew7P0An0x+5DF8os0MYa+ajZPsI+UCa6EVz82JpG8uYTtfXLzEfHz7E3Ms
+eYSwJNTRgx4zCPXM0VwS/6weuoGoowUwg4gVlejxEnmqiwJ2r0Hqc/IW+a/Rbi5
AlKSD+/YuYjbI2ztPEI0GiAa+rr3YT0AkOCh9MjFTwathYqeIi3939WfTuYaDhAR
UZB3/mf3cc8hhJmEXfnB1EKrnjn4DuYK2oMfU64aMLlinoQHIHmYfr4Q4XCMM0+i
CUNfYOLFGhosjmvjRD8raYA4ouMEHkYMcwGq0+0WiAOamkJsh1immpwTCESgFxyP
hEJQsP1x/K51ebiSBd0ilrJVRTbpdY+nhSNDcf9MXf39HEnEmG93WzhlMGZCOAE4
MmnsFs49LHO0IjrwUNpjMiYEh62PycPjQlTG1Nypyxl2sMweb56+UJjM1ic5rHs6
bsa7udJOrnHtAQszOfIk2ZWYojLz6g6UAopPWnzRhPCp34Y3P4lI8ckr6cHGsJlx
MOM6VvufrOOLVCfRXZyWmr6LMQGEofwCWIvwGAQkBBPTLvc+pA/dvCCzGqc+joyd
NgJfO6M0PjiczNodoM7oBbsVgE7W04J2PbIFHdtsFa3nSpwBqhz+/KoYHZ/6rKlH
ziqKu0NPXmHtGgHKOego+VCPClgrOFSjBLcRbaMeivi18HG/lPn2tsvgLEZ9UQET
CUPFlQckD2/pjG0QEpzBMHH2h9jN3HvZCqU4cAKWPQhPdGHLdQqx9e29RwRU82rY
seJG/TuIJWYkbYR3LKo2C224iCGxPrYu+7NfOXIC5oKmWaZm8Ev94ClP76CfOZej
F4yiMXF2lnJ+e7U8Q2rfxhbMZSF2AXwY7DxYoMVX2AKxKoYfYSu5hlQCJSwUfuHo
9xk4yd9IYBs43u+db6CsEB40Vao5FsVkPKgSTwDI2egHjEwUWaop/cbb1yb33u+g
ElCWoayxPyWKvCpu0hZJOzmK+bmRSyU6s/P1uzS/wWS7BbLn8dqZfX+OkpC5grER
09ulSS+F6XD+RwZM+Du/h8jNcFmtiVZe0r+PU1kiJWg/gIGw32mqH/5PpChSkSNE
2oQO/mjwCst63J/GvPDqPb7VQ+6iYD6OKececylElC8zT9Oln457in7Jls9PMAL3
An/oLFzYvTPKEd6gcv7dURzVMOsOHomMV5ftX8DBbUpLL/UlAGZf9OuM6tz71VOw
DwNtRap/cR3I5NGXagpqE0nd4t7AkPViXXV3jwYrqzqCVgSOchyJvmQ87rFucgt5
pRbf/f3Sv3/urHSb69vvORnI9nDfoHF6+Uc9wzPtatvBBUDhatGlReZsu7Zbn9yQ
E1alJQyBKLV+eXtkfWPyvTNJCaoIL25LZJBP+Qf/MxLST4yIrzVHlHA0LTlU1/tr
Q0AC5LjMjqUZmk6Zb93iAIMavUvY7q4IZKkCa9Jk14xMnt/hBZjOFgv460uq3hoX
dniU8UWbuajRkmVapNMjpGAKlbTJoyd47FedoaPIj6qO4rOxdzKskL+R0bn0TcLP
nU/PGiNQgsA/87YGPu7Z34EsaxhvXsqFWF6Q0s0UoqCxUiSkB1yH2psIM4aylSag
fSeqBKvjNJcQ828GDfvei+SR6Gof09GLEh/O9+iREwn+xjY2FyzGDMTJGUCuTKns
BSLpCW0MA/6XyuTGoXy4eEs4FahaBXGbVjag3DzSWUU9T7onvKV27IW9h5ep9Ulc
nQ1DR/OOAeCaCAnh1OvxNucXuDpSSyiTj7lARowIdvE+XbBHhbpcr0/5lbg42dJl
n3dnLW7igl5MrhOMyoMG3t5yp8Lqwjbd7WQ6vM6QVOzA8IWFQGjtsSjBKz7Ks7bq
UefBuUlnScXSUQ3sITdegD9WEQn20DWGIs/CbcCrT6eFG5EKKfOZ2fQqnIOlINeD
G2DK3uhyaEaQes37R4QGJhjk/0aRfOSFBTcwuqGRn8M9D1dQnZLHghf5J9ZQ1Mb9
3vYNUwRzdiCMclO+oV33OLtsdt4htDVGXbpgf90DiyalHiA01JvHjQ4U5kllxLfA
4IH5rgYTWiN2GDF2vnx0nVE3ALjEDkQ+Nkdm3O21t99HUTM9xHFrMTiEro/y51d5
woVh37Aq1/JRa/QGLgOW9a6ByUPUd4Pkt+rM5WavABqQN+b9LFKvVKZq8+zn4faF
426maKYsu/hb156qXDMbuhO1EbN5lC07uaf2ueCAOTGV9mZLhNUBUS3ep6U/QasK
8ItKz2mjNAxc8g+Zlzxg8DXh08Wcz0abWTrwXd+jl2Vp45oCkqZqyNOghAIxZ3DF
CLqTED1oerSA0b41uwE0dz0q489xdEBkdji+6rcd33hztsEDOknWVzpB5fw3uMUl
FnqSX7VzuTLMw2rK2i6CKOcDLUfePtMtNWDsX0nbiwgi5Czec08fqGXodq3wAI2b
nl4HOore2FF4KM5eL2rAXMRy1MxcCAQHchoPnUqrOuJxzxuYTQ1mOS1ogMmmqZM9
uqCBFBMzRyUC+KY92XtAxlHGAYWhZlhy8sjYjA/LfID7c2NjdTSX9RzNq013ZfNF
f3QRDT0x/SFdeEuajQ9KoGNmXAV7U5xO39tDNEtHUtEZH5KEUuvKxv8a/s8Xgxbz
gLa72ZueJXNifdVGQWTALSmgTS1jSLS3mzwTZT9rXzMkOMvCnr+VCMJQMGK7KyKn
u0hlPafPMDo24fWRuPfBlZOoFNUia1U2XzILVdKGgi5CjX5+VrzLmSdCHkAUMY5F
N9uvxIKm4LX878udQa7jxfiJgCoYV4aj/lXrUvJPK7mT3h09fUmd5TG+tKS8INRk
JiprPDFVlm7nQ06emfw+YbzowTad21Lsu1dlYspxC+kVCvI2EPNlg/wkyeNOza7B
j36Ii0dJmGOc/D93H5vYFAtMJqtevlVy9FPVTl5icmBdTCDtRLSMnfCKD5fcLyQn
GgbnnAd2OB5abljxHo/K5ENoIg6GWxiWjCNUkKWQz6yoCve1B5UdahKc504U3x0K
MCKvGO1zCgMMyLfnv1QGP8e+My0NAqHQm8MNb11e5SClf+qp1eFUhrZawdw+zhWE
k9IjkSZIPEADz+V5DHfxM+z1ANnafyBvnguz1LUM93KkziO0bpvnSuRMP1Q+tjKF
ywHutKAC4Q4uRftE996qzKi+6yxzIMBG3Zeu+5CXDIkPAfqEov3Ozlk2j/D3HYDm
fK6DFTrAt8F/WQoTZ8P7mVIJ9JwAejUSscH0UHz5XY2DEKPH8m3cMMTliTnGLF4S
ACUsTOVb6WTaQuR2FseVzrsF64rjEFwt7xkI/r5e6YnbYhC3ibuKEx/B2q78Vo0W
rRsfcr5JnmZHMGkSx+RAidkEfJ+VpvaCblfpeZ58lQRz8hKyCHyozW2eMQsoHWYJ
yraL/c6SRos8g0l5kXxDTQgxFhQwEtYVO+TndiVvP112xvKyr1hcPvMPIS6+vvAi
cn1t/m0+eqioIc9eC782+lN7dzl09fJi4m2txz/9nO9fe+Egy4GAz54ItQxJhSr8
1+MPmw8GLLaGmTTrKF8mrDmNKU1AN5/aqscAQrYweisblaxroxGE3dPYOWhuYPyQ
ICIPsFzcsLa9yqwPcRxz+vIsuUjTS/mwSPurpHiaKithiupBqBv/HHynPbepiNfo
M4T4LJGEV68EblqIlyQJao8R1ULnnf5cWPJRBSbzOeHMk5aLi7aMXmvc69u+jjZ3
mWa0YS1Wvck8TyMW86yPnoB3r8WBTKkOQmRuMXykO5RiSHeK77/L3CgNRED9uYX1
sIS+RaiBOibrRhd8Jis4bMsmQQo1wNEjaZVMvezCPRgdyagSZN380AWABouRIfWH
kgJg6TeO57H9YfZWab7lvb5IEs7Dgf3Opbo0vEUOlbtGY6o+AP4HLFLlpszUfLvp
xUdJNAUVtsB0PR6lsYRyFcXRKTPGj8C1OKT/EwZAedhUAUsSZwQHOrcQkGx1Q50s
fpytLKE3a8U3bKQAije0SxTOZuzC2bkLDmSLbAkgHKnd6oF5PG4a8Dp2c3qBZ14f
Z/sZTu0KGe5T+xWesv3oNfq/o9nUrB8JheXbWlzyvvcgahBj7GrdHlQArVliKY6Y
9/RpV/3znOl91B6QTfxXMMuOGCy8F16jAwOuU+lIECwP1IpIuwSRqZvNFzOQU26K
UFQN6e542oeGmtNpEkzFFhhCBFaAjyCCqjJKedmms1sdoP3QY71p85T/hG/OPkVr
Tp5QotAMPaqfQXP+1hXrw2JbgqYU5zq8/C09Peh8j5/OPq8ZvsQ92mRHbLNhzFoW
1grqw7qUTFEIAM4j6ch7fgADVYTc9hGUi/dZlOjC0Dq5Y7Q6KeQAgxIdhOaSuJbj
Q8YaocqTyc7AejmJg4UEasbXz/9sXWLBL/vEgKQqgR1lv95IjH7wGKKq27F+vLER
3mzZ8liiBeIDe0zzTYgH2buzsRh1ykTgQN86UKgteyVV14nfKCgm4ajdRaxi74at
p0Yi0FSvNKklgBSl7DuW7XFtLHGBeu7pHXgaaTehW7GtOkl6wGcoREtLehvJBUXa
vmEVTLOVzvNth+k9FmqQ0hwDCBdSXBC5P6Xcm/NeayW17VMfuOqVogB6uXLoYH80
DIh1jRKQPyItwTnvybFTzHE1szZPePVgsdNYF/HsM671vwGcr2/C+5/wARGRgCrE
I03ffR6C+CL1A6Rl7Nyir81LZUR/uFj8k10YHi7ENc4s1AHo5C8W554m6m3o26zx
nasTPdR+9HwBZ/Bt9fBwDsmUcaoYlP8I34ayeLlDRKRLb8graKG0ocTbOTJUly1k
yb9zioYRC5CHhCFC3X+XlVUyycEEkonMx3dgW19Xbpju68i2lfjWVNgNLMwNfxkb
DPbhHla+Edu4jKchlasvvfig3bz7CnCVPPGsLEqDJ0rZhcrwZj/3IcT8PVnXwWX+
jGpCJZ49aR3kCVnM5Uvn/R3ieRFrOvJsjlHZMM8DFRo+ECefO9O+pcOHHYA47zRG
72ZbIdeF4Z36kY0Sa93mhHoMT6qsz990Pw6Gs09ja1m6e61Jtq7Hy7CB9xFOuwg+
gxLUR+opdVFIzl5wbCk2HnGaTS8jSvWARnMDhOyGLgGY90PmJWv7+hljCgxzexoC
SPo/ggAyvmv0uwAvGJ+EzjENsH0uHIXlxNsaS+Ad3N+OOFz1mQlV2yGsb4GqKPxP
j/yK93zhSHnctHr+35aI0yOSgg+cmvjji/POZmdxiEtkFveJXe8kCzKs52HF3vq5
VbYSREJ1DnXjBZi6UieuifpuA4idZT1tVqjQI6zdR+G8XngKpwehWHKtfIjjPh43
LRdwOjvq/W/NRynsrkL3g9DHSuEGQHlp2mP/OZ1hx9vExo30hcaxppC1w3KP6yv2
rMyOod+ofGourdmV9U8qAbBec8nmOUCpsi1cKJHd+oxqD+E55DazyS1HULOmRAK6
CXKapSKDBqZIhehovmq8gN2dR0btG9gdbtQbLlFIbGKEBkk3jQUxw/wgrZSp+MV+
mlkQGvxpeN1X/8bs8+g8sjfQ/196tdtr27qjxktzcIBH/wfrMyJ3u1LjTm9N7UzE
Oh0QG4oqtUT7e6TbJK/g3d+6Mbc9Ru7a0EcM5pGrxgnnmm/9gbnDgSqVm5zszdeF
3uh607VSofs2QdiEkq11Ip3PEQQNxeik6C4/tAGSwb2sd/TTcieWvwJ1C64nk/rA
4jFralGJOTr9+n6IaX6J+cjL0gLc9f4DIWtwgoxPwCsS336yAG/tYBRQaj9FxP7+
cpEVDbmudD/GBLfoCDGccU14+CY/XG7Zc3+0F1ErIFCPwNjjmv4yPxpd4AFJ4tgE
QRQjcw7PMnOPqziVdqA41d0N7cCTfXgIMXAU5Y/Ss1ac/CRqEuJxCR9cTRLF0MHr
yCnsR2ClN8y6+IS0XPky3tsE9DE/g4y3S3EL/CGZNHTjUbLF8khQvIEZVnrGS9ZI
Ie5/YGS7xX5UYjjpMKrq020O7vDfSZiUkz7++jZ2Sgd5pSodeMNF+ZTIyhb3Djoi
JckCiQZxqd8VSd0wU+QO9R9QG6AHXXtxSEGM+YgYlE08SiKZwuuseUQyrMJwH/F9
5nWrOlim4ZFlbmE0g+oKmTzKGNjO768Bvjy5Y2HhqgHUCXUdTvPtSOCm+Vgo+SB9
6Mgstx1l3TvnekD7n2rKOans7yjl0+b5JPRvFdnvbB7c6Eo+h+YOX5i/12ZsWs0d
7zvdHVSZRZfmGpg0uAoVscQeDNVlIWSun5iiG9ijfJvl7xNCLAs9mtmJag/koeDm
E3gNzTtxuxWLv6/h5RxCXaPFUHMNeT91cUC6RFhzruSHh7JbN5ZSP1cv3BuEBBBS
dAZRGhuVp3GGsC6y1xppzF6KMN+Ro2fouUQ73Zz3AiSMOJQBGq9h97+1n0kOdo2L
Jq5AK/mASsNHbG2wbD7xXcDspJ1canvo5pA+IjZC6xlWgrWcwHPKsxdCAk+F5sz6
ZsTCGlrSbElPcq6U8uEf2qewRJ15qK/PU9B8uVp0M6aW81mi7p7DoxljEDSOk7C3
0HWCRBSzHJ1mQxM8ZPJJ2GZZXScMT/20K/YXW2TfVAsHYHSNAtN0U475+2BKrdAR
jZdHnyKEalJnar9v3fFaLSoTmuUVOtsB0eAMBmossifwSQK0EqvsKp6MRP0siPCR
BibzDWThpHMYT7wZwqlunHoUBfd6dytZD50ZkzugqPf4zI1RsfADoIREcm/3Ivw1
miVuuD64Vt0Yfk4w1ryVfPfXIKv97L/BAHzADroam1zsNwY6IWSfpjBQw2iHZaur
C9ApHapjOuYll/gsmS7ZgGCtM2cw2WF7YTb5/a7RlWg7S5fAPqNxfckjntrWSK4K
8Ioti/MXlJWZAIvx+22uW7k23a6MoPNcWq0QEnBYf264vEvPWzR1WeTRCrrxOsrM
/bN3Rx9y3KEqvJfrRqKaklIQpwwH8ahgnMHT2ApkbRyGDXVn+rSVzYnCQvLUeNqM
bF55BPwxpoKpR8NpctEpxTgSYZXzmOLfaj7jL5gWoQJo0tXT0JDowcE/lzBxZLRx
9fPZKBS9AWzBjNbpyw1rE0+TjW3MxoUxr2yzVwA59C4/1HGlnJYeRGh4ZzaA4BoJ
keuASmwOhgpVv2FNBpRcLrU6VyZaAz1eYqtGHkIlDdXRgo60GaPZPU5xCm8uwpTT
j97jGOCO9qCM3Ge3oM5u6SjINUFHqIjfaScLq/tCuMoWhc5eIcJFr870Z3vS6yoP
u6GEcbXv6x9jKxuWtgjEXrMol0Wwtb4spOTEUoi0T/mLD+P7uJg3Dpx0hhIREvvn
jwaTSMQHJsTMxiuEXIafkf6xfexXNBOJXAM4S824H0jr18BsnpSbg3/Tun783LGs
BcV3+BV8ZeW5/n7Qm7JX2jP8NsUoOqnRhRdjQcnQs9u4qe39c3msMzJ0JBYUvY7/
8GEn0bLJpCysCxGXx0XCm2n1ehq7OBUvoSD/tQg+3VSutAY26JZFXJFUTkFSkBXg
VqCVnhyzNcormknc347Vi9nCCXXkzVQz7DorK+IMebmvVZOgYFo6Yr/1HhOE6lQw
AAwzdoYq4jgAE/jiwE24Ck4m7Pa+m8LtmDUCCxuXYR//RoO1dOa/QMFlakuGZOqH
KiKQILBZbFq0/JoDdfePL6tKMCZmWj+t6841dlwH/XHxYYViktqYNQbE+TZAz2hk
58Vi9LxFg6j3yf3GO6Ecd461c2X0k93VqzNT2+ZYe2LazM2ownCJUwDRbt/ISG44
/fkguY824wl8ojqUaMaleheHv7Sm4gYj77I+hokaDeLc7KM8X+Mu26YyHpBhg7E0
H1pwH1tYODd1L9btkcG3J9M7K0t2r0nY3vwJPsc2pBwDrXqf//QsCp0+dIZgZ4DI
r2bWhG0uczBQ7KZt5j9Bp0zXwUNcOdClffp2FXH5s3DU7jLdTzvShxEqemEPXQJ3
nE9N9UWkLzQouMaZ8w/01Y4yiu2Vg/Kzt4wAJg5vu2kmZpwvrvYGnkwYqhgrBren
h+UGvFifCa1zT498R2saYqlkcKPGJQ0kB4NV34H34eOXlNw6AmM6llXhUHrVO9Mh
Y0oCDV6aUSJQYhCH1R4VfPrnFqoSrvjruQXXp+htxKXsVRI6gX6HRroaxR8NncSj
TIiiJVOzNWoOuAEsYjM752xXvAm9w3W0iXo70bra8v6C/vtOQLQk1N3LRIguVq6/
Q6Of7C0V5OUCn8FS8daQfFRIEQCHh+ndK4+s/Wc9RONPST1hsyXdEZZ6Oj24W1Nt
eaDf33I+H6MgCUcmlhPwY8XzQZAXa5SMupMqAZQe4MHvtbcGGw86DRhpaOm4eezE
OM3nQ5uaBf+ZZEtVIHmxZQ0bHqc3/59fjQ8KsWeavkpC2Y2SVAV6k3qkM2jaBEcM
c6jZs2EE8b/xrULw87A7re8MQhjirHeCH/OKN6aw5PBi63gGPhDjSeLrbZi2Hdkv
mapxVlJEQKvfN3SNJAqUPSeD4XpMEmMkme30qNuLt2s/ogz4AcJm7eBQfvYX/cgW
6YLIAFdlK1UxQNI54aAKz/Gl7nBO0NnIxspi3XrCTl78x6BdTbkTJB1EVGUdF96i
Z1srFyOTGp/2piCvikxFhBNifvSfqT2UmkxynU3eMg1TK483bGySun8Sk81KhuCF
DQisD1F0vclx5nNoluKs7UxoWA9QsaJ5gtRc8ox51bokZS9JUAJGKxVe9H78XHJv
Lf3QUzdGDmDuwRDBfdgxstvBVGWreV81Pyk7+toElYpqtoAYUD0f7AyuepQLc01b
8ZKPgUFWVUC6Yzet2zRySZOtgf92AAG0LXPrpzBZkECjWuhuG8oMm7U4Vi2EqLlU
NV/piqtYgrTij4iSOPHG5XQtqsYqoyUaTNrz3652jAf5IMRrLxIfdrawAECdzm0m
B3k+QrJ6eeGDK2cqNQdwXJdkXatS/WLFWlxEpPlRnUqS+zSvvYh64SZTIMRzEARR
cL3w1vMJc81D+6dXSTxxIWh6IaotlDTw/OpnqvY5xcS02F5g4ap6YAA7rX1H6HbC
cfriLX/5Tdrpf5tcb8kIXnKZp4d4CH6FcrPDUe0NKuAyAcVvOMLoikb+QgFsFdlq
fUU5ptLDTyJLZcFxzHudhu9Wxqx+wyQsKLuLIEvqnj/p9iE5JanKQ392Gvb+OiLU
h0wSxkDB3sTCedDPshWpQzrjVD4Gkzyd8ikZBhB1c5TmVF1ZcqehqBswbfR5Qpgo
rYJ26Ia1J40cdi52bQEKtE+1kHckmHzA+3LW1iT2mwiyhzEFJyGwi4oJ0Zd8Yap/
8UYCjUPb8WgymHA1FKUimQsd68VnPIslMwwbiPDbQ47TQqcLiN53fE2lta8FEJdk
7XkOEO/vXzRHb1RKCSRx8l0YjEmnByOC3/i/0GU1h+2Z7Qvdyn47kK+WFfeLVFg/
h+MVL2kQsZmLhLQT6CYsXuaS/y/PypwigerSmPhwYATKrKwMoPGzjTX4xYVL98mY
zwoo04Um05rv2DNjy288plnDhb06o9z2m++l+0tjBX+pBg8z//FvjOcFNeox3iVO
caG1jrOX6wYRlBiHe/paynHQ9JwdM+SF+7glBQOOtuwJo4jXA6bPfq7SL2SIDvfg
vHEPXR00fOgYeROhY1KsetETo4Ve/IekI4jQvcg3hBHJ+jPSJsre6IbEyIQe1n6b
T0u7qclkdas1JpPN/qofynGbGR/07dWkZ2zI/5qm3WH/OZ/OK08GQmb3/amj4NLL
wVCMHO7p3eQmT2crf/8z1cdwd5yoSsnW72Ox62RdSFQVGD2Q3wKkD2ieGzmNJivo
7UgVsibAQkCkUvIagEbmz9ge8bLQkZJUU6vgctzHo7pbrykC0Ch7Ojc0sF2W0aqB
TGWuIRqAbXQ9BU3ce3KkuQ+ILp7zxr5l1nnR+m1mnLpxsfYH+LI6yqvnJPkmsTuP
w4Rt29qNCc7yEV7rujIcDaMg4snxa8KiVmkBcK4sFszdhSLD0Z5mB7PGLKHsL+I6
SbX8D6tDJGYDcuPCaCrtsZiTWHbvgk54lyYFNGWCPsj9YOETxunqi52kAxImfldx
FFrFpdS7XQV92vow3IoR+N52q5v88veAaxf1kzRxTcXcSV2AO4GWlr9wKB7rSf9W
0iZqaPQVGQIrtq9iQH9PYXeFKGh8WJxwHUJupg3gZASZYnTowCV7JH46g3nYdd21
u5gB7Cj/wXy+OW1hv0Xo641Nh64WGGVZd9lKCyZXgnd/aemFeVPZHUEgKHVPWWLt
BHBoS5H9xK5SKRiV3yBTqzDLdv567JE41RDAdRo+KfaFYu0XAh4z/yhixDoNZVF7
HPWStcmHJDXO6pvPSqs/gT8wnp6YpqXheUTSs44FxVRAkxSEk8iANe4XYXRBhh7b
hcEM6phvgGkT809i2ZFqYpsBTHsRSouyfFFcmd/DHvlsqfRwSlMfwMimJ8SFIaMi
nUE8XuYmf5dpAtQcXvx3MAZvGmDT5fIaEQoE2Z3LcxxUMrp1rNBNLHDSnaFuaFWF
xSkS3l3DVdbCj4VMJJaP0Mj+xvnUBYKk8pOnjeE4pgH3OJx/mxmsBV/ftKJ4+9Yd
oeKvpznH+ggJNW4ZpaPs3qIcsPmvg1z2O8L5M9lqnxyvIjXl9FkGeRq+uRwj9tVj
AG83PYKASxLhkPd/mE+52ABCqFdSf/uqltWF2o5EKWuNvn8vSwSxi1DTx8obPQnh
A71kOZYrH6kslFrreup4SWwQP1HC/paKImeuH0TPmkGvg1/lctUonmRql/5STeJy
AW0jqzJNNW6uidutnU3UXeg1JnSHCWdKtrH6oWQEVFI17Dv2+5N2IE2IHqtKKaQm
MetpUjhdcz+J5a7PSQp/FflVg1oHIPiwXYXXIQ64dSLz+uKz11XuL3sAQu15BBQt
SzCQAFdEfpJR+p0zaJcRHBhAnOzTzCnDqvK7RlbXd9S1pX24R+0qkDHLQupa0tBC
DRMKTSRsoPi1aJsW+j49abKktPNWzWPGGPgIAuxs+HNqSY5h433PfRnJkrAXWzEy
3rhBV6TmwFcwwUvfGKrO662UtCz123OXlaNSynWjH2P9IvfAl3vsNga5AlY5gHDb
qL4DofyGvVrhhxTDZmfKzAmraOR89ILnKFNHgwjwpxiEbskP+Acq6gogXfZCSuM6
a3JHnMWU56nI92Qz5Fc1seEKkXqaDw3eYpRII8Wv9C9I4RjSRGlC8beHRCgKg1Mf
tv3bePqsaVcGcsB3PtexjQpag1JK1JJYtiB+8LDPpkKxKQgf7pxW9KzC2dwlO0y1
lvq2ugWEJTCSYD0SbtXsfetn12RbJMMhz02hjSR9iDWqaujbMfRibgunAYM7BYZZ
Ys1K368jB4Shcm/h4bnKSMaOobnLb+AadpwbBntea1r4rvJhuyVbj51kjDhbqe83
OkIKiNSiAW0OYdIQEV5MGvF+gvm+Q4TbvoJ9+z4DbhL3rlvEQR0V3ZvtT6IS64nV
Qpj5bLtv8n0Rz6cn9AQohW/H7jKeZVL+XmgP1KcFoJSzCp+Ed+FaXPLYUzMdX5b4
xszPIDG0ToQf0Wkq9EKnJL2Wal/SSXzqpr1XmPxVcJTz7vnQ/nXpRzwFVL1MzOeM
fRBk0+9Y8CmqjVGuWtzV9/W1/AsxmWrUjToXLB1yB46IwNt8u3pw7qYyhdtqOZx5
79XpGjaQvE9C+FRPl7CZpTjEfZ5jCkPQ3dp0aGcm2hhqe7sPw02fbkawIJiMCo4s
RK+H2jO9G4k/0ul+3MpkVfXg8d1XRx1Y4oZTLETe6YsU5QivmVCu78cn10qKtq0C
Txn310xVHt2z797mLqiFFrEUlg6Oc13j/JO7VjcjwTQCWPnL8wEm88mfMDbW4xQC
LEfeqYnRs36T24li3CmVtmnFk1+2V5SBH5+RrOL7j3ah2YF0zCHrurbLpsMS9fQN
Ccp/uDZXzn8Eb9ojlG8OPvDDmgLgkYaezhKJc5Gtm0WMUNiqld0uxoVNbBhGcCB+
VClmUvaUAtmQFZmQuhqVfrH6tDksnq/SMkKhChyv2Bd24oXgop7XyrDYF2JhsWgj
J6Cq55eofbuvLP92B708DMyfi0H6vmxwXVFjSUXGLuRkn1gY4oD3Um9Aw7RkTKcD
gAAbKTyNXJvXyxVi/Xo7wo/d6Bpa8pN4qYzPYz98j5FC08Hu3oa+xESqTK/y/yy2
c3lN2yLDaqreMVHXTovTBLmT6pvTAXKVSLr345Mw2vP4QlmNXjS/ZMVUeutpxsgO
JAIXdY4whFMTjKUphWitTC783JMtoh+LET0EVDWYu++yuuMMucZsPxE9GCSqKE83
NFs3C6LlnY8LHaQZc7PWUWpaswCYwLL/uUA/DVRvQe9u+o646W4U9z1JU08YV/uB
/gvHaFDATqIMVFoo0jnURx43VKnQImyDTYnS7F7Ow2rx0BQRMDHeKLr1UvEJNghW
zbWJXDZUej513z1fuKyk+CZxQfO8JSfT2fxbar0Jv2u+G0MkS41OarFJ4CX3rPtr
CIF55WOtZ/1RDqgz8/QlYCJmB2VqQzztuP5cUKiK8wjXepPOhi9M9zsTGdURfx3c
h0EKjNjYclnlGo38eFJNUy388QyDHSV3MP+iQ85AvQFNkr+JoHqYDNCzWUZfFRGI
bkAT1ZpXMJp9Fi+u5KiZVKpEqu+xpsj7OSp7KcqZsfrkWxnnGU6Kb70d53Wo0dZc
Hx8cEpsS0wkpV0+4YeIEqQcmFbtZyPsO4hoqeYA9jm8ejK4/6owLSE6EMFUtyZUM
k6Nj5YmHgryPkrBCAGMYuhTGONg3/kVcAGlwwwnM7LjA3sZaZa0vFxOazUwkTBXT
/vufTEClKVMIG1OiEXuxiOCIC8o73iiOQaWNxW8B/sICLPHXRpzNCgg6tRcbHhSu
DIdd/J5WruDW/ThPRZbvvzByB5HkDsZRMC993IuXK1Gv2ksX1kgqX/nK/WJ8A9M4
xP6oBwiE5i9+/zf7Stwqbe5F5G172IOGVMJDtsTKqFc92nT538B4fdcbcyha/NwS
6vNkkYPlwIirKCIecWavkSkSxyHLdKrCEg/uW0D56Dn+FZp0OV4MXmsAtQDGkumJ
3u6TKggTSDx2U3A4MtZsmWKGAA6zOhDvJHOouSeXzbepO1MDIw8TrxQ6d0xtrmFa
4R/g9kGPN0S5upBr79hHJMEu0EsUl2jmDIZJIgH17dzjjWiXGInECocotaL6mn6X
iKlH4zeuRz8OOQs5EaW1eKFaP4yg9buCWOSldaV72zK+buKvx5ZeBn7RHUY+NmDv
f25mtTqMz29vksXCXrO8goRwcAtkFKK50WG0RFPO88euGvov4y3te1R+1Z7cRSz9
8RtPo+F+PFbjSlxELlAimerN0x7nvzD/tCf20XWJklFR938ZljGSudOiQgY5KQfN
mXW3Wi9TfTcFdkO/Z3jilnIXE6wiGhviQsfSCEXBvdVQC7e0RVJETRpoFZVmzG6w
YNgJfjbP2Q/EvIEzuEj86AT2n2KdG03hO634wTjyllpR7Kp4KsbbtZxGMre55Tcl
GT+waSjNwTiMLfgZ5T3iPuqN4gz2X16Dr6B1X/cT7kD8jha7mvsZGsXT+4vni1e3
KzEnIE6+hhvlB5oLMs1WhlOk6ceJHB82No13Fz2QvCitWJmoSji7lelCnVHdArTU
clFxlL5kSaKRa+F85e+4eG2Nv/WaGFJ2dKGf2zsIjbAJNGUz/zwg6txlUfM4NNKW
whGm1jxa/MjuPahCw+pHj0FBVxNSGoAaZnzu8R02NO2bNC4UDxS2pz2A0JmShICA
7jUZ9saZLFEbljUTQsmDNJ46rWnbTT1+E8RaXUr0USRInRSGkpcB3n8SecPPIeMy
bTDmhsB7TYol+WSHhTHOJaHbWtcS1ADblVrjZ4aG9kVmw3Pn6nza/lgwSF90KCQQ
+Yd2Lg3HaEQGH/QKAp5iD0UVavzh4LQ8phJHLY5d45jT5fOgH6tvqq6ITSLqbUKX
ktbhs632sV+4H+NpC/FVIzbvxTXQ7U+PzhX0LvqqoEysQZAS3xcMGqFE0/YkIc19
YmT805OvGCagTjOtS8NatSAwHv2wO/1sL8T91fQlLuGciFuaA0Ye2Ga98k79nnS4
H/oDdg2pGTYgx2VDNR19zS2gZTpqKK4BINE04C3MbJ0VqaTk25bSwcAIh7rl7Df0
YQ8YipWINruNPSBZJvVSsfWKLqml6QrQplDk82NczkkmtbZbvDaPWVplgKndTAkU
27WlzafC0C+U8Ot/bx/uuusShvaIH/EtCZCoo2Ur6r/1EcEtet6U6oksxPvPvO95
PPDGN518BcKDvzWToS6sSE1Sh0Pb4EBPPHNXRHUdIHjJA/CAhLz58USnH1GbUc+R
npYrNoCaqCT955PGm+ZKRqJPnEmBkB+u6xO0ZzsdylpajREEqrgVmwBGs96BdVDc
VyRpnmQ3HfRIhJ6MZCicfJNMxtewFExDK7BZw+cbp6kuZxRKCNrAyd9/yfWGr175
4qQmhgnfJ0Kp3TvzqcARsw09kuc4XYb//XKwotTYvm/GD4WQgyYy58fT2NlOJym+
HlCX7hhPtNtoLhFeASvJUb71Uu8NcyZY/W/83499MmAJA/aW2eSUsvllO/2nWEtQ
x4S1w0xVUBIGOlkpdptR4UwcwSZeDZRRkU+Zkg0ic2uAJ70qQIh9o8AQ7U5oLL6d
hZ8SWs6rrK6dVRH5LiHDI7D9RWbzb2Gj28rbjjw9dlEtJbuYTaeiGjERXhxLsDdf
Wx50Ln2rKtudJhAj1MCtJVwT3yOADReq30fFDJErtstgksL+gkGnafkT4O+kaB/i
XtOxaJtQPdHwwh93D3dUgJYIfILBcTFwGGvKSmal6rymf5dsZXD0Pr2KvgBYCHcQ
zOV92xasJZL1b8fFMdg9sArrHawSHvCeFGrKp45KBPx3fN1+hNPOBwYc+6Ip4Our
m6ilCgUEEwRNFAIAcR8MrB4zMtwYCsdU0fdLfJQw9XOt0Wpa1J8e1UaihacXZ8+b
MguchBhmzOZMbiDAE2rxpYWkaC57pvOI8IILI5EMthxzC8vS2muuWJedloxjawz7
MDp9cfoVn9+k06IssyFXGZzaikBrjsk/4V7gYWdcj5r4inFK8LbjDnNFdvq/Gn2I
s1ow1jDAa0bbr7wzQXC5iUji0Gva1Ys9jWNlWVBz6jADeQAyZMPne+azX3AQHyiG
45NCz8TcqVu78aANkhu31PnW1rzwvP/iLy2WYA6Ebpn7QUY26+deckpAM0QbLbCc
XsOk8naUnoQrVZ8b4vzwEZsUHylSxsVu+pn/WhYXnUk0d46C8Abt/q/jnNLE8Ptb
GUHHDCgkOiLgqugAiIk7tnq9jbdPW+Tr2UfgGxwFyxIu+AWvbfQUl3BHxOXDqiDb
+0XiS0svMn4hTeJbaY19Rit54ug3k4cHvFls+6XPkY3brKsdJ+sw5rWjw8+XfLhQ
koSyfQR5x+zpqMI9t7H6WlbKKqRReQ0QNYvJmvlO/w/oPCHhrYSwKC/tpEIUr+Ba
i+tpXnYwNSqdBm0IYk2OiUXJ71bx0GDQGY69dHa3s0lcUYEuRSpoOB3/w+9wF6rL
0VJPA/acJxPjGNzMH9BDWcn+y9UMwUPt2WCR51PLfJYpUtQMoVmdEvtbdauHtxjR
11LjfI/JfNcFf21nc/D3WwQeLPj+BEBtfRXp6Vljs41/NmmGgU2O03W2So0h8n5U
rKeyKerDKiAQcXljw4g7OnO3fA1DtjQjbKdbmIs77KYtmGSlCIchxh2uP9+Wb2Zk
6UbcYkWLd7vMmZX7I51zGLgVk/cpEiSfxhBT10ybsB0CkfSTL04GpNZI+w33f6qR
qdPa9lI6crUThFz9o8+gy6PmLSN2rUSyxoxroiuFpm8HyZexQXInp7uUFspE7Fd5
KA5SwZhaAk+bznN1PzVVR3CmqkYEETqfRUgkQFDNhURTqkM1Bh8AzsdswU1lfvqt
FU/YE6uA8qptBjU0Qvosq06g/sodI1Wg5jmhx4A+SCtMCuuHIsurAEyS3zdiqWB+
FVlgGRestgeJtddKwNXpOeNaF9LYe+qlWvuIpgjssY/fU1yBDngU7riTmJFe/Cu2
rfLyOd0JoNExEHpBv3B4d7x1kRt6s+eFEVTdtmIcmeR8V86F2q6lfAvXXsPtH7Na
X9i998EQfOb5KlOM1Mby4jP4rG+0BQBpZJhUaVitDfSxIXMkmWSaNKIDiKIB4H0b
1WkVuZfsgkYfR0+7NxKNKbG++2bMBGVhN/POC96vIZIEv5mV/BC8VTEGCvxFzqn5
2cOnsq7i+C83wuL36QGcfHoI9P7JqvcD186CRFv+rvFYBl0J0KDQp1XtI3uoFfYD
Jxz3P9uffp81v4pNiXHy7cBV89bYTi310uhKaeiAW4DC6bbeMv9zId9y8S7WmvOK
3HrnIJD9+Wkm9k0VgWw9cF6sm8l7DEcncJIPtXUBv2VJ4LjmuL6fwoDrX3E/Anzt
wdTZe6f21q6T/2ETHy9XARedP7zkkp3R9P+7P3iKi31tPUevyZ/ss6MQUgmpluiB
boMGrSsAOynhF0iooniMRw/5RisqIaR9l7NYcxnvIQQzPFBjz2S7cN2SSlUW11XQ
fZJgLGIqXMQIpk6UKSVOHhUqOjwtKXV/jxi7vwE9E4pcg67qXjjzISPN5L3yH3D8
9DL5p6tCxewugZo8X7Uys7mGTkverTJi9S8mox5XliFLgelAXcWTevAbEFxmThZu
armFHT0mZ1YA/dssSCwyoGWz8vUcksEiCr93GJKUAw2ONzDcyioOK4KwuTG0eBw3
tboyW78Ft97sLPiVnk8FJbaVqozUgycZWwmQLFFtOX60JaDw7O4VvZTicETNgar/
6LJ0OIY0t7WwvjMc50aIqWdarfkas8c2b1UFCeVr6WhL0n/ZyZd9r3Q66UCsqvrY
1ciceNBGvIbhH7kWfPyamAU5EVr2fujAyo1E4PntpIYuPFJ+yJRsFRBmvUMWarKB
M/YHXnZE4PJoCXJl/StZphCqKG3EnWvFytj7Ast7wVZdG6FvWMYRtrO+0rnPpVQA
r1bFLtyPFI+GtYeDChiUhwdDYOulIbJQ3HOa1aMAsLbjg8BrCXjABN3qYvGt4QFl
4y7ja5txxegLmxrvMN9cmEshMeI+o3mtkHIfsVxF9GPFrFqeMO4hxrPSB3ugw9Rw
FICrHeF7mkuMTv9J3jxaYEjhcaDAoSUV5sUJWEf7Uehng/DkL6Rh93sQs+sbCrDq
oxRIoGjKn5K1RhFcN9H69TJ/2/jni3ENkISSIdsLhET8xpMed1mQjs//TdeksY0r
3/iLXQeKGEdB1pCp1IwdMcn53QXIkb+zdyePoU3OJxuBgVwSEseq9gdy8wypDnze
gDgZjjlAaSGQOH8i7MBkI/Bzd7HWOzXUa1nLBQje7pTeG8g2tHafsV/+taNW1xgX
87d6m033V41UVox9I/q8Kixy36pbtlBzd7snE6KlHaaTsP8dpdN3adi74SgLMH8I
dh3yFIzSVBgvKe6MxlQyLQXgyirpJBWFYgfwiqnNkj7dvISSgy9HAnYCisyoSZkh
Jv7CLCwf9thyNuGLBaafJ2xQMINeQ0OWQhyY2qMsBrzWitpjRv2BqLIPriw1m5IT
2+6Zm11fuBSm9pWPLO4rHfAq1cYZ7mopJbTc4ELpsa3em4mV72KFjDUN1Lyo1o2L
K5XAjrx07ulqx5pulQFo+u21dKr7m++xkoX+dq8ROfQduWPvlDSPNSxhFK4S2tZF
kHEd/Mpn0yHCTkZEsLyzdgfh5yHB5bJgDqEOlmvsmMsoBLEYGuWTpVr/EldUY4xJ
HuCXhUGRHYyqULpkbWCG89beNQyR5/RWyxFm55ChXWCi8xZ91maXXBfNtFjd/nId
vubEs8OmLX1stHTj0YpWGpoyxwDSCl0cB4/xg/tLvJHe2R87jBMPSu8zOWxddnM6
3s9EAta1qbp3wO/P7INHHexxXqqc8bEFD/Dco3d3JgoKXDfpyyfRq08A72I8kQUt
IT6xUXeuhQQ5CBzbNLAMVSKi/L5OMYLKyYVrubSCyjXTNmfrm+v9SQMaVuJayVR9
zApgNXZ/bedzsgFEBJv+ZgcTUg6uZH8eTlR2T2w98SzxnPBzwoHWdjroYEDcQggf
dEQp314TYtnWtZZeDWcWfVImjPqKd1QWOf0/URn7gLfnNhUlU5TSQjcb/ZfdRZcY
XkudgsRgyw5GA49zt7i2Zu+XXlNlAEneDsEpY+Higm/HF2hrxCdlG3LlbGYPzmvn
WPbSj6JWT9asAcSXfyd7IJwXiUNQZUduNmY9H/oZh6651/3VqEn4QCbGty2lw3OG
mth7/xnOVGScB58WFN+xwEHU9bMmnXlq/fyEM3mVeY8qSKfRn5HpWkfj9NxXSwd5
kb0cRMBO7Z+ebLjGl7tl7Y1kAczHU2gpRyl8AqVbudB2UqMQWD0Si54ErsiDSx65
d1Wlv7lNkVcWnCtSqYxItX/8Wrp65854QdBdXKfcGnvWxFE7IIkV9QJ8R8eLAT9L
DVtdWN3Bxr2PcWD6vtg9sOw5QEd3hTEClx0vic9Ds+/Eg3JmpWIE5KCFQ5UF4Ice
lrptxh3i0PtzUUo7dfidM+Q2JwP0pqQjb4FoPpuYWbac4Y7ItQogi/yOC7ilFWWa
dG+AfgFDOSevEHBXvwWrcsVnGhpPqQgYoUT4a1dayaKruFkG+casl9/OkdiCEa7l
elU9403p3HwZG+3ttqminPZ4orKiTyMrOMgpmTILmj3UlLB9BfE5cW9r49C5D8Dh
6LC7BGlwhfYe+2r4S+vF0qxtvdCKmJEuGVlYv0z92wNap+DXcNf+Pu7YOpnZ7XyI
IilKCDnIfsrR4+5zu516fFp9G4PMcXsEuKgrr3T/yj5lAaTXxuUbsRYgrZdUfDh0
+f9yvgpAvJmhFBdGNOFd1pfjQvw76O24aVO5L2ATAZiP2JkWGKXlXWhUpaD/tgGF
kDcj/+OXi4p/qtfyIfLt2OEEYy8P/xXkFJOgnEfz8KkVQpDE0AkD6rCUGOeBth8z
LdqgsCWXCPcdzWgAr34S6WvBbDj0uFihvkZ3bXMo/LEG8xFojGJR+RP8CDSIt3I9
Z8tyEYYha0K/KxKgsLxiiqwpFKv0yB4CSaigUbaloT9ixlnkmmOMyGxJzyOOVSiu
gwz2OCN2BiUpNFinbELk4hyhZ4f+hcfqs/qnhg76uAfbMhjpbS8sxRGEI+mbho2Z
saUIg5Wk/hXNbvB+V8NxAcx5SZelSbR7JcrSIhE2ZD/aEPxGv3QfOkz0z86kQehb
ChX1VaB6iaaBFWi4h/xwct9VkX4XgL8wKaQxl19MuBtqqIc2WgwmYew7Uhcqybg3
AU1cmVKfzed/PTBra53BNNirNeZVzcMus47YzXkJ53xCvZNnKPgHFO/RnwndKyT0
v1KbetHwX0A/bAL2HXL8Rv8a9ad9o31SzLcrmsylkVEfzKc0fh6YKCe2CYX3op2P
HmXvkZV9zLZPd6593BXDKWtIiKxlLx+fX5n1z3A9h1vunvBmZnvQF4wOWT6ZTwou
z1wDK+w72pmxkj6N4Du8cnBdGxIB7Bj3WZR1yach9XlTDiHixXfKrOGaEJ0cVo+b
NiFDCgTIQcMkzX2ys34OD7FOupX024T2KQcnNs1xhWCja9S51YIDh+4PkIIdKNUN
ttwhOzI1U5QcFXqrleMQKX0883K3XObqki5oEGciKwQrnw0UlWsI7p2inKptRJzd
9c6hP/S75IAUIEP+34IC93xEEktnp9OsyqbW2mw3euVJW80Ylp1z5Jth/tE3udTU
ylkd7Ep3rWCqdHO3qNB8qLIRZBjsgN7A/rB58uLdvgt/GA96lKKeWXJE3TxBC3ns
5lJ5889fw8QlQRneYgizkI1ltE+vSXieCKr34IJz/kfFiwpLcckCnJKjK38jyrWP
bAiWgxVxPfmyb/pnDCuIIs1ivWufRL7/AUV1SJCIj91g6HlyvAzgM3CqInM5IoiT
dyEOBZhyYkRfptCXUiJx8zGBA99MF4xH2og99uGW2VogxJhCxS5lXKG0yCp9wvoc
R4O152MhNCunp23CEte5OpA1/ovy32uhFv9EQ+y4eKpDyNVxnGml9Yj5ki/2CstX
IJgmaTrryuiLKrn2rc2kWZX5jyDQpTJ3ynHV1kRtqxfe4d3f4acigulg+oZrTezi
es7hA75Ly6M7s0u70Q8tLgovlKEuEYieC4Fhu1MS3BXN5KzGNwxxebrwZpMOH4Ji
eXZ1Yj+DBFLCkkqTNdWmNJpwmZHALIVKYWhLvAH8lIAgUcrT4avd5Z/60pV/0VEI
vgFxAchXnjuKxqiaszMzWahelkiz8Lo4++J03bKjkL+szvjtXzuhbKiZfop/lkRU
BPyQ5XRoNsz/Eowi5cQxbBkfOKxpSqUzjq/jgZp+mCGu3a1dJN+M5YmGPhoBGeAs
r2qgm7Cg7I6hMsklimdsvjsDFML77Og4Z766iZqlkWAOUIBgSGuedBJPtOzNoAPM
YnYrUWYB46MhRzz2EFS47cx7rj4ax9KEYBChczoOT1lyhr156Pa992I8QtcBqSi/
TV4PzTPpvUNX1Fz6Rh83z3jvMhFTJIgxNZWWj5DfccBJCQ11mDigwoLygNcZpEZ1
Ana9pvwzMESuBZXM/QrdmKSy/TeKmxlmAHJKZT4AW8QIQCp+r7lGcHNrnMHikDQO
JpKrQccaQLkIKxfGHDpdAevTAZU4PIUAyKQhXMBn2tJAtyySqr05l4I8UPNk5nlx
JzDC7F0RQeTmk1pmNafxHVACKqLj+rJZANCPLA5mqKZboLi9vIChdEP1OybAoPor
FaiuEv2eWyA28Fa1NUdAnjrhpP/LVWTkjxU9snrHSzZE+alhV9XrLbQjbCFQRXr0
v16es1fx2RQJEL30QpH1+VaPirx5AIGz5e5EmlSvEBG9mXHT3p9n9SBQ5CiXi+al
wy/SVhOvN4StvtXaTq6Ffvqr8fpS/+pivvBPhMS0FTFlXD4lu6WnQITOjQYI8Xz3
W61P4PTtCu4JCFSDBiHHiloLlFqhNSIW9UXg+D+lkD8LTmg7RxrZoObZsJwXD8VN
OW2waZX5ql/lqLW3DW0pn4GCqIjwQOgZpLRZ2wf5pae4ROeqtUsJpHhUYuq3v+K9
2DRP4p5LBUUJMv79qgS/w5aautLRCG4SCWzLxs2bzPJq4V9wGa4EHosrnz2d/FES
icddTH4wmanwQgdu/hj1SDIMSPZIuLKhPmgLVO1bAHlZDWdoI5A6Z3BmZzr3yUEa
6i8LvEfANqm5jgQLG59H00m6MxNBk4GlLMEUnO/6+5fLB4Asvg9ydgK56rCOv2tq
RrN+S4e9dimR/CVviJk1VNZlupXLEOpXwz4tjrviQnUe4lYpw88EmyrOxS7+z2SP
d6ejypsNGwZMIIk+QnB4J6wSU24jN0UV3CyONP/qwwRIoGKOzVyGKbjCYEIzQwZ8
opqZOQt6sgSkgS2de8UQ79Tebfd/LaFLPQ4ko9QcSq3V/kOnsGAeL10HSjtetw/s
GRwK3jf3mwujXRRJcWHun+cUYwTZaUaiZBu5tnDDRtFzK7se8sL5BSeMLkMNxTz+
Ch+AZRuAkA8Oh3g1yML5y4y23mSgyr5oBOPIwCfQ0KA/iHbPNo0nrPjHJLzAquQz
W1gePQJ4/XDstYgyBAVDkIlieLOw5noozu/JP5jG+rSkYHyhYCgbvuOLE4NjS+YZ
5s0K8EfjtDpq5wPzbekwSD5EZ0M+qo40gMK/VwsWAcgTsZrVR4R2L95PaB09ULIm
wol062ySB9zDBKRv4BqnzwwRf2+C9XXYFVazCOcf5x+JGRqfqBMlt5IIcXXsfLES
dl3nPLW3T1VNvlw1zYjUDbTOkZLaA5TSTcE4lQJ3qoocU2XEAelEjpf1lI4dAE+2
W0Kr7scBNVPD49w3QwLtOmb7JtOkLiB0FHz5Xcvvz8rGEZs7Xb62OdzRnFPcdpPp
gKz+SKpiee159yVevaHaMU2PXvOKYyJ1Pw5V/U/ZmqPoYz9OT+g7Nb5Omn44XgHo
1zZg9E/uBY7L8T9oFOHARHTx4EzQhIQQRUpsg56visv2JxVLwPrXUYslWjAHCeuC
aHd1xVE64eI/A1YZlsGQE9H07VZqYvlI++9oBojZNc1f3lGRnJGWETPu0e3et756
r5gE2jDWJejRVPP9p53QQVnqZhkXDAoTWLnIM/OFl9ODwy113DP4/srQton+1Oop
51N95q2UcxR3SmMtGUDYjlR0Hiu56c74TyUPNW450KS/nHiHRMXL3vpnfKrozWrW
UweNyUt3KjSymS0PnCR2mhJrct1uQpLKFSeIJ+UY26oEit0q5Qpf9TrEUV9Tk1UF
msGJTZI+4jR8pVCMHhON0mE87a8G/dtop0tRdi3k7EjLqy05jnQI8PcGOBPtSTD7
oDx09uvzYj+r94aS6Tuxp5+Wnukqt1kSt2kOkxL3AKLqgXpq89pp2UycmgF9ZmC4
6M4YiZeOLCGXR7KaHs4fPl1Hqt1tb+oBPY/4tXrKF2zpESUVf/3Bvv6l47EjaxDl
K+ojMigrwv+RyZpbdL3r97cKbh7ibKOjPsHF4PYEPuMI1SUa2OG+GTwOZSw0+SI9
4uPZrqqmQZB1bshaXCwrEnT3NCXBGPfbWl014ziaSugXjmasY6l3qm34B5DdM05U
X+GGgdrUcWBUuZMUBgFSEz4AA0t7YydKxppZvhMf98HalPpkYJtgeXW95uHPGEXF
GrYATKkUuk/TDsKckZmtV23EjHJDgAf61ZKaMwsvYJ+xf6Df+uaUtXg3R6wroZqS
LHKJMf+M0KuUxtNbN1KhS8TMYLdolVUgGTey3CnU83Il+mr4tUujv2tkhzjW0Apg
wv1h30DQGpJBHQJ1iXLzG5uTQKoFx2Bv7z3xaXYdYMrx/3xTaWrsIoFyyS/6hD87
tKMBPMk4GTgw4H2fGl/DobkYwuh301MRtW04YTB2CDteIYy6aXW/D11/CpsQKpRA
47eAs6pPvEp6X0GICDvk1yTyDnP2breAD6W1dYleXG31AFrvcdpVoJtBftzkNL4x
hN/ZcZiVfqpOIGcJbGSvJgCqmp0zdTnoW/8lE+M0eXM6iqg924jo5R24bGVe2V/u
mFHVHfxt3jGNaL7iexh1FiVKrN5jSDZvv63QaO339XZvAU6P6JlZEzjYuHfDYmSM
i+YOlwDN0hL3kX1UvDR/5F6Wb52SJVVXjlWVPTcGp/1a9OTR8t6xNbd1K/nuneFm
ViXHLJaMW9ZfOLUyKrhEDRLinHUEKy6RZM3RcTf8nVDb77xuy5iwhzUwbVaYLblJ
4wosl9+Fa7Eql3h5hlIJ6036wnsaCCb7JjFrwSwZCkX/yDAPPt+0ltJ0jMnbLv4r
nUdQ6beRhMClHiyDmdKuOGgR+AY85ehs8Q0gHOAbTgg3ZlAYmKSZxb2WNkDtATmR
6zStAr003mXqF4tkc0TfceNzl6i1ekfGUijkDgnKuuh0IxILuyABjVgoTneKzR26
KWn7H+RpTPkDQyjjisb2zKgtcIWsHOKZBbGZc6mYsEB12dHOL5F8wtrRwUsF7B+h
zLPiMqzsDuXMZguohjFaELdGqKSHPAlWfvP6X7cszV3B2dQOyIVQ1CWHHJmgctfE
jLgnulKDSRI1zmmobFFSJWHv2jTqfc9dOHMwNcWeECAHLbSNuC7Uex2hzVmLu/ES
A8NETQ2duCibu6gzLj3t5AAfU4xHkp+nFNKzHEGkvACX5ff44SZ5pLThYReq5LN6
xQbBuWnTSKi8gSrHfV2neaWY914xhINPZqGypjRBf26g4NvA3dHyu7qB6Q3JGB/H
9MNhBfBrkIeLhDiJ42cVd8a+H0jHg4J2tZ8Tql6qJoiYFPc1BBJXZTRpNKCT3pwj
sbPuRexsAblz9qZvwoku8mDO0eamdSwquok1rQzNc5u7YKORATAf6gqci9+7qobS
JCj1ufx+rcWHFzSwYrjJypESVWyjqrlK+HfCkdIQ4lDRFqMFuPHt7k+cf3O/Xayc
E1VAPbmdTw1sEtS/8390WItWnVDQcShgC/irUutTBWPJ4ZMnMnHOx2LSaCOhmbmX
xvz6X+EsJawKPDVn3SRZEDeza8Ms7ABQARqYaK+r6wjZKABnp5tWvM8rb3PtXBvG
IiHxm8GavcJ1EFuTHVyUJnZsrBx7xjr+wjlY8l+SflCPewLBZEtA7v4mKTRKQjzD
wDAsehnVGmErCAB90VtCnQjQ3Z2aRNV2D/cIdbqzzeB39nBBJc+gZqHeJ1aV+U3c
I/a5EhYpDPDcYU0/riNoEHvzjrXUP9sLqBUV2H+AhFnPVbwUT4QbLoloveoqGqSI
6fn6ZL3/xZtKdPxupgzMG0MLjgZhxwxvT4hw3TI7y7Q5uGn66Q2Jf/k/bSpnq6ex
HRtS+fE0GxR72PFuuvu3Rh8pLqPSeMMKMCt+cNAGLCyf8JZ+xSTmrZ4XXcjaWye/
FrSJyOJgy3okcHcdL5HaSSUTqI8Vq9VSDvazvHc3sdNCE/zKHOobNRpV2ceukmpS
knIjG6m/1l+n8GYhyO8gHLxnAQM7govRrZE0lljKSLzlkvMKiNU716peFKMRskMq
RFimiTMVwNmSW1837QfVm6l4qKbMLfyJXX95vj+0RD0iJM7S1a0QFXX5hjcLTT0z
bEAMnbpw9M3czlQINlkpPvACk6vISmbCfpPRRJD901D2stgOzQj4gl2VLJZiLfHh
4XfqKJDPwrIDjG20wwL0CvFJpbi83AGTIUxw9TEg6q5E6oWI721dr0uI+AvI5UAR
sHpSlX+BnF+PFHMFswL8R8oOVbNdDklMpoCyuyaYbQoetMnaWSagVIeq4+UKqdsd
jt9s+i4giPURU+LD0lotORk2p9fr2JhyB4cdFe/B0ssi4T4WLKLApx1BHoiQXqJe
WdFgw69HrjyMglbo7DTd/Jd6ikIalGpMNQc9Rl2pfGbTRLn8yBk7wZt3out5ZtOG
fllaoJvlQsWS06PculJNW/s8lUunhxEoRvDT1ngJhZcZ2Hr5OfOkypub23O9kmeP
Y3EynKiEM2Gpg8MEiOp8SGNPy8+xSmxXskqbFGJeGS0U2eWogMn3SuW9Vr7dPviP
zb7c2/Sl/bzcr26uL+28FRpOtedrnxpY8DqRYo5kwM/4Dque1Ghf27HZ5BPj1X0v
kuafGRLYfgEnkyRsPbtNKI3QBf2Rk+el+Ihz7AVcSBPh0HRfCKd/1x36AkjKD8na
8VAPugACGkUK3wo9dsuo70mpJImMBoBdYJ0L/YRHHvoDFIL36NMUPaDjZdry70Tw
Jk2B0zTxDoim5PeQW0pm1MJRlyAIzXFaF66gegVSVyXO7bxIHQMQb6oDPqnM3dFg
BZ4vKSwziSF2mTytcXEX5EzUXljOqTACDURkCVPVK8NjnL711Vl0xeDyr2LL7pDW
tNAv/RELtiMNFZMjYy5DniqWE75pqTHH29Wby4fY6W3OOlUqpiFbzBN4PPrlNe0o
n2QSQaXrgvL+ykKbMoOy4PYnHEBNUIj2vdD2wBA18bkKYgnX++xnu+aB6TScGAox
xdfVROU7OnZB3srDXtfy+Ym7+1E+4zNNFZ15Apwosj1Xj3EYxDv3JBEps+4UqtDq
u82bNG7Dm9Lnux6hHJKlXe3Ws5LhAVU+IIvd1crWQjJUqCZgPDvOoxAKH/09meMD
zbzlX42U3VCg4tCyN7S5AX/OsI5toSGd3XPFAkTBJYxm0S1MwtIPxkj9K4lZKRmB
cAhdMvgQO67qxtvip05Uqoc+jbaHTfBfrcuu/EHkdzrjZ9BdV0DuBPJ/rALobBLb
EjjIFtyBqc+Up5+sSPDrHQrwzKKx1u/KD+M+KDYBpszDs8J3+duMvTS/hlS+xRu3
kLyaf5LtV2YGtXq0uFiPqobVtvEO0jIjkveXJJdxaEZMW+/7Jg1c1UNNdioLUkXf
pgZlwow9m0n5YhFqcK+ZioFG5+dphzOHAlY2ToVYLMj3CiUNxmpRIwX14Gf+kcFh
9bNtRSYpyh5WnsSmZDAd4a2RKSktS+pl2z6ewiH0amLdXGdxcnJ0rjZtsTiJ8o9G
jL+iylg54JHBoYgrRlNPKyVd7TD+EIUb1uxG1KtS+IO/9nNnuAUuetMPMJeBg+eB
Yu3k8vQ598l0nBhYEFcpKrEUjCZqOfUU3jtbMa2rKnjJ5YblzIBc5pEjUBXdCQbp
xjS4Z55B0VwEZZBx8XAkW3yqnUMLJdCwO6Qx7JErKOnYRVZnxE8+SSLodZI+GtHf
7wmkW0v0bwTRi4husHpJvo5yBrlsXmBGu5EjhREpwrdHmX3nEAY6F46/ZlX8lOHr
/a60twNzuHFTCzpUfYQAdHsn+Mbgc0cc0/iFW4KLkmIIz54DM6QZvs+EtW1i3lla
XOIV2DbknR8roily5+wjtDebbqMEbR7m+HSbjJUeCIPdDgvJBUeOe6yRbD1FilCx
g4TIVErWimysiol/z6SY2Xrpz0JekdHGltTwBK3Dwr7ss0LNNTLTEuyUpj7iVE1F
4KhbibwnlFipe0xYjp/hbqIlfFCKF7StaNwpsQQNJoOH29NV6sNlX8ZX/+OskCYf
EjxDFTMOqTjEvpfcJGzb/cEuVubwXzp7esM57eteRtX/QZ3HkQKQS0pRVC0eGpGV
KEvmD0sZUnMfzbQBscrvGmxXwrC4N/KEd3pW54EcTnZqY++xVWtBzYKNFr7mGKLV
88BeyMIXzHuT5VsbcgzaVSQe2rHOuVU7BgQbKHQSAz8AH4MGL+L9TNmSuBpLJpt+
ItQ5Hvohmmn3A9HihJ2n+VrXVWfNWDoF1veFmtMKZiNTpoFzypktLF1lDEzg4u22
pHVuGQvZy1jgkRUEO2zMhVsnIJv6iNjBiqyrPANnuTa1AUdqbL5iTUq4nb9Ek9i1
JzWW4IW/jc1YKW/4DS0O6djNNc+/x9Wh2BVyYKEgWlAI2alWxTyuoK7LzSfFrndD
duG5K3xzMlZwM75v8Fv7hnSuslrm0s6bkPmS3xo77mq/+4iJFCTo8yPtk3rbNSmi
lRgdnEKghgQkz7I++awkybATrv60Yab/LFJgMcKzigx/CeML8SGnlUXh2AB/Ga2+
KvRGxLJPv3mUfYWUn12xLZvSzMqQ0SkXUg9cUHjuk7L5Fp0OJim2dlLogPlYWT11
MWLMZhR+IUkSZkhG//pBJ7/Z0pG5KujdzbngQGB9UHrVhmt+6BIIhK3y8fv+4veK
JjOz4IEpmqddYfjRErWG/mk3mBEe32L/no6W2iLlwaKf/Gm0vvy2JChW5P/iyXX5
797TWry1epNpOSCsugemtDrcb4BUMciEABdn0GU33fD/dQSBlox/sEWyZXrBYsZN
vmb6V7XdQvApko7eRG6GdQNfvpjuXfLWDFbhKigoIh/5lS2DBjD1+iAScCMdf0D+
YIOeEwWd7TrE8WuewJPgznvZr3zKUfUkz0DAbPhonDCLE/0L2qHXnOLEVzevVaKn
j3GnLuL9bXX9lJjzsvPlQZB/5JyP1Xb109nu9skQWUQUgu8+z3ApApdWKKFhcXyT
6qtFf/m7koKIZ9fweEffkn1SF2C5G38mn6sXN+BLP4IHg16i4AHPnNrNkLghi9Dx
P2ClDfhh7XqaQt077ryDV66NA284AAdSvFfW+bgKV4a+/QvX226JM2LBGgzo8ku6
kVLzCx+XAEkEs6mTLK0hja1vqsEcTWhEwOoMXD+yDBB342Hm5T8FAb4nTXECnHKU
gvrifCUT7bb8nf5PasKT7tLXDrXpLiaWJvNLDg38S+n7neHxARxpEIR1hy57ee90
enT8r3KlALo++9xiIad7QN1wN9iV3+UFar0per7IBUn3dE8jBolQSd9Bl6Cvg2U1
ou19yo4hnpBtMciDvQXSdDmfrkQ0myhqDYTmPjUh0ULBMiMiyemPz6YVw5YIp+el
0uXsC4hAB2ty6GRB7FrSotzRggLzScGcJFJ8VfvTNVDxbJ3iP55fsP5a1d+6dEFS
iWbREmfhZcdV+leKgjHkSWqyXDeN5l3mWOVbRjxhpcKILdgGPdonL6OeHqK7GlEF
rhbuU6TERsBkvXiyaqlstcoJcV37459+T9RPQUoWXZliMSeZhHlAjRd37U5YY15k
Ueycb3dZ0XfVf95FkPaLFAvBKpOB4jnRQNF9uqfOfwN0MDxyLVxbxxOaHvIhzzV3
oLwsanyLCO/yFdMH34x5lMmRkKK0nUt0C1O8WihVBWxKDz5MvywxtmRD3Q2hY+ax
pbcDPM8wOYC8yjHSU1Tlu/RpwRUju1aiu6ZU6sf/8ipIPjJfCNWtuRdn8TsMUzpX
F2SMnemMjQjXBnQ8JwtWiR5eRmvlq/F98JyOhpPcNMby6saKeey8UKqhdP/x7cZ2
qERKClflDWSBljPm62zGS+aCkOOPubJgL28eSiAHaC0Ys2lZgQWfl+yfTuRhAsEg
WGkv4+ma3t2/Q125VtT9Nc2ctZhMHUxa30kZ6TFRrO7pfkDjG/euuvXE2bvXL01X
Nz+E4Pn6eUqFiWREpgS8eFVniBAFYFYoFgFl2jsTMut0HsD6N7HVGd9fZXsTV2T4
iotxq2tmO0FRAYBIjbpGETVcQ0ggL+++TGSh1rxxw7JStgMSbsbMgCqsFetpZ1tt
NzDVdy+mVzBsKaRRDuTViOItJChn5rQ634p7JCHbGNrCt75GzVU3syGx+GqjN7vY
X4nBihvXUFAQLv834RMlWffcCitAHwphCrsM+VOx28BXEsr+o1BolDwxDS+CELE0
sqiUswP5SbJ7wGHzfDgo56tfHmFVuQJyg/umy84RjEY0L+LnhmzsfyitAVKsJuli
vKUHY35A5ZGSkRKqdmQpIkxBnfJoZk0mAS9F7eYJpZFdzpseSLPLuqNWUb4lU0sN
fMh16JL/TVrn9uuXrk2CwI/YL7xLaa2daOGe7FXGpFsDgZJbYgH977m3gz2/iSyg
g47uwLr16IK9SGbLkmIo3WKqxKSwPcNfqjU4xJhTnvx9GgazCJGoeTEutjooj1ma
tUxUg6Uzi2U06piTVuYOddmvV5qs/dvHgGaOcoB0Drb1hCmH2ltN5qTN4u7rke2y
0p3usONhk829gW+QuPdQxzC7gBLFUxtcN0GTMM/4VfWXmKjc9URDwlxdb9ASIQwJ
rnpd+9+j4ugEkZWpJl/s5ihl9E/3/DAmw9o7v8iT+9NI57asXb4U0So/Tlz7BY6S
rvn9PnI+nPpLiyAXyXyWhuEvqBfp7y9MxLivTyYLgXFHsqVGq8/F0y5aaGw22vfC
T7M//qV7ulOLXkwj8wTLMbzjBP2TdMXPfrN8Ga7KjirWJnSrUzqW6ZqwJ25a97e1
l4VY+UgkcDlK8qtwxN+sQxwhW9jyBD4t8NKUqO9PkUf2m2po+veGwQOQcFQYGysr
ipmt1x0Gefn/g3bOIL6ekLHWqvFcE2yQUtG415U70Lx6DortcPaSyrIDmz0tMdAx
1pz93TgSBKRIMePT6Qpj+kdAiELlc7hVJunK/0ZidFp/pAcK25a+vNqS49XetXHN
jPEZJO5cN3GWZT8URnP0WLvCXHbAKxya5/mkO9a1ZzfEq1T/73znww9fcvitzhxs
pMkQqVcX1A2x0wlvhyDft5lewftGSkRR7roUynEyVfW8lQoe4CKFj1IMPYzdH9oz
5BLy9QymvIR3RGSPfdUkM2+B6VQp8swpSLxWetWRr6Kn7MLQPmpYTOkIvilyDKyf
HtBQmjAfdgjtYj+DA1m1qoaK3kGszRHe0ON1aeT9K3WCMFxAdFVxl+9zkb6w/DZb
RXuocOCHxzcCdeeCC3U2So7MZQtjqjA8bIanP9juTed+fLwI2kADiTiIFKVZkAEr
tovjVK9A5JMs8ztc5UMwU1OFVTIc/0WtFMkGPBU4x48adEq97F03LTAfiYPMEPc9
L7GIF0Ft2u1KMh4Fdmgck3oHNQabuGhdArhSnZZCtNtNSr7A14OuTicz6/r8yDGb
Kl+GuFl9Cwb1EcjPx48FoTzHR7LVqZ8wYvQzhMt56Ch2VL1F5QlsMq3BTjN4tvnE
B8QBi2jPMEpyYrck9kIjzIOOE5I39se+Sky3SFqGybynHjAQDG82YM55ZYDmHs7w
sc/Co6xh8TNqW2Hj6S+BKh6nLWqaOk1KrQIOOrcyK9T53jmMHNiXCUhjtSQjQ+sj
tTWmw/wVZGYnHCAmBqLJvBXeHwjXx18SAa5iCj4F60QMjHAEQwlWNgkz0SRfrvIl
LYbbMU0xIxBfrD7xxP+4JUzMbd6uXSE07f0vGCnyvumI7fTf+XB4Ik3YA3peUxtF
w85SK3Y3zvUybKBI7WxjJZ6r8PCtbGOp+XujlidGq6r6p31rjRC9O7gWcpvknP7t
eKj9H4NumIOB5+XeHeym90w0gpdXFCuv9VRh/EPOgwa8q8eGj7MH+U1F7/VIXcx+
hBI8iOJTZ7x3E//HbvT5516Jnn+VImaIhksN2SidLbHNkBWBZ1qpXrHA1hqI9WTa
4/B6MI4ZClhuPbi3Z8M+zWQzVmrdJ6+k1edGF/wU9lbFTv2RmYQgn/WlDbQoV8bR
nT02bEzTPUNl+N/dJfhQ0HlrbPTuAWZwbV8OauNUgrFRkfi6G1j3k8WAo2gem3HO
u/hhjjOw+76SjczasvAS3bdbsSGvIcCcuo3ULhNcvtgaLjDdC8pnROwLC3U2Y0WH
HdffOtW2VYvgyVuwewgAegOLjBJpeoSlOdHVIfhpe8mLxWAhNK7f4XFtzgznNL+g
2EP3cwRPzlWMVVPg7Y8sGlwbcN0ZVTeyO35t0hxKNefy1Ii1cvDmzev21PP/IrIo
qzq6JB3vlNerT5Y6yIrYm3wXZxlzJmArMvK38oCpzROnSWhE2m8pKRpnDRouJImw
8ziHosy+pJni4moYh6Qlt0U8yZ5pgHTfu2inwV11RnqMkWYGotx047EcZV0E8Hts
ics2w8wCnt2XmXhgTsYHVgq/RxS+yscqomfOHPbZSwv/hGNbI6cN9G0yLHl2oIhC
DUYj/kbDAw8VpIhZmp6VgR+tuPwd5Yomjj232oCHSEDAoihJD7UAHgB/CEO+itfm
S7a0zqCxJLRAnesYogb2cuD/E7vbL7QS00dfsmGWxgJGgpFCNEgO1EBZfx4Ir3rs
zkI7KBIq6NGyf9nt2RjtvLaLcviUb0ssLXcp8PLHFZ6kwxO7PGKNS3pU5WoFizr8
f1bcOH6e+3sheDEyGuWYr6azHm6mDeWw7dQ60U7VXMrPf+zIltspubP3FK+jrOTn
BmoC6TtyNQkJxqTkPUi31P9HqzGaEspY351zgwwUYHXYAq7FmgLF9HMMsp17Uz2n
eLBTMM8F4uBj/EusJmKIWVijfUXHzkOJtxjZhRtfFC58JVoN4aDDDJv2DxveuaDE
jcmIiLZZpRBmjirnI0W/1HszYJQJ2ZN0giJRqGc7HMRCfQUV7c/fPweh+7lZDiEi
eKJsxzC6qiJ2POToALguhlOZXj2U8ref6fj+0F/cZtQCTkxpcgdEIppVAqTxd93x
XZ5eXgKoVotpzOfwJKUUyYIIwO/vuNrX55WyEO2t56DO03aZR9XCOQ628vn51hCX
4ceHb8Zg4ABILLbakSSvtNZHZVRuzhyWAD9xNqL86Zjkw8ix8r8RG35h78WRBN4D
Ov98UYdiXthIKwkvCU27V02Os+fsQJLk5R4g3yAq2uRQdG77VycT/AYI/Xa+tM3o
QSiYyITKt9MBKmc9Yuwxf9erUUl3PPVlb5c2hvn/4JsmA1VNVfU801I8qRgkLMe/
XiIVhZLjIxN2XR78wbU+0Afi/VXFKYSOxTEXrifDiU1JegpEsDB3NDVFLQyQUUEy
oKtGVIwbGIz+KfzuM2+PrjYMgPxexe8/10JcHRvwOp5krjPu4ln6bnFe3Pus+Oud
OOXSVug/V4BV4pu4F2btTCKOlPvimYsQ+xnRZr23TgC2iiFKUmje+UtFRQ+rpcmk
4S1n457lfgQeXklbxiAqRs5r8EoaO2YhSue7IYHPdRbZVPIF7pYC6xFjoYkuoMTV
As0E3sMGVwZ6cQ0nFbOeyQcKSph37cYbxt9r8phCgWi+mBQSqZR3dwOK8O/2oKR3
79+3C11TSDGxVu6h2vMOvdfF+HPW+tQN7C5PDeq21Jb77NB3KMpJOhbrd1bdk9yF
XZW8olph+qUWdrbCKatXgLD/5A3E/gIwm/q8/rKIHRtvdfEXGI4vh6Hi6JwwQ5jy
S3MSEZgHR9nshXblPTJXHLTgVmGs+DyUb2WSgDfleqqwplz3KTHlvMhOB3/21jnu
1n63PcdaycE/23sjDG7Q/D1+fH45893/4knZ1haVdYjifd1rltYJtoH0yJsZ6Dzg
9xGBDy1WUNSugmMZ9aG2PgrztiFT25ljB148wmHCs1JRShPVeowmjKlBLUs2i1Ko
8oAugXi9JdxTmzjhFlES0oyCIWvPvQExCac9yULzYgmKsSKKPpWVLhAh1fM/KvPK
qackDqlvVyTnjkEdC57ciKYDhIm4ydrKrI2fCoi2ux0eRrZrob+2sd76Q8gt49mL
o6hp7dy/ejTBRV5Zge7Zq0aTgtpLk/XKeK7ZI7VULN5aCaOVqi4VqodshoLeOZ3A
eC/yLhi8V/XtjP/946Mh4ovkafzDpa2WaCDF8PjkcJAvSHVPyySzh9/Jra5Q05xf
BI1uoZqeEL++56MPPB0gMh7a1kD+JTTZAAxmUEZWM2lphmJMVF+Wwkbs3NaQPvaK
XzXyQxW1fEUhw1cDhGJlgek6Aw8srrkpXLkpLXokKjklJDgOQhfZ+aPEdjtSfa27
OqKvijzW6Diy424gRhk8lDg2jXaLOyxyOXoMIho91iCvoVb+6Q1b8J86peN3V+zE
JlG7YWrWiRCyQ5qtFcG7Q7T7i1qU79Uk21aIldsdfq8tSIFyy1QoMgFzMEtfA5Au
MdW5a04PklnMWyOGhcx5JbM2W2fq90lxSMTMz0/oBQTrvXSjdJ2+NB9dcg0yCg+t
wGNd+Ni77qMmJfUqJJpnFTrVB9Dyfd2vTd1LFpVkGJzHR9jxhO3cUn+6cCh2suBJ
pXLVoqXew2Kng2DlqeNGZn8kd0lmYqWNyIT+jUsD0i55NCM1A5Yxv85xMRYlGees
qedHaCAZq8hlPYyGrGS60y/LQQrMjMFe/figkJsI8XTWd7+lhtDhmdoBDOakd+iT
xh8Fv/4kt7alKrZU9s1mocSBX2GnPXEHqnnUdIZH9KmvyX61m8qGTxoUtxEW9036
kD2lDlYOqayfA7S5ttOBMRixY5mwSwIqbTkTm0I2Z4dFO/yOjSTbYsgrRTFvb0N3
JifC+wU0/vTJFT/iv22UE2vzwBCg8mRNotH/Bd+JfWScKagRc6PquNYhs5pSA6JB
BcQnROQrLZXIWzp5f7PBUgQHu652+TBhKPlsesp/DnpWnmlmvocBLS3W6odQm4EB
KGzkBHYQvEyxptb0MqPcCAgVztkqh4wVVmd9AoEuI5qRu0jqmdJvrx45fIXqBcHL
3oyPbo03ejM0c6x5uRphveXZWmZGSmp1MHQAm/Zzj0/vp7yJL/JOPz+O3aQdHkz4
YNPJ0uSLVAt+wtEFHfy8hDZ6Sld0hWKE4uCsi28B3AgXKMtojwdpplTDFy1bVWJR
lL0m6vVD81EtSpx55pDo/jB+KWDEOnuT/4roMSBwl8c9a7yyFV+QGeRMXjQM9USn
34Q7av+/nukAXZXBrBMte02OEtW8uEhNyY1ZKctSMT8RJW+/bTBDdWPRaOIKkuNn
bOSViggy/yh0HUhS8qINdh3cXlIxfc01sZm8Up4qxHaKedl4I3e/gbA6eyAkzLvT
XQS1EO+uWHJ4huqxm4ehYqAZxoac0ulJSqKuPPUEBvavGkYLOC5YpY6dFANbBeYU
UqevOxt+6KPnJuT9+kSdkUuFOmZauQVcm1fbbbhjQ/sfpys/LpS7/SvZkrHfUM26
S3DR733NhW9zI+yKrYVeKSAaGk3CONLOEMxX4FgRppk2tenzORL1HaI1M3tI+1xv
Akumpd6M+SLMBRUUYHlXjz+xVf6uJcj2kX/Tty9yk9ZGH5l1LG//RCUVwulbJMQ/
kb5GtMQcD+abs/WiBOl4xhRL/d1ohSTT5n2GXqPiZWvty6MDdaMQCwPKTmj+aWAl
aOCldiOSdG8h4cu0Fc5eL/WayoS21GUYQjzUhiGlMgacTcrPC2eQa4EqNVUDu5HW
s+xmnFtAO0qyAYCS+AntOeMsHE15Hqb1Vud9cA2dtxFMwXor5BL501HVReMDSNdY
hdTOPTLMKRcd6AuyTab1JoZzjQVQeCzR0HSW68VnGrJ/wZGJRsV9Rr52qCsvK3UO
Dk2/7zIqFXuxTS+w95Xb6Yo5XlB9xiWd4UXcGVN6DJf4LF28N4VmTlegt3K7tO8H
0YjWhyEWq0IpcV1O4EqLY9dGno81kBYS83LqhxuN5je4mqTO7Scf3Vuo5lejJESC
h945/A2JrzQLry8U+CFDeb1kLi1z6yaBHvhwIOQctc2rR+DDe/+P62BnU0iWJedD
o45MTIbuft0WUB/j2jzUDmY/jwt5EZM6qnARTY8EzKMusJaGTqQ+VkS/8qK9hJKy
d4HM0SST1H8711356W7SXthkztdizQIVsofMnHNIVSUNhQM1oor4Kc5xtUykbS+F
4//D657YBPcj6Ew/5Yw9nvnCvj/FbxcHeVPy53cSQwDk2vC40/BJb8k4ydHKKcF9
H4uMVf9kGbydwez4QQTis0IzBRiU0zW98/tL1IVK97uqwF8dC8EXRqaoP0oyLygS
zIHHPadsl4IAGo36lFJ39nLpZGqbCjB9rLH4wxaoccvXy+b7+kWj8urT2QGRLuLy
6kzfCjqtjA1PO9B8z2mRW4XKyz+42hEhn/HXUYr356tgNozbjbiZaxwCWzEWPbmh
WLJokHQGmyJqdx4ayVZbwG0tzqbrtzDlmQnlANCzW03vb86QdZFrgYAPtPMfJfHk
V5ZRKN7td1lpLBdrWSoiwYstQTzXkxVWV+h0wB7wPh+q6bm1KQCz3EVSi22eOKvg
I5VEc6wUF5xZZmYNnXc1v8Nin/DxYo5jfn2fui94khmVU5CtZ1rogVusrLILH54k
PGFrYRRTB9ELeddls6dHBxdJaK8cZcnJbWeYNjSif5KueoqzCnJudLbex1TnRl0+
DHZ/R0w7Fl5YZmxxsQN/s9cYjmT/u6lSyKJ9xPx5ZC0n8bSc6l9h3DVuFAthwDgu
z+fRGK9UoWpuW2K2i56UNZgZ5ocxo4flR+i5rUt48LOzRAX4F38ltGbkDeqSHSMZ
ryZOuI4ikEbQYMH4vk/HxhS691P3yr7IvOg3NoiDcOSXkvDYqf4T3AN7+DPPhNFL
xXFT0dryCGaXnRVwq4fzqjP/qO8JXeNdAiMoj/8mK+xEx+hn1sIppElXw5SALSuy
5XjI9NFyhNKB02GRczkmZd5KTyXGN22IKltTs+pZn9WHTl6IyKno90ku/YrS4E13
tDDh5lOOz9NG37R+O611Y2l0nBg2k8ksMhRco3LSk3+o2eojldQL47usv8QlCRXd
eukeDdN0h5LmiaB07vxGeuEdFe2LVBdLahRpjdj+QEE8nBKMq+A09SEYgz115/7K
4PDmyYGcuRSEfWpulX8Dndp6kpu5EDj6uQmndbqmPXwpbZRwAMr3l1VlC4wUb/Km
lNHU9v+TghoGE9qOOiUIiVEN0EBN8Un8YW0tYQX2o+t4zolfuNjba4eZVbm/Ch0v
ffqZrznFLMJFyZjvBoEz9n0VOQviu4MN6l5/MAI661uNi9nRF/C864cTosx7c2mk
clXKhK4T6VDYVkJ18L5/ii2TRwnE3lMlXhD3iPbubfHpuueL77RuRYeIzNxJKXbJ
MKhxh+ymUAmjykz+qMBSbOO4KTlWvAaYwWISfwUdawb9f3EoBZuAP1CMNCpfSq5G
7pK0mun3WJ++oHMO0Ex7OP3uuojS51X5VgnOqo0qARRX6/pWbhNZfT9tQmfQpEq1
vefeszaItpikw6xRKO/vFRY46pVBwElF+n/bWxouk/N1L/2oewCUYHB2AVQyODsy
86JLOODSl6/sOxq4Ow2IEWxJmg6Tu5lzZgkeMuts///rUVnKbvCDl23W2TCTpGQE
oAybbCYdhP8NGGvdDFxndCRdaphg6Lk4zxM3BmYCWo+H2HKKLOE/lHVbd4BbSiHL
ZrU6cMK5oYGc/KFAD+HCwo78BRc+8GLZJS8OTDno+R3ufSElDw8mPzHYXwN/koex
p/QllkifX0Q2Xhoqy6YwOxodGhoNsWYGuapAKt/ZnSki4XoXusEg/pzoWYrmokfQ
0LWN+5UB8qOFMIOSxj0luKLbcY8X8Ef76j8YPkNLUGSu+puTBq0dvx5Qlid+YS7X
NLaZx2pcIEbefCKED+pyt5OXSO6rzhGndmHxRrxoUpqKyQQ3hbZJeINZ7FIRtVBu
x+6q26roZIsOxMvJCpLv/l6Y9xaPprhWTsZi2qq8h5wVq0c8ocxeSRuNVpOJnevd
ntSnKSIg5ay7ccKbUxc7TbPk6jzOl1QBwKyK0TYRboQLpq+myZ1GdJqi8qD/hncK
YbD6yn3rX/v0AAq5cGmdI1tZT1R8dWkk8NEVJ6MACF1JOdlu+Pg5jidsbWEVC/J0
JdV7hjcgSrlhLhlIfzS88HjENmyFgUMEtAvQ1Jk4jiJLglFvIPBB5qZhtUqTpRCo
eSgYA7ESA6liXge2OQtFnvJ0alfmo9BI0YYmz7aQvp5u+/3/DHgxalDemjBdTVRZ
yAOwXuYcvzZrJLJFApY0pdJgnJNeLheSoefJtpC7jadEcJbp9jd267nc/VV6dFbR
XqJFJvGx284iJ/MMSih/J+DAGzIwpsdYMHhEykammRvkgEAmRE5s/xh9SykdmLGC
63ZoHU8i8hfNttH8UFH+2aIdfSanFd+4Mll/T+trhNCPURx6c2/zE7m7ByOIZXm/
bVlXM4JALEV7/jxH1XMCKpzC1ZidIumyGL/aCfQtXv19L3wZSJpvuf3pbypmWrSy
MlfoqNjtLmFIgbznvYrniEZ3h07hpGqYC4F5UQMx34urRIwkzWzeYG4akT+HFXBd
xUEymzskUQalwfRm0A41+TwBGjm6aWNoRTqTvIESzuSlgUZyLEk3itKxUF3q0R0y
ILEOyQ5cRhr/gOi1G+O6Z6buCWxbcqOxYYpte4rLIc+sUVVnmIlLRMBCk//5gRWl
YlEogqbekSxXOPMekWcocdSsUxBvBLzhRQKdAXfMtipd9KFIC+pBLaVFHF2dRyKL
ffYbD1+jV65LckqtDGk9Nr5T17KtWWbLg73IBR9jHTDwKQ2UKOiLzII5Y1tDehxQ
NWUOU+j1qpCTbwdLI/JRvIgKGkg9Yv9nVkI5GGtUmZbV4XYzj30wkzjwG/3d40I1
B0/jDnFpsmdspqBDT6q7wzGibsWMxtlY8AdqZfjRxCkwbu581duok1z2LxGeVTZr
E8fol5A6g17aPJX9nKtOmPtCYwn3E9cnP4NnpM7JaHyclShdEqYFxFeBMQhWSyKH
s/ia1O7mNqJ4sEo/ep7UvHfjPkW8cQSQAZyR6I5T5eIRIIXGVB+fSm3oNFFJ5zMY
ofp481a1d7chmhndgV1onax6356ZQi7uIWT81l8o0R9fINJyn761KLQ7k33eyDik
1x7X/C1K9haDP7GNtroOfeys0i/BDsjOqFP9asvVtCsSC1319UAsLm/jl5nfkIuP
gSujTmjNUcalz8xNDsOq6lJA65o6Q0O+Y4whGNBxwzFoiKgyQCP/l2ZF0tIGYc7C
aVgE5mx//zRNiGX8e0EkSO6V2uj0O447Q96SKf5G5zaRQvH2IHgvaU9xJ8psZ4dT
Y3FJq0U40nxX9IzJi61vdnY2AX5qOIwJLOFf9x1+MxN+D4aSZEDayul0Q3bMy7EW
M4UjmdJ29WRtjc0Rm9WMl64ybHxlAVf7n36W2Cb9IcLmBdWIXUjVTXKInPfILcnq
acPYoAxiSEy2RvQSQPXM2uo1CDXsvySrCMKxS269TJfuqM3c2cj6IVovq+Byyeeu
wPhQFvZJ6Mx/1FEba4gTzzNV73h9Vs4b72RJyLoPkTLTddMFPFMXpCSYCS/wtYkI
//TNuy0nkrjYb8naQFLThqXEGhKJmAFgY4LE6O7iHYR2jne573jmFvcEA55rnrA9
UN2w+5uLDO6wAA4I2NpkzEQ95jbJ1mb/Rr+fyfXQJszBO2SbUa3BXAUI6lCEg0tj
C3x9kalZsxHf2DuxtP9ye5qguXGlXLw7E0tfXx/aoYd6QG5DC/54mBm8yGJnDENs
BgGDJcrskaswuHJqvNvYqlZVTeqGu2kkId0RQofOm7nuYmEl276IMf9UnuLGrP9n
iy+tbmeRjPJ/eqmMbdRGKz7IJujVd8cJWBSI4lDBtnNvWtwk5Afxc4Fd2EmG/Hu0
kpjbwHd6cPOV8xtm8dmjqsPUyX+FVJECqwtfLkfhK+ufqOAKTC7d1bamL9E9DdtJ
8zTiMViYk4Yny9zDZlfXvdiSONuWMVZRG0IGPz6eqBUMOKIgM7aMnUBDa0zF/ljH
MCTkVPUtKXeCb+7OAZ6b1FayvpAJd9LvXTIbFu4GqVgBmhKZQWAqHDik/rDSN3Qt
W4aLqWWfbapaHV93Y8oKnV9NrONOFeslzCU5k5IW+rVKbeWx+bKxy9+23TWCDjGC
X7uqnHPl4s51nODjFzua5lbE29KjQ3SOLajEpJ43LngB9j4xL+J1JCAcBAu/piQj
N78tiBQHGAThhEYmhairoScodegRqHETAzchKBHnzpgRv3Cd8yNFppEs0K04Kp6B
9E3urvxlvxvE/jAHzHe3AJQuYNTtkt+slOXf2T1BLENC2q00qQ8ep6yIpots9ZYY
HWFwH8L7DcXW+Z3QOjwYpO/vUYxxcX/fI1ruBHpQ/m/Zjm9NL015vmdb36GuXfYR
PCBY0H4JhvK7SrZBeFfNDiVGfaXIoTxgdLRu3PEM6ylgisjMLhKQZygA8AXnEtyF
F0xaNzcnCOxoI1cQYvAtrtEVVeVqlUKv+8umZux9MQ6k2zjC1je3K1lnDV0nvMZY
0dQs0MSHRTcGPvge0ScWpV0ZxBNI5ozm0EavPhFJlvinjf+Bjo4byHq3uQagrefx
iJWKzsFBlQoZu9hb8cCoMSL/kjHijBqvalhB1CimLmdX308k6xRA3S6r3K8mH340
h5XW8kzlr4qc7IM2cXtuNcyqa8MpozeN1I/HRejnqjHiIYbvWR4ys6k49UuT2bRs
Y75zDftD4xDNrULzMTbGMZaYoXKycMnsbwm4mPzDVoIf22nqOcEFw3M1h1+XTBMo
Nq8LweP2/COWe+En6DWi48VeAjdy9GF6zuh61U9mxFGBPosZ3GrPkU9MIQK7tapE
wnwRtU1oI6l/KPeAn0kw1OTkHEJ82XPa26JZ2HgYa1G0ZXRHaqg98221QjnTSdqI
xSHG1TMRUIws4CdB+X2my+O9YyhBFtd7b9RGSQIrBoVmcmsraodmwW9mlv8lxFe/
bVpPoGGgx1MKrPArusw7OSk21KZmCIHRcMAsUFnZ4BvOf/tzZTMrpNQwpS6DEcSo
mX/QjAzCxo7V6e7m7qGqWTrthT+WL6VQKldVO619Hs/lsCopjzF9Hs1gBrFMGuC2
x635MCXalATDeKWsI665EqBjyyQo2w/d1nIKZhA85p7FBR2h0JZrIDylZfzedfFS
VzhxlrdAY5bu3irU2pByyTogLi5JolozRZIXHlxlO8dhavxR1FiYGkbxel09UuzR
FBBM+Y4Lw3wl3foHzTBuJ9CF48b1wTd0IiUWv8KPkFN+zDJEhykZQz7F9LpIh2ey
z/sUUBfMO6kZB4yn2e4NAmNRMjZlkeEmgan6JgZmEDofhdAEhNRUJolmw16mh+tS
g+iywb4ALgK7bUnLLSwuTjgW1zIglthjCqtt2EDcv2dRSaPPAvKadfFD8x42qeQr
tJK8f7/G8rMKA+4XFChNQDDPdRF0y/g269Q3uOzhuvXvl49NhhypWfRtM+swXWzn
ol89VdHL0t3e6tE4BOete5wTvOwDcBIzdztObtij1375Su8v1qhPwRK7uKXyoPd5
mTsySSV8I+qX1xLnc3BS8Jrk8A25w2QYOFPy6OXo9lcvDIeXPRV8dguwEwnmAP84
IoGqQExakLsTFb8EoA2w+xCoHaFqt45LgAkX+dISXznyYCsC6nFE7csbGybB4YMl
b12nuC+hW0tVk8ibItgeqqOIjQwkvrJWfCeox+wUgzf2VBbxx1OG5suN6XhIJVfj
eZgSu+8K9PUSrjHPusHKlCTIqnSaRxgKMeq9mMRzgrZzUrbm2lyMq6x0n7GK9+Yp
nlRFLuvGQayNibZbuNKY9Nl0bYA7gMjQv2eWgAEz3AaTGfwJf4/7T+SyJLi+Cwab
MGyyfHed+rmBKW6k9gJNe4ptOniYbPLu6lM7BkZ0UwwWrhPoE3ZQG3fwlP9MRtGu
jiGsIsNGiJiJahxUypBXNwthbT9FVmARbeTnmymjJbnBOcnZ+xJnMS2tZRdHBKhi
d1cdfbK+Z4wVlTLQL9T3tYZ28LBZWYOMX0vAmamGJ8SOVZj6V3PCpUn3vM7lg0lQ
KDI+zqb/g3V/5tZOFguJc6qAG6No2oTbWF8zs9U3BVjR/cIkhwljz5kmg68KMB0T
7JVnkJCTsINli8l8j/N0svKccw2U9oj0VSH9JXYaWzcV7lhUxQd4sjCbB/HnVt4Q
9fAzo7WwOI4FNoO9Bh+GEKMuNjEUw93cq9rulod6VrhnFqjl5O+Y4FP+fZcaOAaj
tmVGtgzHx5vGeB80fSgRVaf8q4/0a6YGQe4nofrj6x22vCr+y2IjZ22PSDySmWj3
CL8IO3Ob/oELCrlIgQiLlltBs3Vr0gd6/ntZpFGJoFkx84wCQeW2k7zATYmn25rB
2rtszfD/K8Hz/Dqxni8Gs/2ePLjCvxWF2FaMUjxjYkAuf2rZpQYwcC7ygbcQlJGu
f2ks14mK4p7Ith5RRIlBA7XW33ZUUH9wRj6uCHSYlG0LmeE+btueeiTYw52h9NlZ
NjGJ36V6wNfelAM7NTED9jGMaRY5IXwX/R0/5nXW63CPaPz3JfuzHT3LRoJgpVx2
21AqrL9LHvT/8+Dc9loMJZoGF93XdehNFtmhroByQxIhm4i0h/sxi65YMutlDnSA
/8bAZQja9TBx2XB7Uy7/WMt0BR9/fWTcMKv9W03K1LMlneR4U9LcEez847zH+F4v
fUFNI1mtW3ADQ285AMMAY0Qi+ch4OaWFygFD7ayD5Dk32Z4eVYIcG9wr1iOM/N5o
2XQsYQIdE5W3iKpTTsmHdtd8zC9TPWifjcYh/cdsKWPiWp+ST3ggYZxJRziL5FHz
PR4AGuP5RHC5UvVTjQg4L0eOb1WH0KHPXkabNTNYiOF/OdXE0uV1BI0qZasAW8U7
PNGR3EUJSQx7ZgxIkaKykxyUYh6JKv+5GpPrYePPYsZ05j3qWjCl4AZHpagkJvUO
tdoZ2yIqn3roE/PMiZTjw5aP3kQty0mAF7EzByx03xPrfkzqL7BbXozmeGv6wBur
XCaReH9vda1r1OJVScm1t8M/0NiiMlo9hg14Wg8rwD2/crE5cZuUYL8ppj3rUujy
mlc9u4AVpvjG7xHLs7xzn1DqO9C/J/U1IPhN9XlPMnD5kuNi19plueHWlaEzc4h+
B7qIMucKaOtWsopgStGLeGpOpy1mfuEZeZgjRcyviSvyu7dE88ZunGAzPPW7KHSz
LtfWCf6IukB3pf8SZ4IYc3h5h/L669+i+wIapY8QxXCyo6jU/fQtYA3n0kZztvfs
0jk4FeW6f7Vj694a8LTsB9+vUbqe8Qxn+pFdbuvAq3LthGtqqiG/dB98t5gU1ciL
2OKUlZq0CAmgGIQw3b68b+gGsvLb3qRXPWbGzKlm8Nt1PM/xlJh3s2QQ3g2/q6Mc
8SiQ1o0rGdLCsmljvMK+IdlzATgHU5be1AlX3yfnylzZ7BxoFgn0WMTrzl21/5cz
zMBgNzJ/hNZV6QaGXMGUZkHkVWM8eZAuhiKAtU3eQ1FwRfSuVm9YYfHsUbpCuMEs
Hr9gnwJ0PjZZupEJg14eSum2noEBrzeaV5CbIXp+htQboZhmyW0TfllPXtPcQcvA
uVx5Wkbxibl+kDVM4AFVWIiUh/vaoHfcYJ5w0TDWebf6k04UCVBOVcLemoYRDsaT
lu/t+MVpNDgdEGhuNV4z7OihTuz088d12gd8/j9ZRB5jzUxCiiOA7WMaizVjcMVk
mOUDdWhNV9aPKlxvIBs3bv5/lnW7JXhzaY3MstCXRDtWnfrkbVYDCfqOgsq/Y5i/
vTwCvlNAuuEClLTAWUCM6T3AGprWPeWK42j/tX/GIsL4o5STZdPnSKfT5XPfAlJc
2wZ1UlANpR95r4GafLameAUmQISFX1snKLrFY3SmSOWFR1ehJX14b8xGs4X3owjA
U6ORbR8VFYHJqX7vcni9S283uTeIkgebRKNg4TXOGWco/oHW/jzGE/eHBt8i+Ri5
6G16+95Ns5TKT7bSEMgvWIbLPStTmS1MOBswLony6DDODsVfcQuG6k0aio7IPzx0
5B9ymutkWWgXaoYDagCe4hw7jqaEvfRWWKyX+NSxzsZsOvrhDwlWamKOaizWHb2o
4I1W3PtgW8TKhXx2qXuRqAwvjBu4o04oS7s5gbmpqEQoWFTPJNT5WsVPL+ifpRJo
LmuRcXd+INkvcitEXlENW6AG32OU+RqrCZ/7OeDDd07sIWPf1kWdI63WbER40dul
d6X4feb2zk3kvj7sviUbtEqhtyLCw4M9SM74JtYMzpyO+I/uFz7tMfP8Bew3gdv/
CALgAeARl6yYjG0F2qab+LmaCEumpx4ZfE99AdoFaPMZioFl8ZYSuNnbI7+yhXv8
u6rohrBe1QBwxWAYFyLCceiFkOADpJvdIVCT2cnxYpJ2nMAelxtgRYVpaCDxe0aW
XgRHLdgBI511b6ptrf3mlzkcc4P7Dito9J5WUZOjyFUenkhQz6te6M7jLNPLPPSA
pdR+RZhxuxCE2dZX4na7eaDvuuvjZ40Uit2dFHWjAnjLMoZ+Ts2lFRQNKhC5BTZE
d/UQxPPhQfJTk0YvLxXMaMoBsHou6Z/xuBMLoB7DFSt0KDkYjlgp7lpD2vScnyv5
SYM1MmtcrmukgL8SAnuHKwVbfU3ZNm9F6h9nL7t2ELKlkSjeH7JfXNwFGXOe5S3i
LfdDUUDzn+rnANdxKMIfkjAjpweTBjGyaTOcs6GCFr+4h8a6b6rd8DCNyHuxHGyo
AXxWH0HX8DdGOyr9F4e3I5YTxm0IBG5tjVxzylSpzBe0rrek7Yv8dkIlfgKT0dJG
ta6ZZ1QhrHfT0BREkrKD0dE+Io+ev42nTUqCsBmcg5bVMrp0TxfcDmkx3ScUpCi4
MadGVbQS/OLE0495GPQg0tDkeFKt1pA/xfA0mXiUnaQkqU/DNbMuMir12vqdWLfh
gCTIBEdJz1D+CZJ8zgFif06Z1Ws69Tr50uRbMpSnlKm+bcUv4tTjMywflcO0aWkn
0zQlAMVO0CFDOU4oDaeujXdYp11wHlr5TeqZlHfRWhvsX3902t3G1jn6qdkh3MFP
KCr12XNwkN4gUYScqjFlivv0cIpguL/bt9GfNvBze6eidwOzQ67D5UQBH2ccBeys
3l+EWa9ZbTMTAf/Rc4RIS3BWKLCRCYAyocmmBqD34OtwPe4dh7hgAc9o1yMkftBR
DvHl6W5FcxAm5S35Ij6bUeXnIGLdKMvPHY6GXHHG7AJ7p33a1Cjnh5l4Fnftc6Sw
XtgfrtfDDSkcx4FJn74iyYKHX7IoGEUhYUGVtpa5NF1RRHV+HF8IE2OWI98l3xSD
LiE1upiEy87T0AL9zyC78y1jIh/lMBlvcQvuJWkN9EID7lHk7mMKV/PuiRl6jlCY
pCLbYvS+go4Zvl2lS4H3NkzWubiE3WHkhiWETgFcdWzyhBDtHsyKWYCbsZT1LwRR
P/IVGmDmcJ8HMHMEBzMfT7gqzU0vuQon773x04J/t59GUqhufYzGoVtUo3QNe6Nl
bVBm/YNL4BbK9QPrxQToKI5rAE0l5RySRQmOj6l4eSDEWFf/zz7+9v6MdINJr3Wl
jIOfCShFtGv0rRtGc6P4vyaOfXM+sIn2uliH8qeXrhUSktQCB2oOVxxc7czJsiMJ
p8m4GsO/8S80/Py01rBjN8PfCy57oQzPHgXWhprZfMGzxAnCEe4Mt3q4Gt3u8GVC
veAQNl5lPBB6HtCdawulpoCHub2853nY+N4MVytbNiI07kCY2EvAJP+6PBlaTARE
w4sJlxf82HYhQe/p4AAnoCqI8F6O0hOaUqqFUsL6RzgtdfZMsLcRJT6YaaTSAy1A
noWR8ubMSifamSFGi7AeB3ze8992M9wkXkL1Lmx9ciCdf1uTqfEzoHD9qJTal4fy
Jwj753cgHQlf3T+eu5+BpYwpzMmG35Vy/Tdf8gGGMAMX5Nwij1z04E+4pXmays4S
CtakQPOaQQMloI7h/JsY40J2YQNqFzLS9HVy5XY02L9gd470aVitcqEP7HTk2aXR
RkmrKPKZcA+B9p7/2fQEMB337q2GZdufi6Y52x0FMzcVVlcgnaXTYhSg3VywT5yd
OH3bpEvGuSCepoFDQ2K0j/oKfd3uvHODPg9phdlJyyu13U+lzijASNqXk5K2NlzK
KvVgG/xdJ7CS5Z6I9WyjsqTfhQQ98Tt5bpAQhjtCG3E2Me/qDZGAvNbmmwNxVgKU
1byplbDy38GtzGA4kR4F5zzlFcT/uQt2HbtMIEek+3PTq33oqIucqLp3ai2NGHlG
sJXrK22q74BgcjRFn9wFfKJD/jqi7973gJhlDyYkmI7b4A3PsHvNPpDkKEUYeeS5
o3q/dsk6C+prEFx9sHYvQ1kVQErc8LlxiMFgWctVONhZI5QiT1XQ0PAE9hh/rGUc
dRjJPvCyH+LQDx9rRaXX/7QlEVECWCXtErhM02XFbw+p0/aOwC9CXy7TJXXNcu8k
vCqHhiB5FUWjnTXN9xZmUeiFbFw24jEqCjLhwTH/5oJc533DMNs9KGodxiu5zX+x
FwJJof4BP/VZQbeV21a14RV1nd3m8X7T5RerTpVAnM+mFkZVPipVH1tNcDK6n2yr
dbT7cf6RNcYSq7EnMKM7zldyomT0K2/o6DtAWq3GkxGbuT9/yWnGwRBMhUecydcH
zMn7fhYVvuLzusktCDKK6Cw18svvo2WH9D+TY3a4fBteqDu0UEsNzubVkj8i7TX4
r0pqTX9v2vgZb5GRvbKqfbgyqRGkPoFF8AEpThvympQy8fOW1qqzSYA1g8qNIKYA
ZF3pdilFnHjL/HlXKLgsD2EcQl6pUMVfpMDd5EoGfKs/D9+PIvbjMKVLINaUOFqY
Ep8sb55tj+/LTldMB3A8ef2yVlRNGRQVPmzp/SVGws4c1qYy0B7uOQ2w2P1hVPAX
75ea4bKhfAwACwdW4DAxzmGWFX6EtiEJkIIaHPA7NjuvTJuFFvs9UwiaxEfamL80
DzCk65c8B62taDd7e1Rap6s0GZuwxKHfV6OoM3CKJfFigR2dGwQGNfqmc7pAX5cw
A794PvkhcNXasXyPAeyUTc/zj97SnlyWxEqhVmQ90hwjfvuG2IbjktT9p5sqq4cN
SrmoZJeBvsklQe3qD7DUU2pRRo3SMKlenYgCm4Myl55X7cOYjdX25/tqyT1gjtYc
ReFT9tEqXBxO9JPsJgpAQErwxbKxuhmvn1Nzffd9cX05pK30rkjizN00LYk5ohRX
2kpKVCVdSK8A/boNYqfZ4uKvSaX8L71Twu8CS0FKaSr6uJV0HHPIDhrulMvu8hJV
1smJ5Vp2QV+Kad/sB3vzPPaNKWE/9PTevRIexcpkm2V+ReuExM57TSwKYmpbjdh5
G4arI1AgdlgGfmVJe12exhb2s2okiLnfzBbFyddvswyy9KqA4yS2ZH7pWvxrFWsh
NJG3l4J8XQZE+b7Ge9xUyGobVSj89DVwbZ7JHIXQyoSfHyWBi73zU/OD01WC9C8m
1cjUT0C+1wBoLo0cIoTq0si/8X2hSXQwYvtrmNJ2Sfc6SXC0NYqxmZaAnfUvDlFq
cRZFCBbfXmrC0mGz/4pbImT1Mp5Siop2TbYM/h38Rvz5wxBpwtnM6YCtDvYINKzj
x9zP/OW+TKBblEZUZc8KueZ8sFPG2MNrfbIdKAxvYGSPnlPdwrV3IP3FksAHv5/H
bZBBKrIQfm9egIo41XuHCoy3yz2+vrCg0yMnxaJ0dsFCpUGdnJjmZrdWUgXLajmN
URldMAh380oM4Vbq62a+ga0K0+hTFyzJRARMy+Ur1H3rBmroo7o+ulcBODehTktj
Qcenl8E/A2erv5pZUHhPKRKJFCQuTkwsn6oJrJxbzgmxexrTZk3kYItqVfNupK8X
H4z/U+/lImWCyDalHaqPTODVaOKTsQjS8MGzW9MQ228/ME96y4lNgl/sbEFEr5cv
P1kUahPUbvR8NXkYQeuOXC09SNII2r4ZNMenXKRWHoV+8DJeRWF6on23ZYzn+uO0
FO1jnPX4QfGIbmttMYEMTqp/xdBUqroFu4QI0GTK/Yj9ZzqZJH+GhvpbzZDVF1DR
PxvPfw+OadsaJ2EEKa12UepNc8LpN1X15CGtvXJqfYaZ6rNn1sdMJAL5k1rqKs36
fFIJ9mYQ1yU9XnCtOluYmn3QFCaw+iLvfNy1zUrRM/TBHyiy8PqPmYLWH9QCoSew
qrILmqGnjZKHjD2g5ZId2j+QsSjdzppPR7m9OnQ7PvdP94sLbyr8yJgOPl41Qn1Y
O8Mbpi68h1Q2GpaSkcW9QIjNnNtucN852PYKegE1yudijk6ufiKr3caqGiQreInU
jkWMiKsNRINDAKxhf0E6fc63JIGdnYPzAybfeeEYsolTfWfmChKtE8tUV8jOLS/x
Z6TTriWrDw7GtNWbyeIp5Tli2WSUmhyFeAlrKcavMrtp7GQ011hbCBO1XKRrAvgy
iSDyx5F2Cgn7tzvQMIT98jqSmsFKKpFEE69wXjMuMB8Kgvw/JAMODAFA5kLuVEGB
6AjuQnhCy3X7sLZKX2JCR+fwY4u4cI5QhsnC/Xvj3QwAkAmwSqnxH0ZBTFU11LYV
WZ99fSbyqZ5Ou7pY/NVhd2CNHDjW0BRt4GSrOoD1NSnR5uTPTz3m0Pg5/zB/JIGk
Wmnx/n7hWWv8mVAvUmkt6MXq5rDOrrAKSRq8Fv/ffV81vzWalGy4KlPYFYHKp7DC
3s20su6tTdD8AFfq/Le8tT81v5cqfBWX8HAvy4f3wweCCJmoninqylzR4lfa40S9
j5RolZx/03lFw7nt+JtZ93j6kpADhv8ydVx5hMPkZUwA1RLdq6hN195mkLrsxEb9
IJ3x5TFdClnTzjenW9rmAhArmc/4HXSX0ftrYVuiSe5WpR2ZEeJX/GDY7qH/lpR8
JLogkn02S2XPqHPr6qutlCzh4M7S39KHJD4EXBYtV1hbvP7yytCQTDPZL9VR04Ra
5PZXSC8jEHjHmAMPrUPF7ELldNF7D6Bing25XzReKu0ts/fr2WcODSkuvuNjZOZ3
dxPRgZojcih9NKlFWn8XONR7eWYwZHenjsEyd9KY87SCe4Ze+bEstgn7SDZpgnaG
yomL7mNyQrXn5CEVSH5SZ9WZm2Jnq8SUKXAjBb5FsppZ081H81R1J1XlM/HlT9ym
zonvSpJ/jVnZ5TyYBfWluJuCRxfDWBoZlY8ZVuquP17W5yJzGDcySrkel7mR5559
ncAL8m7b0ZZa/S/hrVDVWOd6QMSKaI1jr/TZofx5PAbmq9NNMca4DxpqEv/E2i9T
Phk4DxhoRaQqhWOQDDDjo5x9LAA2IZdQBLOQrVolI/zae9zg0MuIMG0malkwl4PQ
uVC3uyBpuaq5wvFyHYIyBH9rzz2G1CwIlX1GbK2SDL/P5QgWllAO7p/IFrwgDpZV
UI+WLGBJgL23EFMHyXgY/48W3lHSAcOd57sykKmsv4wnC7Id07Vg/V+AdaJfTCGa
41VFuNPZKdQ4lAvGnhzMV2m0Ob6hLyQdNT0zTA0wlmXSXiIKWUrgxiZ2eis3iGju
aBlu19do7dw2FErkRZDdFmfF5cTAwKfJSyb72OBTM2xD5ChMTuc2T3Hj0dLBHyb3
ta3C1CYgcnZmYjxvN8bsW1XhqMsMLU0n60JKtZZTv8E/bLYzK8ZG/ZhzTBJId3mR
OR3vU2lxKvKKMlskbTDol+4ocjewVcHU/nb+PLAWtk8wYkds/ytJfxZ9g1lggh3u
gdzvnNbHksLxaeSBE2cJnTSnzbnvEyVsdVSjFmKJpxb506TJeesKbZaOxlCdivyl
xzS3H9sYGrzL2F+f7x9Y3haHHln4XklvWwQhDnm5iNl5WZiZ5F3QhSZSKkv+z0HG
mFKKybow8iV22kEMNAOL+MqvbzhE77rFgniOWVNy6sjBWGM9mvkhhC14YbvUg63g
YdpweuOO5Lbkln0hHdUub7DdoVtsYGOGBqdHu33ScAtfH4nLzDoZpvY/N4b9qXOg
m2GG1Eo+NepXMQC4u+PRl7jBiVcog31a6eQl/4hN4ajqibe3uLgdp/zw7GGU0AdJ
H0JXt9H6yaTO7lp7X/ozG5x8zIt8e/RleyZgL+XOqm+OYNXHTY6dNZRUp66AwVsV
bjalc4ils3LUZvtj8es89u8Nxg6kVwn2hTJJ+K7RmWnCBVnV8SceGkxITD2mckVN
dh6ZKQFuApN9x7IYvb0Ch83eS61Sb75cIRao1feqpTzhI/0rYQLVGnwQOIzP8WRq
TvYtaS1rXFcAqmLEGApPTtfva9GR3lUgzj0SAYxPqqpEvS9BzZTUfwZGZQgIsbEL
2x5ZluRBn8f+Q8ta2scKUmSO7ZQ90MJKcmITHNgBxa3dkMRWGJ1ArUwQicFehgl4
BMVMeyCT+okFoX+Sf+MBgO2Dpa8v7he9wzmEKz7mRnYfx2Y8Ym4HbbYjjzoX9tij
G8ctvEN+5PkSR3mDvsr+5HZF4ZL2Y9oFxK3KqoV6EAuOpovWPgEOdMR5Ks7qGaZ6
Nk0Nr92WYyXDuSFK38kJuTxeeDMDj5Q1ifpudO8SIj5lxkCAXGLwzA4UnZ+AVpMz
gwzMHwPB+06VtdCMve00TcGg4yhWtEeFg7sv8PAnOUYz4VyrzrHhO/G5vDkGcFLE
l6HG35rqFkAmS5UG8BoleNTscBaqvtw462XJ+LiefnvYBMbSNwxsQMjc6LuIhUoI
CtVinpLLfVMhun4Rm/QT3yvSp10EZQ5r0zMuRZACnnERAiJOi0ygvIhm5g0x7FTs
3ByBa6rwGeqiw4Ahsk9YKp5iEhIieSzfkBfAcDhFutJGS1WHBbqnTjCj0JbH3x8/
nWULtwWEYNmTChdZFXSlKwyTo4pefCIwHd2fh6mPg2BBO3zm1HnztqK4oWEV5l+l
sVm3RgKNvsiE2Sca3lr8BHlHNVKsgyHRakC+qbHfnWXIfTp0pQBlDL9gPR/qo8nd
tDanKpOXUf8gy+ybVoMQvpBLy47pJKItFj6DjypPKZYlOr4TA7yQxtwtpzpHrAOz
ouZ08CS2K4HFOKX4oK8Y2G1s0gzzUJvSntTj8zcglmSla+6rdS3n79ln3cbPN9EK
aKx4GnVOIN+rmsAGSJfL4zms8V26sRKDirmVdAzwL7CU0LOQTYWZzuKlh13a2dZQ
JXHYsnRR0ZH6r3OnCocT10jDUpuJDCo2VPKuQR1BKFytJV4we+a5cy6u9aNU4QHL
MFKqAoZ1YbX6I/HnM/Ndo4wuIXzhck6q+V4pXxnmlsJWTaeLrslY707jG111ICCY
mlC7CJ+kIzzu5cynE7cB1ZwXo0FBohBqTtGg+0W8Nvx9y+K5qLuIxh6dBRUyfdPL
3ZZ63r2khOu5hZbZFaHRscSdE3i5cv/j7XpRba/NHJovO8KNgmNtzyDccnthE3Uy
hyNbhTmCaO+ffhpOrD2f6I28jUyb4g0ChBKDtsUBZGOT3isZGZi8AR2xfeaRkVYi
wPoOOP546okoqiHZOsGb/25QSX7cWeYNsuL0vHplrWyIPTcJdqDePeZ7KKjRaJ14
SC8ilVTv8J6GFd+HDdxvkMIcKeTI7M5jSAVNA9McvdlCR+zxnvE0tPWLNhnoncYx
2wQCHhP0XYnKKF6umN7VyRoxk5OLo9hDzjP+s1mLYnRq6i3u/4EyhcVDF7zl6m1a
7GKpDHLplpQhpNhabWA4lfrlZi3JP07UV3Fgr1wQbw6I7yHRjdbTiINpJlNFBFKz
iGocBFbci6XoBc3veooePcSqchBn5xQFKUSftClShSfm5Iic9OL2VFQFti+gotQb
zwJU5VNSGy0tKEvgnKEshkJSIg6XEYKNMNHY2rKZm8ZMz0AGO6+96MQ3cyn4WUVn
nJNlCXon+h6f5wBNBwr2q6cuMLE5WcytIiIKe2lUWS+3CMeP/hxXvUWkDyRltR6G
tpu3KV8hoI3YifA1AdzVOyuZuRCSeBfjxY7TvqZoYIt/oltX+CPbb0iiTZWby4WU
j3A+mAevtuASnyoO1mAWf0rwdzlzYZgMvpkMJnBvKM90gLAHokTcQtAl5XGRnZtX
3YIaoas5Zm1Eo69Dmcl9dCiFTT8QymxruMTlT8/hpT8hQPZWhTGAaVsS0LQ2cYoX
tDuWD4AsJ1blw6fM3rvFF94OZgx27wI5NR5exQZ8thURinHP9PEopp4qbt7imqxo
Z3Xr9rTGuLcM0DXS8CMn9r9d+QPMZ2qey1I/I5Yq6lEFPVPn3Lxu5Ig1fPvh87Td
kIKN0Akg6uIRAGl/ZrbiMw+AWVJKA+INuj0stJddtsuLDDMUFQfq5mhuAYDEcsze
EH6IeS+edYtTXlVIipZuTWfPwwpAZ89Q20+P0bQNxR0LtSq7iR2wCS0v4IEIT/C/
B5gshguFRNsXYNYBGMq7aYD5nOaIS2dBUwR5oI6Zkq47CefAXaWohYIeIDjDc4iV
l7srXo5pBnjjVPu7wmyNwfYlnWFSer/fRrbBZayTvL7IzA/J5y2bQ4brQllulFDS
gnBZ7mYtlgJ+RkoMp3Kd2ULzsNaa2c5TXyFM1AiLXDbT6jolnlRcmoTAt1BSD7fe
hfvWLSHdugTkKnYRQCeKG26ikIXbRsGIS5prLeiMpsXBJ5rHkHkrAIzQxV+1dGaN
BordST58J5rC9iYzZcigkhLLHKUTLOElScFI0IcbTihrt+L3o6AOAiRkju30Zf3I
w+evzVmM+j0jAqKBX0Z6dCGeQwB73zNyenOqJXhFaXTTid9Q6i5GL+7R0nFCQUGw
AoRiqxUQfC+oOb+V9Cd+qi+WNtzytavDOJdEgy5bbBU4bAsZhSOAMVW8EKRpCCBk
oYYlY1kSHK/CBTKeC0uSMjblqYM4q991/pc+NBNt9hjVKLy5U7aYkuOB+cQF+E3P
PvPUTjp4fQarPcG6U9xqqWW2ziwy2ENuGyIJmyf7pLNPiaNtyE6j3EzoqwO7+qoB
6u5EVB7MSsZdyiHEb5Iv1FfT4DA1yDQyE7bmvsxgDtfocTpro2zLeW5pfUSLZ7hZ
k2oJNxHYtNWBxG/aSrOsh9r87dv3UeHmlEeAao7wqFN8h52Kumj6r/tDXqKvm9zs
9GyFZ+6obKYO7QE3zsZ+2K/sJbpk6heO+Y+M3tqjn9BoNWrtoMxLMmb6phpXjLy3
DAxeOLwn25DVdGqGp4wRnaXaveH3KcoDeD5QTNXcOUQjDEv0s4/p6/1pBSJlyevJ
pwiXSR/sU/4Mv1aCGFwtmxRUHoE8Ex098pRzCHnSGOzz+S54J2KXHLFQx/c6wNue
NcLl+4tfmGtqvrfamk3c0AzbgkzO0s0kvziQ026gY+qUy/4a/LBKbnjNfEBNTwgD
DtZbE3pIHfn68luKi2QmGAt+Tez6blb0uZtD60JKtPQYiuQVEMzx9+7dGBMzLCD1
TrWpdn9pojq1pOGR5cD9gNkYExq7Q0lYTEZw0tX5xizidaKsTniudiJxJO7LxLgG
Ec8k05DCKDisxQKCakNhRFMWyr93jIkuBfV2/3GVztj4u/xNqTSNLjva49TtFQar
u8Ob8JXDQ/011ESKzWJVhekN3Q2KBkKbOaFIyVljZsjYKKIIbCXFe74AkR8dyyw3
t7dEI3pwi6BlmHYVBqgt31jeDMv67bzmMj+V/YGAC6OfBy5F8nbJ38JlP4ExUKsb
ksJrzFyq/tTWjRGC9pgeXqOD2ygYcz6gsjgG1RbiYzXCETR4+8NH+Sp37sR7O03L
GFCGcAh13Q5Wpfz877nicfyMQmwIXXxT19macw3/eSxN4i+JonupFoZjLtBAv9yq
DdlpAegymgybDxbVlZBGBHA7u9lWxKn/0n73oRCJQK33EQpMQ1BoF4AJJ+nIGkvf
9SZlYPZOPegHbr9FROcQB9AZm2k7ZsSOXKTCORlVh87+ZP3MOcyzt98K63/531Vm
uMH9KP83TTliLF7vto3cTJZiBAwDJG57J/V4QUL02Lqwk+gaoSfKcQTh9ZiehSXL
V+esfBoW4O+AjlO0GFXHYfRDM83c+kCzcufdr8aGUsY9TdI4Wi8ea6c8NY3Rnpw8
SpaDSSeH1zebtE+/8RVnFsFcDRrgnTXUipddUs4p2D6qgcHIkUUOeOqyOlFBvvPh
BV4hETD2v9ocs8UC9Mg6Tcqk3HT488aSX5bD3dWSSPlELSWL8VGkNVYlonJpOsrw
VyVnBFc0aFyifUxT87o+DDBxmCHhqzW31P9J/36vTqBx0xUTqnvNaKqVA+aXEXPO
Fz7sJcvIQr8vNlFIhgpuSHynke1mnGo/HlhXcTNMHlDiOJ40DrDVMznC7Fn5Qrpd
O/EBvDHQpjj3QY3RUY6PG0PHewYT2eTakEwkQbHhYbg/agTD4K/KGPwtFhfiSoRL
R5Vp6SUkmXaiLcihiN539TzDBrcTW2z4Le9Jv3pT43nLzcaB7mVPVNGJU3CVYQYS
Zp+kXSvlRECaUklcwYQIPX6ZxO0TPLwOeV1mLya1ed2+tDMOAs0/YtK4D2V5w/X/
niP0KAmal7EBLStBAef8p1vaItY9fVoHolpLKbhz9kufo4rNFzQov8/d1Sml8GJN
r8yuqwGDsshkZ+EQ6TQk7lz5ZOcmZD04yM91aszdXtgo34GW6MuFZaLoxe4OIqjM
aGgBE+nHYEzbE9sOpsNmsKnP1EUC3KR74edFmKoNBnizh9ea1kWayKnnfnuARVsp
zsRjqjJRo6tnbka0yK0eugmFFUrQs7y8V4AwiTp6unLPHw+KXrSFEzGceue5RWQn
N7jQgzql9ZBg9LLMrjE8GTt58fU07ZlQnnRLFrbd3x1HV6ubRAyFMSt4S4eaeHmG
vum1sOWQbvm2TWRz+c8ZkfQEwfUVS1ScD9tpnPF8fXXJR3m5E8Iacx7S8WqIQLHZ
xRfZH4Tst1TsJV1swWMbUdoJl/JCtNdyVnmtF31rpNZ5aRac1t2PZuO/fxwobOf0
0OtwAsQ4IgihAY9gkoxq5Ai8jEb53Cm+tdJYfZdDtl9mn/zhqokfAqt8X8H0P2uO
yW/au/82gd4u34omIidrE7npTu1Njx8B91gApPIcC46eMoGJTst95DFl8EY0WkuA
icyh3E+g9BKNVyYj0cFk2uOFTZi7Lf0uJdAnjOpHXRN60hfkAzavpCMG8H7PeOQY
8kyUN8gIkBCXUQPKirEZPt5T1+bCWW2Ux51gCYrzhyrFWQq5cNtPfYlH889BtY17
jgtgAnx7z8heZe0yA3ObQCHIFvkIAUR44Jhrt/1YLdf3OMp2sh9SRuylLcgmNu4K
2S8y4vqDMNGUpqBeVkC0b7BpVtOaNNGBgaP2KiNoDJw/F64f+xc85Ur16cnM8HSy
cANKeU/gOqWUjS+ShJL+ouGpp2EzrOuDAqE8A0EgYMAIHEALJRirD4llDlGqlv+m
EImeJ+ml532KzJNzzjxciouEFQHMFDOsj+x1dPeOfFWtCGX1YOhLZY4I5mifHt8q
fG6mLIdE6NgThrqH9SwFWn6huGHNX6pgsyMY0EFYboTN1h1msEhLpAZ4RzMhdpQj
OyN5BLOzBx0qhkHEPECVnZiHjNxgN9qE2zgtI1yoO9JAJ/+QKHIAhCSIeyKjMnlZ
aPmQPC0Y9Wmx+jTqEJ/5QjkoFOsnygXAUts3V5RIqvCJhhrEkSRaUW73x9LE9WwM
fP5OFjZh9fEgY10i40Ms3/Fwmrs/CA47LioSdelnN3d+YlOPkWGqAXp1tDRgdV0c
1I7J4qU8vS+Mn8vPaP+ng7kSeBSR6AukLGsAwtS9z3yYjHC659tw+PyaNnjVvu/R
CST3I5v33CQj9Ohn0Ont45dFIuIHX5o5p9lxHmb0Ljew54rUmQXgBHNlb7brJcSa
H524+yyyHioZ8LUGcaaj3TtrB7ZLpwJhYlpR1nBx+uTZ38RVMdOY/1LKSxZz37HQ
4RSVSa5wo3unCyeFtUAOw8Tr2w/iYqcQKHj6ShxfxuYZWpVICyHDXPPlP9Mm6Csl
mh4+aR+eXwE9+JBXwrJsnTVYJp+khpXvCErRVfqYUYpUH9YsqPiDQ3jqVwAxvOmW
rHF6NvrVVRMEDhdU4JOgySEr6I+nR5WuO2Pt1/CC4pshWHKqNI4l/71u8pzuZZR6
lVo/2i9vqNQPqgWFOCpblDtlo9D9srDJILA2/5lmpH2NXutn6UyziaRMiSJw5y+v
PQZKnBN5uI8V9xLHHZR1MPbyQXH5ihi7DRRXM1pDKqGk7UdMPlj2QEDB+CNQpRMS
/UAGBt+WDG+aLrqlvPjBA11fJZtYIho1jAkIgKi4NzAJvDGDTW265JOQ8TSPCYSD
gDDeU2Of28ZlHz7gIham1eb4ey6RxKSQOkH/fdhU6qn9t6RYHg1t1JPqqg5x+h2h
STtpnFQMtsFePZWJNgZ3Xdor4wrQlkua/K6wCuUmnFup2E1+qCFoAZRIPH891NN0
KYcHXByuESQWz2Vjn2Y/lGxxHFhBHMN6UmTiS9s9U6UiKGsCNxIcPLD3bQ3qyslC
V3KcKH5YQWNo15G2N/gUmqmo1NuhwPnmxn0ZSCV9HGpAIEHrHdWNk4yKViy2ogkb
Tt4jaOVdjvwZ7I2cwnH9lf6VNIwanXN4iJs6AxxAbkAvGtvFfGWF5Br8/RmgVNRc
Xu96AQ66Phq1MxOuuwwk/Vco0ab4LqjRif3N1g352x8EYHFQaCZyy3H/UgOh0FVr
ecMEfphvDaeq1fhdCsJmRt+FLJc+DCIUIb0FA3+ulw3QJgs/e1nXyb5OvC1Q/vuD
lBHUfyw7Fgza/P/fGOk4UafYYEJjZ4Y2vMfmPelf3IobLdaaGmvWTB3S0Sw/aDlc
2V5CvFSj6QOaEpEcaQeP/kqnciMvyj5dGTdg3R6XfV2Qf2WLXXCKhBk7tiPdwmfT
jJBasueOVid9oulOcnkOXTNQw0vmMrE2wNGYFqs3wRUNFLSNLe3NB9UdlREkBXEA
OXiSL9+q24Fq1Epvz0ayGuIl8dxrz4TgcmB847bSMR3gUM5ASZEO8Lj2PqpPryXL
X5RappHeNIBsrltVmKeu7FeP2zR1YQuZrO9sT8uDSTMVTx+p0e7U20FbhNV3DJEZ
+S6LSfpNKUezXjAu+N7+Ba4Y9eB9Dc5LY2onh5aCrx0iHNlCiT9dFyNS65R2XZvs
GAEzMRIQk7aGhp0yDL5FxCZ4+3Wd/l2laV/dGBUxLPNNZUSlr2DzY3GIZHJVuOa9
NZicMTk4Qy8bR22tooDFmsgEygUAIaWvV/8b6cxwDON1QcCjhpcfRPZmWAWOHayc
lQVFUCoTr0o77Au/dTVTH1dWrHnJFX+OCd2JGFjFdbKjNHs41i1QK+kE1fXfvenA
xyFU4CFbEcHbJTHwUL4s5gCHFi7dZFdlDZBQspGXnipuBSVvIpPAFeYmRtRwvITG
oG8qu50CyrLdtMKGc/1fypVMVIgtUfywIv4toX7hLed5IPjB/sXXBdfiQbsJRsvl
stEBSiuxfpJ2vxzTo37J794P7OEr8PSDJmlcaAGSuyJrjSk5HDN2YdaH+yFgidv0
Y6PrwkrZ2npWeCt1YgCdJJ/9NX5EQ1F761mCBNCYfABQg4BTaB/Pi9SzC2gUmNgs
P1SPPYjfYYRiThZdnHpjkEJWznLkZIt5lvb+eWcSXPVFy413qa5Fpe+4tF8YrlUj
6hnY+5C+uxFm4xvJ3mkE50grgQLy0SMiQX4kDR9bVexKeJ7PGd01xgAlg582yHPX
KktpdSy0Gfm/mkoEyAsLQbi/l8nryS8IG0DRJjpS9iH53IJWoOSPZDSfISq7LSXi
ItfwC220935at+Cjpy2W8Q9sA1fRna3flhFEO+cBTy5VBYzr2CG5qanN3C0DSOgu
FkrWPeQ2K0BrLc5710PKGfr7TT7Wl/srSYXVcJcLqnORWJmUmEvkExAq9rz4ASIu
QsEMgQcyoU+borsWMHxywsWlEQ3s/IvKqMasYdeTZOdiPuFtgab6YtC9SxMO8dVV
erPTsmRh6GNEQktlG0VDT8aOZu5pggPY0nwvPTKF/cTapQvtDM24vmW0GSfREMmd
TUvleqDcO6NAgkNG5CtZoWUI+t4A1gpIEFC6NajfLKNi7qyZU+HDSqMAvjrAcevG
w7fquQJXy6Vpx1WkH315CAed6S6+TIyire22aObHlY9hnkjQZ/8HjxaznQj2iPwn
HFuwKLMysouhoaAwQwj4VdTaC8afEtr0cRtqSK+gVR0PbOjRw7nHSJCrQNX/nwoT
X2ammqwbvAq90LuSFufuk8hJeH0nxU0Yxjni7Oo8kUqD9RqdsiN+Ir4Xv2lYHf5f
RD2TnSPqzutUYPswiGsaevpf68xx/07Fi+gHk2kwVN6ItWGnRQvuDqAGMQTkmxyD
9gniLmBa4Xuut7q8TxcoQnx8Y0cnQugwJVvQytON84xHHkEa9ISniKqyQzEuWBZ1
VWbeaTNAoIETTGoXk99xHW+T/oF1wsJuImgLt1llarmojEnVi+7wNOgYmXbwZfZ5
ss1gCJu/HvUMOEc5gfF4VoxJZ8VmrA6+34896nm1jAlAN9YOfyVfR80NRnhIWfNw
ln5iRAt9W3sOV8bcUP/sa3ews0RgIXPdDuSGdHauEgtNwClRClxuJFsJ7pPtEaXz
K2s1T3di7KkTQ+mPpUAViLuZJ4PzYDClzRrJ4DPf2b/drY72cU73wW7JM9wI55cH
EgzLGq2+KK/zLb9l0pMnFEVlCQlXMtLObc0YZPm1u1uNZswDL8ZbMQL2D1FcLqJw
AVvN2kUaa9iPwwN7xMABtFWP7paRSh7Ot2qv3uzH3Pz6xcgLy9N3gJPsi2kCkDS7
9bhxJEcL1BYrHWlKIjryDZC9sqV9zxAfmq2v/DpweAU0SVnkw3KQVVovDhcGHQgZ
GVOEB/YJ8NOCAdC74RNm+cKKnkM5YVvcbn17Dj+DLf3ZgUhDLCP1RGTKHwbAL0l/
n5AHKQSZaHv8unPvo2a10nSrDpKvBTuTFXX+kBFvLPxhqEnEKa+BEgSd0a8kLUIs
qAQsrCBdiI9lyW+3yd9cD++l6OuMuHi4dN3huF9gZVaEqEcYC4TSfSV84wBk8DCJ
7NTZgNT+k6SAP7SB/Ji39Bp2j5Nzz7PFVKniuiFzuQ+uqjaloztByF76gmVWY0T9
K90DsEqmYdbYZ0JV3fiOl8DEfJfLfpMdwj3AqelXrZW2rNVPxR6I0NXjT0vX0AxF
0W1hPLvjePRjunr+Ecyh4xaKLHMZGpY/RvkSnxjoggXwlI5jCKbSU5Fqq+8wefEs
yeOG2/oRLAn4YQbDFmv2/SYmP+ejy8qjDMxXJH4zSmo4kdOnhB03cARzqbvW6uUP
KZ/mQuG+lg+jsig4H9+onHLg6g5qY/lPh62sba8ToCl3dlzcH46Ogvsx8ZAtvVRD
k1fOPkIIFT7rS09MGUqvoGZsg545YuglA+Lt48fUpiUUhT7DZuYAnqhgnIrlKS6W
6MZbi/fpEgia2wRMNDp8yJqkrgTCkNxq5ZNs9upqf8AlgWfNXNdFE8ERBUZh3PPi
4lGwW4wK3WAczLEoykYTEp81bo/6xPSxEQagODy5fffSVMSUshIcYLAoAz23oh7R
pCR/4jLb9dfSVXakcGlrETZi/32DDZ35UE6GCZw2IuKAi501f92211yirJyi8h/e
XKrX5eJk+beMYCg9yH/X7p1O5c8FsFB4KJwUbXDRCpor8nY/IJoOjo4vYy9crsUY
fp+NkcEOAi6eRBN+ZwCMI8Hyv/UJi6ti+t7XzMuIVKkf0WcrtlaKna5pGVDN9hbD
6NPzGgZlbN5oHXFTN1GlcnsJ3FLLppwzjTmGRwSWcYcnzquoRKGFypaS57KgaB/r
sTqmrj0g1qI/oSEH3rb8fg1tIo6bov7B76yuw1OxCX+G1fGwOLP/gYyuAOkx7NlU
hD8lLhjb8T+TffeFwR8tuvkrgQD5kW48qTRLWlAMEQRQU4z+puc6eE3DoToa+pX8
rwnY8hUYG/v5lCrP6NRIbr4zcdPQKUifM7NAeKhdWtt63jGgvsjgkh8JueAFQXJm
JGXHeZLBPZGBZdk8QlKtIhmp1kof5haewsnV8ey7o7/c+3k9923cja25eEUGk1Cv
k9/fjgKu32562PHRA1FzRKn/Sz4iIvqS/LkbYKvFSgNqhVfwuhxvMw8KATi5hEtG
qewVchdu5hkCWsyKouqkKLeb3h8N/35X33cAx/oLSZSlaxZDAu12W6ZpoXco2iCm
tkY7Me79yQnFAkVJ1wgxhAvu0kYWxdfw4ssSaNoU73TRQo70OY/vYDaqPzbcQ7Nm
ONF7dT1dSK0PKPnx94jVzLnPQfJgIYQvoi1tWfYyQ/7nGVtDrWusV+PPyeLqUE5y
9zHl4H7r9TEPzYNamvYEa7qa/MxeVLY7w6SV1rPZgMBCh42FHiqkvOJExSgkr5Jh
azLd/THTAZ4aJ4RjgTzqiFCVXp0LDt8vrnEPNqs1idHxCq1yXU2zoj6hkXVRfAdt
MajHVDrWzhd4I7lMSiTMZuWliuqfKw8FTsYPWkc/IpYxwLpAgzCbSE5c3fXQQIf3
U2OkHsluzkKhrvjfN5yRpO58GTg2QVipggV+nry+66mIddazT9vHkR6vpLkSVLaU
dXe2SgGJ6YkJ9MVEyFSDMxoLjyzaVjAuV9ECymgW68e8eRiMFkZmlChYzF53jaMB
bS508YMi5AHe6v+Boxp/CpCmpZKU9SVfDenE6fH2UCNuTRS8n0hhF5iZLq7rD/7F
iDTAnDmbe2Tx0YQsE6k0X8ij8SnnlCzIsxz+Znb8EOTOWg6ngzKVRtxvikIESNtF
5lo+oGyVzU+2W+/E0lS0ru9IsAhN5Qf4qUs+WYJ5Hz9Q8dSlN3DVLYWhhVD/41ln
ZJ4tCu8y8z+AjthdW6PYwVjPvrNeC/IQM6Q2dwBxVx8pFRdoluDR2jARXZZVqiz0
RBFZrU1AGd8lAWm8J5CE50S9G1hreyT91doCd0jIL4RHB+oi+srK3lLQ8K759v76
uEI3dMUukweBzWve1dz5kNovJKP7kV+/DYGVWrxcdGFsh6alqp3aR9NZW0xnLwgv
2u1S7X4fMnH3JXUAfwFqE71BhNXWz3RaxJCnKVtJYqcITMGIBoMZuE4r792qgHyD
ZBVAFfV0SqojUvB2LPnw9e9bCOfQMid3/tIctF5fXnlr+gKh3g9LHupSOZ5APrAf
3H6/cicnkZ0Xdz5D1cmVbmVK6+TOlXEs/+OTlxBcsgGP2T/kYlX+Udsj/URmLXQo
PRUhYPoaU4KO7GUUBCFS9S6SiGtArKWMb2YICaWVw1WDwKxXsks/QCJ+J5+ingZP
CcNFz7yPhuuDzxY0DGa5ax9Kt1VSVH7XpuCIR5EdzVBzMJA2ziWRviX5bsOtYvlH
Ka8MPk0jLDASN4w2QUAcxNqilG2mOwTpdL7UjwNV6c2QgIfMv7yqPHNZi4PTBkpk
/+aDrmYMFbdnWresEwVbpa4Mmzom3iIGyrBR+ydoiCOZWkcoR6d++D4+tnhV88bF
BW5ZNK9/X4wG+aQNhZsS19otzL75LNe0H9L3LBtKsu1Itq4AdeDOdWk98pVEi52h
0xdsUxmyoNtCMKUr2yZeC/uKFkaAavu23hWpPKy9sttkzAJ6xWJRxY4eWE4xH1/w
iE0/lOIczTiiymQ2foXa5fpcH1yPeUQdLuIhgFJ0K/ENrNcOLOe97ZJixCe16Esf
LYkn4I450mQ32eclS7qM9z0zNTHS0cqJ6A13vTX3VgGGgbmdpXuKM87sLX8NZgE1
kbC0sdH1rTbSvIsOZhsCSeXsJMk8yIkbdKbFVubTaTirATiH+uE1Xj5i9Zeal5lS
ioBF/ZsKz3QZacBOdqnSG49X9ARE6DMImwgHozy6UkywjelSVTMmTe8RTtqL9P7n
H/pwj1OUT0kjFgAYXXQJPn/cZSJlXmMwwakIbOBlvVqfiZlQ0238lOJinkkFzlyP
ug8UeLphntIUXZXjCCnCy1zeqsl1N18dzkPpYg5ju8VJAMkIqbb6uQisYVu2aqag
ROvzJ1v5TOeyT/Zij+F4aReAHONQfuwr20sXrZztbcSc2BJUm1NCFohGTU7RWCYP
wB7zflbSsv40581XIuragt+r5RysYGjnXpNnznYmXR73cjJmRjudNmrJaJPac9Tq
uuaI1j6Z8wdaQl1eDfp+UipZt32ab2hxsInkoCQHXV3jNoHfenGlVz6yV9Z/c9yY
9DCHx7DJQHWPimaRCNNiyArXxvX+UHX/zsiIYtbKwGhOPzrmJkT2FZ9qXHVw5KD7
M+K9AZlHHtio7BtuxVpINv8zMWJa1hw+QUll1YsYVt3Ho9UN18LvHisJbGU0Vf2z
1jm9Eb4y1+zfJpp4CWTGRnXgGaTW9nSk5Z8o8lU3i+A7picEg5tfrB3NRAInOaAa
QmCiMXiw3xvXtdAXDkwwMqqbo3RlQLoKuRjaSehhl+tDOiaR6CZiwbUJItr4x/Zz
QEZ1hEEavDy2OhooQ8EKzYxJ3TKsEndWDODWVlMnA+BhoWWpE4ZxMY4KzuqNqs08
b/o7lE7PiEvVdzCpjvrRMx6a6I1AkTqv0nq1t+oyAR3dBWLN1MED2177GrCOAZI/
3uQrRI0qaoKkfJBid9veMx22KZLrYfexaWH0zDLhopywdQp61S8paGokJND06RHr
8CiyjgNjiBzZwgu7fjaim20OtQGdAHAIuv0+asz2ynb/vsj5IHdI/F6TPkx5O3Nf
cQuk/jt1gtITcrd3ygGwA5SHj5JVlRpqDYQBJ7b2fq75Lzqi+aT859NUngULIsHE
o5zF3zE4nPNJybGF/RzNf4/mQ59RMI6nc/UT9+Dala/iLOQHfA7mduB+GkYkRPKm
2TVdh8Ay422U1ejtk11RS32PM8xZDQA+UkCq3lAUSp6E3oOPixraQreck9dvhlNH
vQNakwqLaRYGz8wHhzNMtH2awJQSv2JQL9BFEZKuDU3CTlYpbJ/S9/kgCo66z2zt
RN/M8nbzhro6F9s4Yn1S+jZ6v5oAV76gHBwV1r8+N6y4ReHWyDzWq+F96v0V6vrt
WP5ITgGZ7SVxdIC7w+PNlIQe8OtrapF1WrHGOJJI1AwuGX3/DPdCllUdOjre/QlZ
CDBZPVtx5f0lszaQUJ1ZxT9lvCb0oAU6CoBahSJuOGXzC+pajZ7/sZX+sLmtX6BS
Edxl61C3Jeh8sbb+rp5iBLcwaF/01BFFXH+EeWSpLPks9LLht/upMKWy8fuyofYG
d0V/P+wsk1Vi69+bcvDHKlwgIqAKbbzbdZg9dVliBVQv76KUYdbgUXJedGfdbtpg
JQum9v6TzJz7qCzIgbmbtSm6a/X/gQdE9elJ4wBTZ65e32azZMI9CMlUjp2StFmC
1b8eQ4yC5GC4Qcxyw32cgmDKHXKHwDd45PkXhHKgSvrE8FaDJmhZvIGoz760j3tv
LmOVPOsBmuvdONr0HfZ+7mMBQrpwHJcTbRqmlsccPrYBZvff+Wa/evt5UofA0IH7
+TGuh9UfxaNJ2l7FcOkicku8U0dfrCHUWAQ5ntd3AFW3/3HjL49a+fdn+/b0QzAV
x1kFhhQ4YD8MQ8UKEP6+Sd0IyC6+816wXDnjlflEHAuDDXSzvos6Henz2d9kMz0r
SypzJe9Kl+rKtfAXogEADZ4veTkLn1wVtUhelauv7wMi03s3vnbZ0bwSf2ydOW5Z
BvSFjMo60Vc2ZGtUtlYqcLLoEoQ5u0bahqJqrE2MWGEDuRPrzNKdVtTe1IFhyIwz
xoArGAT9W/3iy70lmqyMexjFF3RMWkLT1NTEDqbUGBiD1Qw5blFTkvuYRH3PB/eC
rnoFwfpM5gvCNM/9vyoRiTPGtKVZ1Eot1NOcFQOUgFvr1+eQGXXisiup3/c0Kf7/
3WdiU1k2wWvOAw0WTudAAPQnzWtjQt440WWunI+4TDnIz0a30UuVLQBwwEUgMZGZ
zlziEEZGlztYmz4wEPFwAbsOJk2qRyNTuRpNvFanW9rfThIaeNQs/qUO4yhgLyuG
8GeQLp1hQdxCa3cnBbHg8rc3xEAxJaIiUT02zyMJPAKyQIZnhXYMwBvvHgu25rI9
FKpU7JoydyCzSYDupR7lwyF8jyPtAVlwzYNAz/HKJQ6VLv2ewyWSlEfqI6MG9r+/
CX6Rt8OmRGW6SpVCecBlVlZv+BY8r7WyP3StM+/Ml5A41Cbxu/9cc8T7GArYTBxZ
8CPd0bHbcc2n5BXbIDlhsn5y6mun2eKtlISbtugRWrjfwmtzIIwDMd0nQ5Fi+ZMM
ZO9WagazMLziN8mv1dQwXsCaYQgO3jib2qEC1xzVwOT+/ZVFLHmKD9Qi+0sj45Zp
MhfkUeDe8cOYhdswBec5k4P+KWfU8eexvQl6l2zvLT+M7Z5v1x3eSOMNkiT1qmgR
jQg8eopaZOSTkuzzrltfJX7skna37utanV11wTz30Xo9Hoh9lFWzQ2kY1KI5BkW7
NWPlClvy3nYP4dznnET/h3QLHRI0Tozj0mLRR9LX+8qTIB5ld/VTuUEQu2ppH6h0
rGCNcI+mXgz8ZLLzsm7Rm5jwvvr68no/eCShxZzoMF67PZT56iveiqQy2ak9hX+E
NX2iFP4KSPpVZhibnI0PxPmIeZHus7z6oI3TPe/bb15icUgov9cizh502e534zX7
5lrvNaAKR4BnDLXdPmjuezbaYDfVPkB6NgMpuHAchu2XMszrUezAS75Jvbqwvkno
ymXC4yjKq48EzaEwW/FeDa/rb0c8RMorBOHNfe9wWr3dsdtrjyNHWF0or8PggUD4
L9yECjY/RUTuvN2C16BxhlKvFuhCRcQR/GWozXvBkkms4jUsuZ+gFAt4+Hcb2Sz/
UG2oFeG0R3TWpZnymmFlhIg08y+FUjOnvkybPp8ysCc7TMvL5mfc1AXt5reGWkf7
tTHRn/SqE27NAuJn3Blahz6WG7qpjd1dCiD4QuDa3mipvlt6zzu6OS7UFzigqK90
xHyTTYBsSOuApMJr9AHFsRwKS9M940/T5hbzUwX2ecBqx804qXBuSW3c3lT04Cab
mSLjQqzjun33NgPdAKEaFa48YEY366JABUv4B/AvkeDrCttw+1TQGryCg34V6CdV
rk3DvVLw7NjV7DDFlUU2U+vgrU/9iZNkdvLuLTj6hQiboTMc+mynOKdgNOjTPtlA
JDR6lsEc/fB2YzdLKsgNrTtCcE6IpmYEj8D9VifhaQLYzSMkd2DcPlEnO1vw0lQu
xukmxNsMKlvmi4ZfievqAH+aFusq1sylCp39pmq8MqzEczJ+EsYQ2xco+JzNnwQy
XhpC14Ld+ZISJHqYNfmFh9KDGUY5h+KkeVsQw8DhadelcFqptwKfPiLiVrVznxEK
a4uKlXeISIu9Z0s1V9lJpi2iVttcKSf/6XD9xtdV3qUF851b2KP/k4ypP00tFJk2
fhHY+PU+ZSMQA/9I+XdPVZhTROJuDW4ZXVPkA+xfbAojesxWwq+ToXcnaGlbOCMM
4oF57l6KgkaZvdIXStVZUDYhrQxSBgeJkPe4HfrvMNJxGLzRWlVda1ejr+NGOB+H
ccwhAVfFZhw7cODnAs/WX9CZdS8xBKpfFaOKIcauO8FR3eCoUQlH4KWkGmIw4C7Z
J1LPPImSsO2IO5y5PZGqvcyCQ9BKt8k4J1Gds9bhemD7WX6PIbBaLPJygMvgYYBn
n0suXKy3xmFIHGwkQ9bZ4IQHNaGV9dY+HA2bvDVEb8MxVAnJkn6ckXUrCtgRMcyB
F2imhGwyYUlgoQpwAPmfQ0V4drAQle9OOc8AYFfFWStZqJn26pQOHvh1E/YalVt3
yu5tfeTRdqxickPfgHZORbz6vGFWkPNSxcG2Zu0EPdfs0hoCXQPDOcdl5JkjlIFJ
rG0cgQ0xiE8VbAis+chIhMQBdgwgUBLiE3hfDwd45475bqCGRHm2NwxI/0BQf+tA
0QHCgeuQ/+5iaJRFyzGiENL362KUJlblIsK24Tbms6pLI8ZXW0QjTsKsKt1u/taA
Aazgk6G6Mj7HyTlZpSe+XvcfVvZTFwAbt9ozZU0ZnnjGBFkUHDd5S/jsdReaSPZg
B3hmsd9uYEUGaCSwvwBHjbhzHm/znV3+ipKNq1mumG0nlBX9mKzjF3T3aACOzllA
jWMLwi6N1qGMraiqOW3JvPcyNLpmJVXbdR5VE8UgqvAoPN26/kO5ptnVPOYcMQM9
fwNROKzTFtS3n1YM6W4SE+hLsKC7sM/rvGz2fMvjMtBskoDDF3Ck7T8UAgZJMSH2
AJ7nFP/G2YWqBqYTpkAN3pSGT6AyajL33827pvXEyiNwJ/et2kZPoprzPvsGSxsf
Jw67zqoGAMO237UlLjt1e7K8dKeadRKzotZopIiAa1clVUPIJKqUS+Plz6rvBOo9
CI5is/xCEH4ZL8fhf1AQjtZbowbaIRpIqtWZSHhgTrm21+q39A25g+MpgUq+gtUN
1QKrm08t2Riglz67TiPRl1z4WuqfbydmxtBqGgKndOw7tqB3cjGqpwqG5jIsI+qo
Q0pAO/ooFr9uiP+bk25d96PhTGU/hn91iAFnU01E1f0tEyj+amXiJnIr9+y7yBz9
NrH6xu1uhpcaMxHF4TizYPkvrBTeofB+jAcH96RJHBu/lRoUxUZRg+Wzt+7czZeO
tmeyxBRk6+61dCPmOd8wgzadkrnAzYGxl8eqmds7nAwr3dVsS9wwa6SKiHBIa5S1
7Dwb0vh3tLZc1QpMKz6EQO7WkfPKlahFMeYutsmZEMIm5hd8wobjr4P/KqA2vb4h
pg8aiXkVPvOzfmP3+Bitf2L6vj+sV59rqf7lub1Y1dqjWa9uVUEwp2OxYU5OFQzx
4BcbO9aIJ4syWNu6hX1WMO8AY8m9xSFFXJZ0z+CzDs+gPSlJ8nC0XHdez/gBWzSs
Rq88IPV8mkS00560K2XcWNNmCtXo0MF5FzUPhUh0NtIxJmfyWLCEcZNjude3B9fA
gdgwJIXJRWK3l/pIcI3/OjnAYXX3g3Hk4nQPplRVUlmbID6uRhlrl357g1AU/sBa
x/nRHgUGwlLUM78qnv1tINkfiMKCnq2R67yMh2ymdxvDk8JIp9reJBBOJ8zqaxTc
/U6Zc8o2Q5MR8HSPtbJj617RfkkJbipgj8YByFNpTCcv4roXypFU0bnEns4VJxK6
uQGB3sukEMnXmEMXvwBSKFxXBDw1ljhtYlF2eZmwqdZuVHSuAs61+zz7vyoMLghw
b1wB262yNVfjrdMusL102KwnzRqsJiPgSlwHbnT9DVr7V2YhZcT11pyDusaLLu7A
Xv8MhpYLhKDkcXhl55RQBgEX7m3uVOkqID1ougjU84GMbg4C8XVe3/sq8dz8liD1
K3nuudQdqBB3lg8C50RdiMeC+OxxipOqVA8i4VGUlFS1aJOdMre0S3vG33Ry2i2I
qfpOhx4bU/dJpXJ+MEGGu9Wuz9vASyj/I0w/4Zp16nRnjTzrkMN9+dYYXtMc6dSt
ypUlajDfMT3ruVjRPhiItq44zFBEA46HF8+PjR4fEKeh9RS0B8N+Nsk9XUnJb483
fsOUXeE5NEzUxNWW3mqTINfh1rJP8sth1ZLQla9ARDqE6w+Y4j/z9GrtLQoBHfgK
GOi+7G+jybLlcGUDuFD+HFgWhSl51XSpS40/gwT8prptACj8aLYOoMTIVqIBVsma
/bfLU/p8+W9QfoNRktAdAi4crnbycC+S5yrVEnGrZ933o1ZTNY0lydhBbZZTNNuS
t2q39iLKpYDLF7qWerVSdh4izaZo11jboDARcqqFxXKPkQeBXWaNA8VMvvNcdPH4
/1woLvjzxz2dnOs7+NHfOJis7bzYZfY1wJ8V9Q6+TgqkNw3zyk8P+HlW/xsAVnYd
ZymoFvJfZdMhZq0Sjw9kyeh54JBN57LI4RSpv5DtS4VTb4EtsEJxeUxEhPBgbrG0
j/YYXo9JJF4M65gDewo7RXqvyZW3sdPYLK4BlV1EdyviJOCFlYCao/+f35lHmj1M
2GvTTZnN3QjiKDEGVV9rFEkMDCG5Q/AR8/u0P7hSwSM962EALH48G7dtu/n2CbTT
y5DT6Ik+Og8CYLa9aRcpyJsheGO6BCVPbdllojg/avIGWcSFHCoDyqcUDkSPrSPN
MwWIqvkUZCeW/S9TLioQI2gPdWsUKbHvJQDs1i7ZVh69FOJ57OhVb+zhz9FvCCig
C2vg1UU/lTwUEFBpVr3UIuuhJIdsnm6nSrxOTqeJnswVPGOW/rgbz6VdUgDXhKQc
lWK9Dvbxq+4NHDYEqQjgWQhRnT5WWGqfiLuitNt+vGBcgGSiSuxRUPhwwM6xmCer
U88hMtEZxvxAy92zIP21asy7c/+HnJojC2l81WtjuN+Z9L79yRa4DAKkHdecCXH1
9fjklMxzSfi7t+ns+RBs9+Lb0b0jh8mDSufvXc00/yhgdIzRS9vpJ3uYN4nLSmoP
XU4Udl0Y1bkwhnKrH4LKeS59zc8aU9xDOHgsR0wpq9Y1q159ALGILuJCan68g/oG
7lBjBAflVzPm0eE30KToew76wUS0I7vb4k2zfptHc0Ujz2yXtaqAKt1f8kDGLJW3
pZUFtvYniAnsxgFN9fifAvQTe5/4sMBc1rZ/CY8/qKBxVCvq+sYjMYg8yoZ8t5E3
eggWJyXL2vdhGGM55Kp3LpYpLlGGhJ5jX8TKakjSxOGCSk0zRaqU5RSnD633DzIE
Pn1sFl9PA2QUo5Cc7mnYAEQH8Sf7JK5BBdPAAV4rlE8v6ewCqEfyTA49KG+V8BDA
6BU1Bxnl4hrkl2x0j1nKyD7BWB+MtxDpACMZBMXmvk8kw/cppCiaHxchC+fm6Hpp
n5BZuad55QHi0ANpAxL7Y6fPTN9zMUPRc5YMjQsS/k2weWH9kM37Cd2bVPRM8wlE
rurm1AY975j+GmXjRUho0amrT8/tPZj4vQJaHLUoVpMeK/feeov/8upZZtXHY15x
U7E245cNFTLXGRP6boKmmlVKhFeLHEIjtD74IYvkBgWOsMpKcZmXl/3BCKF74Xot
hW4Xx3QTvzulsB6WtN3QzMIoexObc+Cne6+SqFgL8rVF6EqAYnbDJb4TkKRyG9KB
P5v3QbU8JsuW2ZNC7vPWDQRWuqGc1aFcrVGOWj2mjacRpZgbFM4Gc9K4EwesLJon
a+Dye+8il7qKULvnjVRHxulxRGMpKo0Cz7o3sDezuulMaxwjuU+NMTNq6L2SVQN2
6+EmkYEVRIwGLefNeuJ1CG04vESV8DZZiOeuVMVNat3+1UvUe6fsLYHO9IP7CG2S
dcFbi5qROhw7wUuUIyimKKoqqVzM3vCVzLDJGgQhVaII3Gsh5D6SZc+KBcyV0qRV
68FtRLoaw76qTeQUztxeRCTS4GRFVP1nJTvLdbdT2puLyfM//q7SBo/rgeN7hETY
VRTq/4BHCyeeSdom6kNRLouAuiq0V83VxfZ/keo361nrVZ8+R7kgho9K9LXUgHwn
C4w9S/pDSqyyWuskcz0TqV2ZpDC8uM9Fog3tULREIHaomqENrfodvqD5RQEkWBkD
4569SQplY8qnluWe1jmZLsbx3cxJwB6rxXXx4fN2B+mHneGpIdgB7TX+sPXdXz/l
YU3GVqnZ1xQ7uMdBoygBnp2RA5VpRQBclIugV0P+BMoNNpObtxwUSfgnkBzWqu9E
NqMXduqveKGMjnQ5x/v5yMRikM83ce2jgCFkndsLbvKiLVQI/WmItfr7AdHY7dG/
48d0vI7wVtGykOPc3TAJg/YammXgcwZmEojT7jaienMDtSrP4ocoFm/dXr6ZGuNx
7ouygBEjzy73qCmJ3g6zTBqGZNngqe5Kg7n1rWxGOvCNStOk+0Api/Z8VfWu2/mD
+QtjGAj1oY46rFrtWp39AGOxm+zLPW0ZEEn+u3CqCAdz3egUzmVj6HdVK8j5Cz+X
lj4sKfQN3cqtAYf/ZwJPusR4yK3+smrHEe9GgKAGKPPBKqcfF8h4KT+RnKc8qgzB
QxCRH8OZ9UPkPUhUr6OLSWNRqZ/LnSWhX2PdvRX65OB85l/+ZX41CFEv0gFEKMzA
EohQv3iTEDBvppky4nWmROJxBeyIW3rhMqI5AXXYNUnSPFNXWq1868S4rHyJCrMj
vgp2Y2V3aJvkBUACbQchGO+NZTNvd/kHngtbZayCaGHOYnL1OL9z4ZV2NsVUIxCJ
JRatVupuXxtQY0XRb82FKGFD5KYTxWysScWq/QiZYTkMKm6lytoIPf6RRFHOVl33
WOg0cDbgkIZbVFe20rpcgEMn9z3RgQSNXeipSvIRib9klP9YTLsGBzF53QQvJFiE
RBKfbTLvEcggSGsRaWvVX8r/CzKGDR672cuUPVWHiuImEvaEiIztdtOlq7c8Swyl
a7o9OI8ZMSbxCKv62gjpJJ92xPR85b3K5dlfJfdjHiYiK3MBV/joZq5+2AF/sXEB
GWYuLpjVN+mAFcsgD2PyZRdXMLRLHKl9EfHf+eBxqnn1WRg6xY3v5bhqr0Y/UvTJ
M+xjULtZNW+e9xxEGEI1G8uSS+QvR7q9Iby1gCgl8d2piY4Q04JsT2wR+gqctiKi
DKKSa10/1ztv6NX44GR+sdTT7WcuMmdP5P2I3H5D50jaHD6DvUASHdvQyy6PcXXG
P4GdAAAmfhs644jP/BEEDh/wm65vXVpsyJjAozkZ8XdZUYf65wnhxaGgwZgrd0EX
c1tLUvXflc/kVIkkBNUs1xtVN1R14G+hjCJbWBybqmxAwBTqwhbpDl6hIPFpT0Cd
dDwXKfgPPFTDQpH9KkHBe93lx9DL/OdhQMoPZYjoiC+Ci+w5qLEqf2wP7UGLHMZw
PzjJwqrgZEhKHfC9hZ1syy+qdQ+nhjALLWjwBIBB/wIm254IpXb2+rbJVxTZm/xw
O1tDuvulrg3a9I4PQK/CFxN+VNeug9013tfhBI3uSA90VLoMofklCMeAmvCyrWMm
t3yGgKYlk7VnWrxO9LIrCq3OXHgBasWwpfJERpT0+H9kIUQSsMdzx0eT+6+TUAdE
eZcSzphedEDkV4bX90kCk2N+4ACl5BJ6puwGVP2CFdHe1PB+o3rbYv/npoI/x+6q
PEy8Zl0CmU/aG/79Q1M1+30OBHi8vJcmAekeTPw5EUvqL/CjXkaY3JAUdKll6iev
1CqsL5a7fgyJEHphvGeJs50dQQEIdcdaZlXPQZTrExXIJOiXySzEu87EEccDPGWr
uljgKsxFSeH1K5issjYw5WKievVpdNuA6wDZB3fev7weSV02siSue80THIRUlgKD
zfsI1mB0bZXY25iOdkkGljjtM/S0iKMtmj2OVfTGw7qP+7ZtWAr/mkzTx7IcKQb9
mFF77pT0EqXxwebUbXfEphm80f7IYS36kEP541wdpjmnq1cm8ETh/H9f9ZTf3d9k
N2+rXKuhwSHPK7vxyLZJ8/UktsAl9zrUCkpSwHM3bhUaBtLUoW+QAHvCfyuzPYUS
5itWcYZEyFX2qFlT79n63QJ2YPGKoHQj/ub7etXmQUoX5tmcJwaPdWUkcdqJ1G4G
Sz3hyncJxKB9lDmiAYvRshRm38BJf3RKRD3U8wwM+ca3G88lRHAT1D7A7lxUnxOW
ZcgEGuSzOwGyeX7y0t+tuBZPeUS/vnBGD9whXHEsg81ZC2Xzf++j5tQgs9s0ssPG
JFM4+OWex3TiwnTo/3ergMeZc6XG+aD6FHDkxOb+B0FzM+wrLpOTqQMWJjNT9Vsz
JtdocvQYl680DSlTv3LIPgN0mSctOvfogZswbUwttnv7lGkBMY+zJ8HElv31FX+s
faUwHSZZuXa21ehN0V1Dq6iZvI3Qqv1A8/Yo1wNpA1/0oHwUWyPkvNDRhhDu7utE
KkOFyBLtuZk+GAuUgyysgVTsfrkunH5rC4uwq/2zUEuF+DXmXLbVK3FEYPNDqJrM
jvxTVLxiRXwgSevDaAokyhm7weX5E3HtIduBPFIJTfgm71/H9nFgoXMdvYSU2WUE
5JVc8BWSEQuO8ahddvi7/akTRP7gnRdAlM2tM+B86MqLwhAK8ILll5XcXWxi9L6K
fL7racNHwtY0YI74DTxKc5eAJb4Aa9URWIvowiQVLt4AdEcD4rnMwoVmLqz1TUOs
NKmaX6DLT3rOlAXSd7wjmQwxAopqKHvTbiSk4Dgo338MZFMA5O3ZJZXkpmPMwD1N
d2l/MYh45e3DC4S/TLXoW/TfZPlqsZdswANB+3ZsX/hME1VMiA/R3elPttygQzNv
gobHC57Mzx+SyaSY0JaIiMfME30rC6jX1VW3xcRNWY3CLi7t6mxAofiRrkNW+CVG
VJRBKf/7XFf5G27zQWMKWQIfCoSkwIIr0dFSuVD9/tWzEuOZjkOTCXJOq1DSbYmH
Re+iRXMppMrO0M/cD6j4/FXinKRypA4/GN7jisg+iII7geESOSE5IR6zUMX4fq1x
+mC7f5JUeLj0RLDOdq9sLu4VWqBlWkmzLgvVJj91Y+JRza/7+88D9yv7alGaxbsR
+1+0G/I8ie7OVzLa7B1vdBHP3SrT7P+cxFc1oQCKx0+HdX34ZXYQSEvmpfjmduDi
eD8qM1uyqW7CjaqR/35DOUaZJ3Qdt5ayheD10WDYWuJwUnSwgEpCyL5jq2141Qcx
j6k/jcMzzb/lQ5pwdJVSpCyDELv8k0MkQLk3mw8S1EBUioTQbqb/NIO1d9HxMKff
yo5N6ZXirOG0r5ejvUb9Ctl2zxJddVwzxVMhvMlowk8CeIdLndgrcmSSqZqYY0Wl
WvqZuLAJRAqrxMRar1Dy4Sh2O6CVvojjYY+5O10l14qnaj7lNvGa7Q9X2ZTahfOI
754TObN2jQ5wZmajEDTLBSI9Vb0eFbV+uiuDyeBSM38zuQ0MdD1VrBksvLyC0RgK
sDd+niGm7YuHFBicovfEMxGkXExofvLCtedzfqoTXb0z0PUv7MuH4d9iAFLxPsBc
priaZD2gzp8WaBycsEQrBR+QaKkaQJ7xT30uPOEAmxDfkKEZeUTwBJrFgbVVIxBr
ZhMWHh5NHvot5Os58cLgoeXISCdegFI77xHckyznRpsP5MYdbbq7ZS3QNBqOZHER
J2R3guX5StwQyxmN7iqqa0CpTnF9UgEQDzcN/UK9H9IxiyV7sfQNoriIwb0ZxSuo
fMtiOC1uyhj8w3Gj4nZxw8Vw9EBd7MIvC8n3ILSSRZatvpKX2e9MT+rugsDbrovS
+eHofcMWiOGgDUiLKOKLFkpqvPxdwofnsEJZPxMwMzJHjq6umlAOq1bRYRlKY67u
dGT5uvlAHmNe2XDDxwMV6fEssbVWHiwPJzQiOj0KubrzsCFL+utquZvLhGlvDU9T
A5/QPeSt4bI3oLhPnc+Bhol40aMA+MjYn7HvtLzluovtCcbTaw1k31iB7jEA9rT2
frGu+kpLxzKMTweRguaOusdPpt7STDk6FBG5elF9FIrdw1Fm2DLBTQwik71HHdWd
p30zj7xVxlNYSuMbZd8tj6WYHlwzEXGIcRn3L5tTLnRITKcgEsAu4nN5GTfFutQA
dW+SZeex3U0dVLxQHyWK5eAQjduku76GaWjBt2+3r0d8MjpbCj0P9T3sZv9BqWVN
GpRylDsNFhTpTru6iTmS/o5LRDKyqsVQW0BhT6QboiOt5EYvFVvDN0sTmiW4ksw5
8ZAAzpw84ci5oJk73naxDxDrrnTWKerHYHtWKwwOYWBPyQ3s4ORcSLxX7zrOg8CN
sAUARbxBrcEa+fAnGU1HvPH4vN1HuwERB+zBRzZsumz5wSNoFvjQV9A/YVNj0FFu
T9nETaiFqu/vMqW8OyczQl01/sBWTvuoxN/KGFQi613oWlUK5qKJLHtHGC2FB7my
EUw6kjl2swII/dHIb7s4lYaPCLomuWg65RGyTiQ8xiA/g5WGBnc60pMhbPr8b2Df
zA7mmWZ5LsFCXIT9edZeQv0kqNoG+XmAWxl4L/N7twoPMquVyHi8wyaqJGpp/OU4
zPQpm+tEUggACSA9KxueQui5v8eBqPIeg2xl1KO6kYZTyWoAg9TKXdDkn3dZcvv+
cHQVT/eHh1FWaq8+GgrUPhBEBmfzhvpv+WhCjr1qu7/SShmf9QQU0hHN4X4Hc0e5
tC+tBDkWFRysMywbZjh96ZUx67rCbUVTxZbTDdYKUwpGMtvbmkjrXVjskeEZRnnu
pnBgNA/G1anNf/f42j3Chc+LuFGpPtMJpR1rUhbREKYFTGQsMZNb/sx4xZJUxT52
giahMk+wtuTgEY8h8nk4YHgvI4gRM0gkrtr3V/rvB/n+11V9lWB+l9F1D6MAsdzT
8ll3y1EK6KuKnJt0XG4P6xg6637NBXzS0hdv5o59KwWfct7YMQh3+cdsVXjDdakM
oY+e5N7cONWxwg4NfN8qeUwG9+IHNpHlcr4EteXe3JSBeAQYnsJ197qhDJsETpi+
tl4ZY495XssTjwHT8pAqej8z82MsTnNofWCQsGdE3+PaXm6sZPy1L6kBUVJly+WE
oA/cb2r7KafJ998PMkX7kHhTlMCKvzne/rypYLIXSvZX4udm3yq+7d+P8rrVfol3
2jqq20y70/Uiuc5JnzOiKd0RW8H70wWfugYnN+jhmo75HDC96bEGRJNrzblaTTDy
kz1NRhxtoKTk4fqPqlUPdAj5kWYhotOT8n6Hq7z/gkeW6Ps2hKBZVhTAi/oDWXHe
IyMdOiYN7X+INdzfx5o+MjEilzQP9OKol21AErZ06Gy8+mvGqsmm21NU5tdSbAZr
x5rseUkGd/1zA9ySi9IpX59tOSFEyshsyLZ7hsWn2KjpA+QWcW7VOLZUL1pCFKNl
uRes5S169IgKrIr5DAzF6fHFbLDiK2+8XZ22bLWEuLA8FWWN5ZBcwHRNwl/h6xzq
QjDc8Uc8wr6az6d9oJf1CBzTyfzn37beCeAnyeOMr+gHN7OeOE65LDQ1FdOSDKVG
jWSGt8XCY3fFTNp1iOGogzrGpDtW9nrin+LpGMyNKvUC756WGhCsi+6XQm1N8XAU
goZZfwG9Ayp9yi67JJXvGmutHcMVZi6AfOrh1DKjf9UbrXoelbE9JJsMxRfcliYY
X9ovKQZpLQ98ruDuiFKZVRBQR4gK1M/qFNEmO4nf2zDG70w0Z24GpnbdFFjxqwVa
eXQXRR0w2+nduTb2O1YQiJwy4pD0W/MBUQvKMShC9xP34pV6Q9pkVVf/Z4fjzxOZ
PJ3aGuwMsQoB5/1PL5q4xh56WeN4pNzq39SCOepdBBjbS3O7hnIY7CF0H/RWpAFR
oA07g8+XY2ByuXHF36QLQEI1RjlGLsYg5OGS0UwgSaOhRj5I8m2CG4K3v8EYmsFM
ndpCmk9QEBXAiyv+Myfh7DzueYxF7l7UL8W/P4rwlZzGEeIFhOx+WCSp0VJNKSy0
I9R/As+GpYGkqVjN4/WoGrXASxYNLIsR+AY9wq7/Sk98mbAN/geTHRdYc457w/Kl
/nuSjtbcANZzaSjqcMQ7C1EKrWiFIgZFMMra+YcYy+fVRe4megz0jjUsZhpJ8we1
P7/Ur3cotByeTXBgUt6TV0mvfItrD7UWk9+YYnqqymQKYKgjZpnXLSGIyB44O+Gv
rotdve3jKwia1nPmisAJItop6jhbnWEEZeKSrbZPRoBDi3ihkz1yHTIKEjcFf1er
lM7Kw+huc1ODMR3pHFcy4D5THpz2/Z9BYO8ySgT9lyxOrDA8fhBlRH/1mrJNl3ie
z+9vjdD9+KCn0neWpAzMllwpgUbAXVr3R04o283TTkEWTyKZisJH3p4/vuX9C2A4
QnrRzmmmsohXthrEVBNzxGL2oD9FPIjyBjnvuzxqtehUMI9d4FVEZCTI2Ujw6MEE
QTjFvnwE0R8UqrqroAhIVKyWUJG4W2BwZlsmaPcdKMj7Z7AxhwETLyr3BzUAGcPs
UVYfuuoN4YgChwEDpnaecXtSbkI1C0DXw/5NYjw/HJzGEEoopAzU8soqm1xjXCWO
Mp7Q1bBjjaGzWi7RasoKysUDZZdEupjgpY9QG9nQ/wcvfMuBekFEDlY64y8FMvjn
lwOlbZFGX9PMd1r33wBL7bwcCU69W9OYXLBycjP30s0WSjWQQtucbJhnBuMtc84Y
Qg/3L6NqAflzddKVQGPxF/5YqjlIZVjDXKQ0bdOT70C/Eu86Ah3ZCOQgine5Qdk2
QO/gLcDhiAfcD7H38a9BCRvhZ/pYvzfe/8fyE/7xrYDUhBMjIILMPG2HX+LuMwUS
RQXSSn+dteSKq2OVG/XpnOqCNJahojlkeZzgkMbLFbfxGG55QgSNFFrymKbZUE+0
lnCth+62hndNR49Z7ZdDLJ3waU8YKp9sOatHbzUiq2xICKmAoANRFZ+3ESsa7aTS
iZNL8KNWc/Lf7vr27hTchqXwAzgH0EVtjFNKD6c4ZCDrT19qKHMcmANlR5A3vlzM
aq1zdFIGPIoVjRyL52Mc0hN/sJ35hYyrg184Ug/Y98kGnT0TGgsRE1gjzXeGoFv0
PFS4YHvxrJJq/UyV/I35xQO5ZoCPtz1ofzE4Dj4l9/aM40BB8xvZqwpBYE4kInUG
gk/X/8WGgBfDNAuMkkadbtBJRVwREglyTME6zjPagH4PQxkRm8d20w/3y4wJ9MI7
yvd4r7qa5HoEcdNkf8hABaXqBDjDEWF7lCsR9dNYzVQJqErbNstkgIFDDM1iR1L0
hhW83zIV5PGQq0ixmrP4seid3NP3xgDhMCah6Rg29aBuNrejD5nrfwq2Em0gc9P1
+1PLVPzZ6KheGP1Av7KU2bFKFSlv16l1nEbemOqM2pwVT6TiwUu6x8rB7AG5xl5P
pe5vy6JmElX1StkS6F39rYNo/pwNN8CgYQ5usqDC8gZhm4pVNC7Wg7Q+zJfCiDUA
M9C3rqKcRwTu2Djio/F7kNXlAIG7WLBZEySY8tlyEUwFwpFihC1axv+eH4KYM1BX
GtxpsIuLK/b+2DSz+bKOV7kEZdAqW9JteXoBVmdNuGBVFxNmXjmGllBxgechCX5Z
/XNmswL7wDRTfi9122y+BLJexLc1ebHKmPyzSWeM74eNtuo7Xshv/x7sTTZrU1lH
/DdpmYPP10UiL241HrzHd7iGtglmgX1hNWJY8gpeA4OpYqydcdBXWwSUbMOUmdCE
naRuyR5n17eS9VGADMtVm1knRwGyeRaGRvIRRLY4rfm+NlG/i1jo9QRJgMa2RvXB
q9MSIYIY4Xl19jHUzhUhRiSrhwELBpDK95GvO8RI7W2S+we/iKUfZbt01VHCp+Ue
myXWF5u5qpw3aH1Gg4C/Aq3aa/Abkk3oRMo38hvokj/TgmmqJe3e+OPpIat21nYD
LC75XgwuoyV8XgRTqyZnjnBrT2vxVxkIAaJAfNU9IWUt4JhREtvVvaoOdEDdeEjz
sHB7lkuoRv5TGnagNeCQxu9AhqokNNN8CthCEsmMlokJE1V/gi9nEan9iaHT/rQA
9ONleVMIRS1jCnB+w6fu3nmoZFG3a3I2sabHuA6r7Dd69Lbp7zOxKjUcnIEVyw0X
ldJLXrtCw6LgG9r9vG8BUuBLIoKz26jdoXn3ZoxrYblm8lquUEGj5lgslffpE6gy
Igc2hkTA7QpOBj5Kd3ed3maa/V78k/Cn4I3G5QLy6l3FLZ9hHfRk010CPZ4MyjGk
qz5bqlRRhSFu+gJywXB3oWjBPS7nmaKiyq/PuPWtAiMWqTdq2t2xi5V8XcUEMf1o
EWLczY+/Zch77/uouVwD4U/ZnpOSUABCvgnbtP6YMbfg0F7OOhdQpiZoWIFtTnXy
2heprWgYVf9cfl8gl7Jw6+ztOqX8gbAERptCiLNdlGcjN2JmMMwZVmk76ZYXjZex
6TK1dwqWclPM2tSy+hTW1bIA4SN7lh+QyrxlXB3DIyejLY9Mv+HDI7jbT6bHc0wY
bftLTPHWSc/wDXYuRCGqNlf0SVLGVP0bnVu0yxYMqevbXD2G7NMV5jwaDYwYWe3u
nomF012SAozyocXhd3uHZHtLS8EZL0ZBK4rwxCtL3V9i6nfPeioJUqI0ZDc6hRrF
Y0fmkSE5DNyfyU5DhWwFGdZIPbz42yYZVXa+DpxLXgjMddvcTx+8aMDrLW9mOKbZ
D0mfU2+vfKqGE9SaaY5QM42cVU+EqkrWhjtrPw247XRsI/PN3VJjESosy9YufNgH
wAf/7KneqvGIB8n7/pB9/PwXvP06W5+hEGRD2Snp77N/VBG+fHd16JsLDKS5Cgve
CegGsGVPqAxJN4vyGKRe1EIaN9m4o0vO5vFHa234VcyZGNNw5yiWxaK0Acf/dYm0
ldoAcb3hweJ1ojX3fepzUjIgSaMS2xzmpQLVlbT3Gi6abdTEzrj0A9ySMtLStPa9
AehRYD0ygurDg20sp8yCFoa/xDiCdvh4GfU4KNQ+IoKj9Z4ojSAqKzaYC+FAQtI3
ZWlIb2WrfOpQauZpDPX9wazoZTvniN1WJxBpHs2salNE32yJHsDuncgGIWET+Aj5
9Q++ooXIkbjmdjIp1O9NamHAOSAJroSQKCBy9VVR+jZFcYk8rw+rp9u5eskT19Vb
xVd0APyEZXmM6RRGb6SxMe4m+ll+A+sy8EcIzvf6h61nbzCLG5yY5C0XaIHHs+T8
p4Wyhort8eB+10wzxaZDeGwCwuw0gs1jkd/NyiCnhI7WjRgmUI6sEUoDdMVncMTd
oFXEMTz9DKOS9As062o6pFEXaKH0vSv5B0bJxQrC4LOyGvo8siWx/0XRWrBY1z5P
YzUnJBhpMH0WKDb867/FvCBAQWFbLSeg9hyOz+GqHxHVxa6W2e4ignn9JbM/Bfzp
7GqDFdNyPygaGr9c7H1nuM03SCUumgf/YZnPulTIBZykTjMK9iJ4aj9dFGelmjGs
09EMRozIfDkrTJGG2BC/SIE+QYxfx9pL71qku8BaJmi77rY2l0JvHYXlRqepZVMi
UfM0U/8wFgf7FO6qsSso3VP1M9dRkGR8S/mddvZOG2zeVe/p8TPab/bX0x7w/4W5
ldQ79oaNa3/STrsHM5oy1NjFWUAtrvQpXvg39A+pSh/Cr0+HolpgPJcexxZY5ZU7
8EUU4LgkdQeYOlsdbConMESwBMg4h7NTKH1jJM8fvR5YbxcYzta0RUZnL65LlrRm
jkfNERD2COEsSEP7EhV3eVIdM8WkqlVkh4q+f9aSLulhu0Y9FJlJalkDO2sN27AB
QdKsZEfwCEKMgRZOakNn4m03DPVQg2j/6zJ0vW+1Vu1j02Aua0JL8iSNUOmLEZc/
PTgWPjG6xJLGtn59iFFBRycrh/oLZGh8jhzCy+zU70Df9ZEKdYVdmU4h6WFEnIqs
gpzWEQRPL5dmPNHSl8Ycp4ndRPWpBOfTwkpHr8NYvb5wUvUBcfOE8aSaHWKA0s1V
lEEOCl5jcV8AOzu5YjaQbgXI+S69JThAffAmPovIkqX0ApFYkN744e7zGxI8+qq/
dq3fcjoEXdAXoWO8F8g0UZjX2AnqacLX7+y/C6TfbsaRb7XRejPogJ7254Me3RKY
kh8ieaSObLrduxt+APl5QyZCEBPog7w9HABN6lPRwVkV5WoKctqGj5he8hvm+SMT
l+/+PCIK6dEq811ARH3SWjzIi1UBB7lq07hn2L+V3jq96UY0KPWuVH7+WaerEchs
UqdXFh7Vhb1D5nZqm+K8fbjtaMC//CHJcZzS003QlhYMc2lJkKpqcf2F9N6JRjX9
en9GK+p7rbH6ogviM0gwvh43Ub3UyycoMcKktWMSsnqTkX5oa+BarS0YBlrEpLL+
ZaH9qMhywaW5Bt98tKLVaMl9RXcdz3n0o/jwxctDl9H6tsFsJvTNS6gJGzOKIPZ3
s/d4pAU92WG48JPNibeRMMoyUl3qNSYWoMa9+W5hySdOYSiwYBJKgjVHqDM81Gd+
25IrmEIHWrgHmumNS58BVc9FLVHKmOXKdUQmHTM7ykVOZ73UTd4OofIyNQYWJF7E
2uPH93MQSsC+reTPVsrddX8ZUSzdIk+P85cyuiBXJxEMmTQYYHWC4i3QplJJlzxt
QxygA9miDdm8bTkDVAQZoHX1B8rAryRKbOODT5SJsIIB1+/FTkQNj8GvvZZxvA5h
+AWSIuvuUk7uPtUbn2TFLGXy2kiCRP4MHPseQLxqZEQozWTzudxq+sPRtUmcs1X6
sfh/l2EFV4+kQ2iGnOpvs1JIGapRfZZ9E93qnFbQ3tVl6Q06yXH6TgOHh1xJ7r9S
8kBsH3I4ir5l2iLOgxyAUawQrSR160qbf5fUtxtcnuOUQk61WbpUI2L1RVZ6ZFXo
ezlikqh4VBhmECojj72b5cWtfjxFYlROusHaxB3TS7Od5xTKnad+DWk2+1KKJlZC
DrkvY1aTchxv9kgbDg5F16FMFnS68N2w8jtinzcX2PtDg7PSJcvMHx0m5Fit+2gk
w0fsOrf/j2vGS+sXgTQvFm38QkjxjKUxlzjxjLXkXrrplYGxcH+V7TAvXHlwJGEK
cCS087WdnBCat18Q6CzSPyWIsjldU/8IrIZ/fmP43W9pT0mjZtsUA0tKGe/tjhyC
q9CZ7fK40pMsXLSRIqSs2DqOiz44cW5ij9kmAmYm/d+DIbPmfopyQC2iGc/Z8VXY
dgxhkk5yayJTZoegGWI+o9i1qTFLoGUl3Lc9Odl8mFIpHpbeVZz7dcR7eHqXtLap
svtEV1DPaX6X9aEnRs+jqLDTM2PGkDvD/NW59XCw7Qi8G6dSoPC4cwN6DVDMWmMV
tvDPGkJIlWRYVavntyMqMREPQxTE1FhAVVhGB+KpqfEpZVVEWjHynoCt3Cz3XOMk
BONpVxEQYAZ5hFip5AsBjx2CB1JR2uBDeOkUx4wAaBSGXAnrnDOxE0SBQKj0EKLO
sHsVBqvhSu3p25+zUSedx3L0oI6JcmZEPmLNf9/Ku72YpsogClQ+lEYzAlOnidzq
n+e7WGELLulyo2T9e8jfyL4Xpf1hmrVY9uE9UxXL1pGwHT06a1FZRTM4v8RFi2Fp
SXhQqRO0rwJSx+jFVjfffq2C/v0FJ27Esqlv1M33kYp/Sa66JL/+4Ps7VAUDAslP
+vh9aHCR1NWiEfONNBForxwVAvv6r0K1ms0X8doaz7M+47QQg7Dri4V1TZR/kxv3
N44YO5fe98TKrbniCiKRDrzHPGlytAOozTTuW4djMjDu0H0YDIDH5pmnB09X1fBu
JWxT2l6iMp9BMHYgxZf0B79oOyxfW2ySIC7JXzpHrx8voKJ5grbArFtTgL4H1TkZ
WNHPy6n6PzI+7ZwIYxi6Z5kllYMecJ0gOEaRMrd2Wg6wdPFgjqh6VuMkHF7tU8eW
uQ5h7042Z6o2DqvXUZhj3en0Ehz4IdM5GMoYPjQkzwXUZ4IxQj5sBZmyihzNsxAK
f0afVgi1S2BwbmZCiYMoIp8TPdnajq8M8vGNUZdJd7UI1OllKyMJxaf+VCY93Qrh
NSdQpgPEU/ZwI9uJIB8u6KsyQAd4wOv75gdgv7t5ItdQzxf+4Rc6nzrkwjTTTnv7
t/apIMmB1GGF3QNIw7s03ql+66OI+IzZySXrkb7jVBqQzbKNZSwc0aeoxkJmv18N
Vmr//F8KV3Hwzs27ZuY2AaMyAX4b+OCCI7uVo5AtwY/qEIX6ktw7eI4jouUIhKHl
W1R35LdFipApxFybIB/wOkVeFT6lRqkTg3FjVnIWAtjLP4kZj93PL7WVlqs+VyNk
qdQiEAx7Oafa3rAoJ1LY/Jqy1Wq0SXDHwGt1/mSMBCzI0bEqMT/FF5leUVvBqNNJ
DQN+/kiCTLQXklPNn4MsA1pfVcKUlkGtm7CSpuKVkkc6hw+ZD7icC4ZdOLGff7OW
C7DyvnP3oWyeJhXo6qWTwXPr/Uz7hK4uFwmNV5u8GXY8H8/lAhMM6JGh70ystK4t
h1JtzXm6I2hX0r1eTcqyhg8OWi6CECF737DSL5/F5dSSp40ykDJcZ5ULmn8RWTOI
MI24yaUNxWq8bS6BKKXDtDGeeEdvGRbKeEYnsH6Aip6VFULuzBh92jR1sHOdR9Sm
BPsXLY5PRXKiNmBgiXAL5S0BPvTHI9AYCraKtwErtI3pZ+muRsfr0ZUQ4I/4qfly
gvuBD6UhisDaVCk9VRhBXV2rIYSqICtPQvAePRt9c4I0rKkL5FCYGhEFii0W3kG8
hstKlPvq1LznY9LlqxRBAIkh6OuPhdTJOIC7QnRF59txxTSUYHEwtRmntuxQEdC8
JIfwcGhC2ei3BPwNbezUODcHJSCB3qr9sIY7CKOzzM+rxUqjiaQ9oioE7b5V2eXz
ZbYq8bbIh4kEFOJjCZ2uDw2w68EUG1LSHH2cuJF5PdTJyCSsp3DQTIj3N7mpCDlR
PaFXHYKp4D+t+11TexKCiarNWj1XNzIAl6fEjOhaE598PSt4TzGzG54hqx/zWOxh
2qF3hzNmb9vBkvHobFXH4kiEELo8cpBTHlCclZLcWgusfZ0rdOOVbrDU9Zm6BumS
tAMxnKSM5xgTfB/LTeQPeUKnNTdPsmvo6Qp8ZRjjAAmWSmIDX+mjrcK/H44vp3MW
XZmtOgV8dce4LvQC0+5pIJCxBnlS/71pMlyJwALgsiuhLBxBoNZgw0/zrIc8xLp2
Lg2L3pEIb/SEu8fo8rnI2cwGP2L4UMIv+cfFywhyuImytPvw8lUnVNHpUCc+q0rV
9vrTESDe+HD+Nuk93HA0KHR1RQvRA/xKBVa1L7Y3k871vTf91lqb/2PdVLiZxocI
k8R+mBgYkm5KxhtAndJJvxa0VhMfodi4EFXtk7XINemi3qLltFA23C/oV3RzVJeu
3nvGLKIBmFbll8LfZF+ahJb75th2RXRm9XH0Fh48FOeAZMmz9r4r+9n5yFVqmoJC
UZ91Wqa2szRHT4NNKg3cH+QG/rq7a7gtr5+71Rrmk9miPvqWz/ajTW1NrJv0Anqw
vDs5ZD/Kc2dUO9yFsnA0KZnixPZRjBBp6njsQgcnIMkzjL64YeYr3V0pyQ9Gt/xB
8WbRSfjIganKTN3JcSTW9lrvc+odopqBAhgViJrX9bMRPIX68xkK6i6Gvo8eUQzw
Wk/UzMiG7erwk6NXZCvkMECD0GjxoY7MyFhdcls2RGVyCEym0huWdwpD2ADXbnHt
ItR116HDA3pd3xFTv866v/LhIZhpIVs1tvjtI8l70rU0sbRi8xWbP0+b7JIZZCAP
2P31vpSjTJ8I7ThkktYxhkQFsv+q7rSAZD3qkaL3QVJKXZDUFGmbLovXzA2yZ8/p
0PaNp+JkcuBGYzyD53UHTwrqenLjXHroBSGd9hSnj/AURptWJjFidbwoxtyhCUBE
HKt4T/un+gjWYX6ZPDtmiN6hf8UBSgfmzMecveKh/WPRfcIs07S9UKeBBzzeZ92J
SwE/T1EgQNGiBJ7gW9lsllhJ93WO4n04kmrMe8renGu7BxsswWpYaqX71XqRCk24
P5qlJOWsGM7U0hkpn4Rcx0nlGzR+EQ7NBXz/K1kY2p7jYUE5/7GeCt9pNaYGqTE9
68jtD3ty6vx7SB0GmUQrDyjqWPMzmhzD4tkY1cS6OQdH/NA4OEchb4XfXrzimg95
iqdbHJn7gm2ACdvEXjpcZIBp1Th4SalLgjMONw9HDbb7u5CXlyA901tfBEmRxm1D
YvNldtjJfITiIzbiyQSqYEemGAzqCd0+T5CZV1YgaIY8gSsXSbJYEgeL8x0y1ZiX
i9t1vaADcHDvks4Gb7fWZQq+2p/AmhQYPSqfrU3jdRPA50bdw5d47qq50kmd7b18
h+QCz7USej+IXk8qFohV6ZSqPitWE4XJ6v4IGKirslZKdHjyc11bmUS7eKz1U9qQ
87V1PkR9GFgo7Lqh8hwOL2uVql1VHbOd+7QXumzjG3twcWVdWtHf+PbNCS/CndhF
7q85t+/8UZQgJuv7J6Wrd+FThlUIVYDxrDS0BPrApvOFcBo8Ba+aVipi+ZE/XY+T
HpYDiMy32ytGpU1mvC1mp6i03EExEXT7+0+gOtAybWBPRj8KawBt+WMl7swjYCMV
945JHN0N0lAL0C9jbI34ml/SPcdX/M7cAaZ7z7oApt9GR4yblonlEomXoWjpy/lf
8Vl94jhXrfcdYb2s/FgAx7zLO1mq2jHB9tWAizAcRzN5pLKbSDFynxohUhhlUWZn
bsYe/Cx7z29/akFfiH9WdOJeAj+1hJzWiS7vNwnxQ6x0pC5onDjl6p58epBQOCrq
kQAtvbx6Cd6Xhx11eMP2xXpamOj7Mx2w1+z8Q5vXbVvv1+QGNXEsllSnXEuRqkza
6APKAsU8+B1REMutFEScRp8CZJyLjsze2yRwLXBpH7/YMytzdLe06Ghq3Cf0eBNX
/TmubYI4/ZFMYqx61Eyrk41Mo8DYynL7e+J/zGmTLHeBSBaXxM02mjpkYN04yFc2
gJNHT8xdpUOZZ53uZifSQW4TnjWiQmvGhkBmD7zAmRI0cy2aUnezH/Q91h8+3d4I
/i2WSfiCMIKOSamG+zyWn/q8o5m516ekwkNnVRkbHttBaZqt+bSMxEJGifU/bqfa
ekw/zyidMgVIOvHJDKkg9qULX6QH2m2tg2j7zNCznSC7QifbEhrnzQfhmrjgDOuu
MgdwyQOFvkP/kbUJ631xaCgEZaxvigm92uZht3WGlwkKbxThAdbRYjtBxmfni84o
5Bu1yEivqnE0++tnYw+5NN72IVEBYQq1DtZOBwS+P2ikJq9rh80h4u5tlf7aBs2l
m7krWtGTH7mrKsVk7PTnPCUM8VLbioHfzeS7Q2MUAzDJa1T6Ne7pfkbZCfub+Ad5
AR1dg2vAsPDeTrgo2RW3hMQGpLxqrpavfbjQ20iGL460BL9G0M6zbbV00kBnygBp
j79/qMBbHOPk/MUyTZyQRLj+3GppehBEXU1OB+BtvwNB+g5RR6out6T6mbCSYYYm
hU1fmwCE3ycaT4imhg1FAoERkp+oGWw6q4xMwvszWaFR2lZpM5UytazO95kcxHrn
B4y5d1DcUXo6Aic9Q2fsA8ppmchlJKZUBbzyDR3x6ISIc9jk6zekewzksuO0CSBt
pfaY/ArTllnPmGq9ZFxla0rpU5NjCiQZ9B+f8h8sEgtd8bHCz4pxUSc6REHK1X/j
ojvFppbKFKds4HCF9i++4DBseXm2ANhMswyQmcPdMdjjpqyEIsqpn40Ly90xqLl4
Bw8jK4hN7Wrfn7GhQJ8Kwx9Nx7J2wKAYi0gaZmE+40BiVhSGvGVekLeUVmxnevNh
Wd/vxAsSXYsJUgnlaas8cFD81o8HzZpcwxZWVj0CWUlCXq/k+jkcCiqbzOk5Ylzi
dFITcpFoMdZgXPAlGrdX+sFfriPiFbjaxzQtDKat35pYshIyLCLYJwH6wQx/Hlk9
NwsJeaLuFd7Lyb/JEMYvzLhmybHufOXhe1TKkHgfMXPke3mV9GXo9V/wsgTuyUUg
l4GT0z9Cy8C5wAzPiN0oZan4n8DBX9BfVf3BAClb+4lTCihuKLghvcuMUlRfEXy7
S9LwnAclu+J+lU8IcVliP+h5Xag5JaAeFwgSlDQ0oNWyXVnepcMk/t5kOP7AeUt0
59S+4Vo1lvGKVI0UXTF6infcL4myLhi8ojM+rlhHI4rgegOd+XMcJ9tYjbJ4SdKs
4B9+l7au4rDLYFEc9+YtyExn1CHfb1i0xOBWOoIJBI4tePjzbKkqfsKMyV5wr6Fw
4zM5ykkaLyxXATBf5s8ox0y8g68rBiegTSOp1dJ0QoyleSfOBihYRLI++9zCY9Kq
4n57LHMzcgAAaze5oFyldZs3cVPqoGYEHFrFv46lqkNTIt6ib3jYtGW3RhVZsvVQ
S1+KpwMfPMPSvN66x3YXCMHjBWYScq9FU5LhLc4H1rbpBPi6DjMO8xo+YOs1dKCQ
cphuqefsOW9C977DNYUZjDurdh6+ncjLWJ+WNukKSlaxN2WOsxTDh+ioI1Z3lt/k
n027HsJlGAKmAIRRk6JsefsLmCuF0DYgZu6X6eGt6zaloru1oYZS2mecUcpi2sxZ
5M+H75Kr/bW41IW4C+szd9luekdav6OD9M3FJqa1g3mjLClFuKgrlZG58NzcQYIV
IK9QFXtRS+4oi5ioslaU3qOH6Wv7f8o9qMNLZbPyFeRi41ourjhXwg9WuLAh+U6U
KFbNcOX7H8Ncbxnt1mdkX408Zij52DDsFXKgqV5cMMor6f6g3z3w2vM5e8hhoYUv
yI8+EhASYaEOzeFSO6Ap/tndR44xxYCsLhFj1KJNTWKjgweSuu+Xe4TkqjnC9Iko
+3Q7gClqwS4WLGFQHl3P/sanVH4M2j+OQacPZ+p/3olX81Zb4QyePcA+8/DCb/bc
Pbnp6kf0sa+Bqa90IvwpfZGg/KYLLxDqmc0O7buYgI4kUjxnHYVDv2HB33R0ZDtN
FZ6z7jbFA5Hs4Qs5v4hvlDzJ8OIXJWMJtj0fNnMReF8eqOvfndIEFu3SmbHvhc5H
EpiA71ORkIlbLrhZz+mLFzIueuLyuDktba/3HBYkKLcgAAxUPZWjYejtO105PQVc
GtHGbRXmrVrzgCeDMpOCirg6poj5frA6d0uHU6JTBy3A8EuaBBeEnHn+Z8Z9K0iw
KHcDYrx5E3F5ityi0dW6ryyxDijBLtg8aCCHHkeXia1XN2ao7BfUVg+H2NAh6Lwe
30Qeqh9aae3C/LxlmEBoFJAgUAi+tiO8Xt7+z805AxTaa3fVDcNcRzpiCoI2WCFk
tnM4IB/jMq5Ndlm9bfVIHJbxa+32OW78meakkas0FiU89AXJf+r3znPrQwU89w3H
Y9RWW+q97QaZqo+qbf87ZPm955k+QY44/38IgDVzY04tsI3elKYDp8gzwfXuazI8
hn+Se3XbhJe9nIQIlF8l9tEIQ9r0w04J64dUxMFIspVB5sHBYg1WugWXM9gWBtJv
yADBpVd+MiHDK6Os1GOh+9p+9cz+9p5HQyqEl6D3BPBRztECdrdhC7ik5InQjR25
mi6FEAYjsVK4NnNLjHLn24xRFIrBKd81xTbBPvJ4NWf4F3Eq4Sov0yHucHNgJJ+i
S0wyBZ3k9lZNmTKYHUvQ8J3niQ/fSfk06rwvT61t9Jmn4zXqGEgPO8X1QNsSzaNV
L+p4qoNsjw1ujfAW+RCU76iv/UHpzZwbNu1pV//eLuM3Ry5puaiGUIssKDJqI085
/maQaj63KhV3Ylkw/N1kvSdEMGlTNYDZUBjut68az2s3u4T8DYcFnQTRBFHTLs6h
J09LVo2fu+cR1VpJ3yq5lCajWhOe4MqveusUwL3rFEDCNVYWcgMFlTAsq/OzGDUo
ssKGnUnXxTGN3Dedg/SK16FDIoHKEWlWy7RwRSeV4m3OLGJ57WBwSTk0+TuWB6Q3
iYII2Z+M6B5qm8ADSs+0nEgETex+U+ibYqlgNH3s320yJO2551XAsT1W4LYExUwi
grfTs4sBLhLXZV1KO4/2m4Q6I3N93FHkqWR+rIPci0vVCD+kZnEl0ICWCOKu8U/Q
lXggqirkciBEW9Tgw/BXQZL80NdK23qW5M+bGjTIL+50kwd+GsFXrFqtXu3Dc/nB
8q6xS4SrtRf99sQjNNskjC+ylGhvm+Ma4z3iPcd4cJp0tIEVDG60I1uO0OviOHeO
IAmuTNKiryRe9P+9d5/N8ToB0axFSwipTSa+mDZjhQ29n7tFpyZC/MQLvJGsv6bo
ydxyFpffsUEukBcktArhgWNa+9gXBtPkmJbySQPiOcJ95jsZ6gUD81hCcP5YoWn1
Y2ffXETFHgzK+CXs5fhdiMXUcrb++v+Tbh49ddfWKkGVt55PjkBl638WpFjDMqJD
xgACsqmKcsa+dKGd+EMvAbQLi2ZSWm2BVGByUfdue2Azt5Vctn0j5abZqu224ChJ
ecbTJvFsCAd1Ygfiw6enBGC5PoABZLMyGGSitUuCL423jYF9J7F3+3DUEV1O9UA/
iJvTQ/+T91DLx6a+5U1MAUToQT3Ifm9L1yI4N76M4lHHpjGdaewByQK7CH3OTOPO
BXqFaWmA9T8RDRBvLp/1mO1pfUKqWUIudjdyghUgM2BI4rO9Ng4xWv/9EWtM9+Xk
V3fJdoI0G4osd5+M0NfLyBioBJiWUA0BeZF+7BKtXd3e0Ec5jmXxW0mqeP32enE3
2KvO1R8FeGCSswxu1LRaenBh5xSdyfboQiZKcO5moqwEPataDNCe9ewG+CZVyhqd
8CSMaojgpAnh9yz1YUgM1H9lIYXFQOCm+xAi5GU8KU4XHrvag6slk+5mGqorzZl4
B+Z15e0RjJhwjvuGjg6vsNxwlpqzgooqTdWrG8qP6aWOO2EYENDAgTZIR0CiphzJ
TbTSsuQ8gemObb1zb7GsV+xcAwkpLjSj6iGlvASteXVyw1C1rCtjXJUyATg1I2aR
wPw4xgafvNwLYrTa6p7XblC/HYVQKDnR368XPDHX8o2X7dGtqQF4zMrwXsLP71UX
Y3LqPFsCmY+20P+bxeoWXvZBuxsbKFDjb1oO3mCI7O5eRH1Ic3cHCvvSKSPaA57C
DKNv/Hnz+zuBrMa1r5s/i8TzGNqvkuat6/KE0Tj6us5nvYjvLru88QZflgY+PyuU
//NaMVU11RDUd/w/TA1hUCGg5S0ntavF5YRagGkaWviV0baDzw5XAH1xLbGkcige
9vWv9Rb4wh02JgrgX27/thCF6SYzNwt/z2BmPxf/b2UyFRlKEeaGbpLfRexIJdri
4yKof5P4Kf2mqciRKyYeeEYEFHXrueSbd1UecJD6TZdsPeXQiuELLg5b1qW/66nd
O08xMuXNJge3yX+KQ6DF/d2UZoq4oCE53JQB/hUU3wNcBw6VUlSX/NZ9xaV5uXMC
OJMQlpjVlVrxkbbxBAyMu15wIk9INGWhUb2Ler03H77yH2rqidGlGYzRb9fXIwth
p5HZ0GwBg1SXc2nwesNr1CAvf4cOdbIxYdT4yByr0Qy7Kk8Ct9HeeB5Kmpg0Vig7
0t7TvBvc2df49IKFm5EjdYfPSCKJc7GCtZ3OLs0Z8XV9oqJtJRgb84VDeJ6DRZNe
T69tIPDxjE/JwpUmlgEzdLuJ/k/ShmdzXHm2J4s2M9ggrmlnB6TCJJEwew4onARf
grbdXXLpB7DqyPAi02etD0+0CM7QGTSrzskf1p3QmS5cHOOiWagYRjNokQoyQVM9
KjAY62sHeTiqOPvFbED9eoXNHhj58qsy3ix7Q8Ef4gOFYzkgc4h5+DLWdGLttrOU
0CKlENYL7jsGNpA66Skw/aHXXqgfR2MYOtHMML1Jrlzv4sT5HPeEOf6Jr9ZaTk6+
8653rtblzpnf4YB+FNUdqifctD/91/b0G1EC7dKgM3es6xop+XSKYxT5E44/IgLb
LPhcddNve0irfduAAeDBC8lCuBts/HR/b8/aqtRTr24PmdmcrcHm5ImdqUj2DJ93
9frLSSuStxLZ1nNfzPq8QvBKolk+vGAiC+Cg4g2+/6mnih2jJiYdabWkE+TT3Afy
O9ucL/j5zUrvQGZFiY30MVaJRiWGPuCDqGm8Bgy+dO38aYHwrdGsQJQRuQJlqMGz
rGSCwPahnRvIJQq1Hle83Ar1MUkduJKRCEBb10Vhkd0JWRI9d5OdrYICbkQR0tEI
Js8k6EBpp9pEgHxLFMXggXljTLmXSwxX1uxtPp0Z9HaPN+VMHBhJEj38byCWqvn0
E9gUtHN3Up2x9lxeCnpAnpPwtvLD0E+jz5KwKgOmsBaDlUB5f2lBgk5lOgr4Qu5y
osBsDclzI8Xl+67s1m20xwLmTgeEfkwXvdW8WnHFZBspfX+qa39WygBvqYh4D97H
BmXh5seO6JLer+9b8ZNHvXUs9JUZiss6Sxh0rFCzFaTuKtE+3+PgPZ6ccvqnFePV
w+ipxEPu+oGJXZzdUE6pGVAXakWcCm4klJ31CGndiNrX81XiKKBTXxR1UwNu31yD
eYF6fz0DaLqAThjeO+YI+9K6vumj26V0zVpvLvCZMvf2iXd77JvHIynQUNyasi/J
Llk79zH18FCvNSS0QUoZRSyPrrKzwJ8gHzGqbjpfQXnhVtoA+VT3K0AiC2X4M0sG
jyKxJS6I7gKobd6hznfByu0BdJT61Ojp1KgoauOwB4Ocvlc1/P68zNCCROLkuUja
FxGNdpYBi5F1XZpHL1jmCKiy9oth1Nl3KUSrijfJumKCxMaTNC1Z5ij9Zc4vC6Tn
ilQ4bInlsm/wfVOD8I7bcaJ3kcbz+Dg1U53JRx7RNzWnYfg3PPcF9pMDWg0mWUwo
eJPdwxqZ/MaJOFrwxQ5AmCDHOh+Q+aVXRYAsJ+gjudvidDqed46tb+DAfQOfBRkm
1l9MMY/G6eViDez9YDZdU53n8U95kTF9OlWEqXfu+gh9DmjAXX9EcWYGZOLXsyZa
PiuevyTvZpFN75WLjxmZfpnG5jMPxtAW1t4GJnLUBTqfN8VBNlBMSC28G/CTn5jV
GH2F6fBIwsiD4piDa1KO++RnJPy/uzIfjAxOu4+71KA95j/rYUMP/6XFQWuWKcz6
eoRhDosttKsH09KOdg/RENcpqDinURtWMRir0zuLvGf2pAzv+YY7X+mUD6AtqFZ7
o5HxHXBT/oz/kDitFMSypHS/Fomi/KuA0R3OsJqYH23UEFpfke+Iy5GMLnE0V92v
djYsWEIPb92oPumQKfXQ86vtRXisZXbKjrOQG97Tqo+ZtzyYzrG+NekRaYwLXxXf
AqY/bYyU8szNgEPu/7Kf265Qx2qUeb0wIxK2BH3fZ9tJ5pPNCTwTh64P6y+kpk7M
O+dUoEMYadWyyZTaDhIhGUujwRjTfvs6kJkPlEiP3h/yKnWAEW9SqCsCGCfAdQjy
nK9Dy0UdbagkwdDYyZ0xajqqF4Sp7/Nu/Lo8ztkG3h648b7we2xLM1aCMpkskVkW
WJPBt9xNcAlaMlz6w+cvWWnnykja0QNZMk0GUfa0/UKcwuON/6M9NTPHqxAXfEw7
Ob9Rxse16NaQmOj9sGptKnkO8Rs1azYHdm1W44LSUGO6HrBfGNPKyY4H5briS6VH
ukQUY00sZnngux6ov/8clE1n9iZ/4OGslmkmtD9XPU/Q7vQJm7z/JEi2/TqZJXP8
ybI52q7Uk1eMSRahH0tCRavVGcbX9ofdzOEDVu5qoFACmQ4g8boYi9zC2RWtbv0E
fvtEfnlt+gdyK593Mv7HF94LXCS0/DYlknn+k53eIlqCjip4aVkQ7+TYfHCdlqL2
BeIVeW7oMprqwLBNrbhzq1Y7nqyec4KCCaz4Kjp83R0ocY986UAjPaM9LYFi9HJS
zOqZ0pcOPGY0TTH9zR3Zp8YeLJx/Orn8tYlGC7aq+a2LVjEBNdnlakqm4qG7yIDF
q1W3BZ/FI9ogyHORILcMYtlrx4QRYbqiK9z8LOZ5/jJkXl4qULME1w8fTC8pHOQk
CEASWzSpRpiGbqKLNHxkWQq2yVYPMn1ousipRY4gEezGPqys4yDaLcqQYYhDhRJc
FFveTiPWh6hy4u27RJNn0cqdmldgJCuLmIaLNtrrOUxeDfQFnTy8pddCvvhCruH4
f2DcEDb0tMNZHX+yiBZWQLbewt0KszlPubgXKmdfYOAIbVHqcgQzeuY6tWKuGh+F
aY1Z/nn52GkZQDMUZhes6H/4NwV4s0k1gM204rpASOdjMZO9vPwF4kudb09fv+L6
pkfSugJAEMrxf/sASao9nRgQRFJ3Goy4nyTy31X29AJ979Idtwb7mWHjKkudbq/r
WiFl+jTISc7AY/muUOLlRk9HOxoNYDJw+/iSN0Tl4ODToa8D/NSCzXDXHQbG27R2
+BKgbV9uCF2AN75aekZsPHsPZ28CQXrI8BJbgMacsXkK/RLKr9myHBJJSGO1nQK7
dHARasPcu59jU/A3NRDQJd477s+pZPrCfhWCDMZWJzH7e4aLx9aLpwQh1IPXlBEy
X2SOx4Q7UPqM3iuTWbbe+V1WElPyqtGjjKhpjdZnMtq7MSZi2K/72LLzHZdd7Urx
vBXHmUKf5dXQVtj39nwI9BN2ciD4kTM1otYMT8/M35ZyDIUNp7a4SFxjDyr9zaa7
NmUk+MZ7Wyj/dqXfSwVMUIDwVASDuaulFoWOS8rbq/6g1KpbKDX/p0mEV/y0HX+d
ls+Dlk5kxGDyyRwhQLFAbVM8UfpIuHKt9Qc6WUwB84mooMwfEWiQYlt+82B2qPeZ
/IR2AKoZRG59GBgauwr1d4gUyrt1Ini6Fg66ty8D+gfif5pfeyuzmFA9sYkD1RIf
0azkAqEi4BFz9Ymg/7NCR6onxtPZoXoea2rLKwIMfFGl9AEK7kYx1EPJCi7LMdEU
3yhPgGUn+LyvOXS/J6hoTt9MUOlIAwMOS20eR5DYH73JeHfA2QqeUEKA7vNWc2IX
QysK02AivkA3SB1V60DcITo4PnZnf1UmqFGA4mXRuWGQasvA/zaGRkTdUWtCBObo
IbLOtHN2lVPpZzUtZ9s356J+HOgZSBpVwLLCVSVGR9RS+8aSkyk+wwQTZHr364Kp
ELgR5dAhzevd/ZFCupP3jL0thO1YKStA953s9ncVPNPYEgh62GwL6kihgIZbDxfk
0WxVPQO/GECrcG9egimX+neY1ycWgggx6c4ih15DFo/R1VDyxOvcJXV3yxV+B1MJ
V7hOhiLhKJ0fx4Zk3AtrnxRC07KZHbP3A1LIg4vxe1Jrff42gDmKfQFx2TJw9rCU
2+WTKMiHmobo1Rxq1mfV74q6voN0pmG+c2OlE1iVYq8PnMqngWuJtuSk40UkdsCy
RxA1I8+Vsapjnf3orBFWgA18+9R+tqKwN0e7J5Py1127Oc4/pqw/FMwOQtidoK2w
gCr9yayVHbkUP3q7/7pb7SXVVaiwObXXs+6NbSNO13wpJlTVMUEP5EprelwQDH/S
lU+REvkmhr2zIVDmeO1Em8MfxIIFpRU749UMDbegxyfq4SR6duvnnsUb/7fAT6nG
58Zr9XQPqcYGb1ihZ2kRQGZmryTd2l9o7r+kiYobdol+WHfHhiJt62clCbE8BNhC
/oAkPcnfp7mMeq6T81qobs8+24ioIowtnnJQ8/mf4GxOm41EVh1dcJAKfHsGJAnu
omHzsHQAh2qavRd9hLHP9OpcP5hUBHHTjzVdNd+I/CXNFq5QamdkiQTxrDyehsEP
LQkiHm/9ySGQmKdhja2TN3Cs2q9p7tB7OoviZw9xf+CyBkEZEBKhiDeFElsF5CF1
n0dw7r/hSTP+THjmFQ5sxCj+CuQqfo9rIJeBs18swO2VC824cwlhreIjXB3Uxkzc
0cnczZs5SS9PuygKSVM65YoGWJP5C4i7ZcTJwAcMlMrAKOGH7sf60WQFhEnyhznS
eGSWNxJxhtNLvAeYpBm9TK1RUnFPRc0g/xkUlGmvyUmD81F4nOncLvr8StUHqMNM
19VFN1pA9d8eAxAZOvyGjapEg86QSLR0uqWSc2/EVufEjG1XGzODD8Jlk8uj62I0
8Xuh8Qi4rFm3OeqWNILu1CpktSP32ignZ4KdS14dqqgkue14F/KisXp0m4SKhsuy
mpemCA3CgTubDI3Zv8ym0fuxW8YzjRJkd3CHiBckqadoC1AB2MnvWiOLNG6wrthv
t8mPGW1E+Vm/uo83zEhthfK3v7K/GYQSY4LaFh0irvjbJqUMYeXDxG2FLuLNHHot
FpGSwomZuEMY1GeLzhgXlQ4XZg82DEc9SbPS8MeU06rny9DmFJsTHH4IpbN3/VII
Qt8SZWroPZOOwowlS1vQA6LF/s97kasd8WL9ql+YZNf+R1mBEsknbRoJ+FIEKWGs
gGBnP3nouAsteiM7l9XpLic1X4wx6B5A8cqmr2X5rR1TbXXPssSlB6R7gGNMURrw
4RQclE5lIuxL5SFG2X2uFo6/HTHCSHaXUKFSUcs98GmEDAcvMOT1GkNgPjEu+D6j
irpPuCkT0tZ8kbVLZ4LgCKxMuJqGCqMMrlUXjNhHhqrm6UvyCMWKk/rSLLlqY3oH
f5tCsB8mRV2D9ZPHYjkSvmacMePLZalqMbd3/GIrMJ1sP9n0Kw3BjhSn6vF3jaBi
GjNO8TuzjCZrjnSVnRiSmBKEg1RPR+J7Je6pyn+gfvWqvLB87Ta6+lnuSAtLOklB
R6+rfRJndc8GyifVTfGODtxI4C/MEeJNoAGhYybzJzTOU7lu3jdalvlh/FiI1k5N
TwzCFHnkzMzs8QYr7PRz8wIOz+er0o1fyjfrFZmehacKtL4yUJbzo4jmk0lxvt8z
36JTpaKzJS9TogK34lu6JJEe0Uoeb4n+qbRaJA+DusevyhGThOnm57YoyqCzMKYg
81/GT28rUv0FErvYs+iMdBlGA7uZQl7itaIPBV0rggauK9uQbcWm1dnBWFktxzfI
DbieubNReVcyXlQGDrLAWoNRsHBGydl0vhMVB5xdkypLNHodIUE7wFNY3fXcwJVp
wqruMx1sNjj8tPb98EPyWgSF2Z1gBReVqGQ/OwKRcjPRUkvUB3Q80Nlh1U2Hd8IX
ARGydFCmH18wBX/zuUxutAH+2M1uti6bYzlnjySdLTIwkXYsvafnBu9DCRGjPYgZ
zfQp4AYyHxa4zTTTd8omJBtpBqJ3vxFy5+PEBJPy30Sm29JeMfMqtTX6FDK5nbvM
wuShTGYZkybvdrm5ohgIunehJfaky1h3pRh8+FlD/rjeKy9syDi11ho09D2J5OS9
T3JTc/cN88Zvxwh2REgkUTC1r7Zt81gd3zUzJcMBKfulu+EIM3btfvDmwLbLYWbd
AW7+llxHopbtRCkT6o+F0heJahKUYa2FJsryoRpDxg0/gkqhHWQxryQ4yYEa5L0/
kARoEabvqyBtw8to2XFzRUzrn9TcvYQf4MIef9LyEb8ZggW3rk/ndVPgIY2ZCFKO
3VaDMdiCyAk/j/V83Nk2HVplwtaTVX/MkIOz6djpgaespX4P6ly1CbTtSVTR+Odx
AHjYMGk7lcRuZhC0Ae43zIUDRtEYbtym5tzbmTVJDpYcchBuhEM401XWO55W3jUi
IQiBZhxnATwm1lluCIIaA/Csh4J1jCwauUsU7gqG37Q6wHGTzoZYYCusdi9jMJsR
/ovurUS9VDNx9eidygYgBTvJ+vrvlmJREnRUFD+//+zRYi1UWNH6euLz893HHecb
f5wypsAQKuOa2eDIy5wIYqQTdJlDkmFFhbPYDk+paBPOMLkjBCenh4xV7HmukRNr
sttnYRSA4bWyy9H8lwwGM4exrFhXP3TldPGl4oNT6NZtRXHyMeVPMCIshwfmeUo+
2QXqCEC4mJHtnbooTV/dJDQqlf8VQao7iUd/hmnuB0FmdBGHYBT2Qs27TXN3vdlu
n+ACuRR1/u5aF+DL/o+LGHez/zuIb+m0UJhfw9ANv1i+VOAURmXyNIUFbczdKHD0
k5F1QdszMNAYWUu/KXOxyhrqIf30BWkZHfQtdOph7jGHIdnhXE2oCB0GOmvauLuH
t8XjPw8VNaK7DJKVrWQ5FzbSQXKPdfpCrwTanGaqtk6Ua3g0/yTjbRHm1thX8cjT
WQfVF9ZN4PZwf7kf5shmrF+8Ok9u9kmepllVFQ6kGY73PUVn1C4EKVUV0LetX/Ju
VZ/f7PUGUvDiyyUaj9Z29+ryeAKD3tv/gZuUylcGNzMqJDaQ/QJeFYjuNgLN0zoM
udk5S6SZEFvB+Mde6rULhw5+CkOSMDSs7iUDwfiWxgC7nvJ99A6klAffswdx1C3a
r2XP0BgxbzgomHpX0wjcscSVS89XWNQs4tfEvBuouZW0N/ztYc34enKvPQF/nHGo
hGZACzSsqdzclHjcOFY3V9cKkixDmsYM0a+dHy+DrNK4XsreGFZTcqWCy1pOeicr
a2b75EbBOH399LZ++FZGeU9TvklI1PFjW0XIIOCIT0kYqkltOpV7T1k42VuUl4bJ
Zi5R5GQKjTIVvNbsiu69ry9bI0Z9J3koYKFdKhK/jSoIS9m9LUc4LuU5w7bFw+E7
mHf6aMkwo+Kd937dPCBnYR5ZrgwUAmik5fvTVRfJmrzYr/SojS9px0pYZIMiQF1u
5QT04C04DRSxpK+f1CPLojF9c7RbHxOgTLFILn+R9RNMckSuphUML+hqhDT1s2dn
+W/68i21pUqIRRgrCQadSUIoMfytIuc/Nyulxv7xyT3S5pYp4hubrKpTZWAnPiPr
hp5RYmKvhXSzwZ7sNS8mJ3f5EuIf6O52sW9JySng46KBOAspE9URcTGQSI92OE1M
jdp7AIb2NEdGgf2Uz2BMFgEEjf4Cx8/4JC7vCePlZ08NAxwvT4Nnqqs9HAoLz39h
Ez9JbmYLkO4Ac8AZc4IXwcGF92kCdXbQbZDVA5UBVOiCqqXlDSasZ+plKr5KhRdq
d3QQb+2jxTNbDyihQdSms+3nGM7ldCtYDaBh3bVhGPUWUq2KP0D3ELADHwjPzjcI
D2qd8OFrQX8PIV5Sdf8buYJ1+ysHur4p6Mxquq2ZcThwAkhvzvrfKbxmVDCLWO3/
XgHVld2yDa1/QvoAG+emFVndMOsYBO3ZprhruItKsEYpgtQGAJ+ZnLTAVngWnzso
BtscqUC9VqMxIMUxG19nh12QrR6GRJx6Aelaf3jhkEfgNXb6jEGC9c4LkFbvR8DS
xlilqREnd0UBqyTIlEuDj/EJLKBjFukY8K3i/ytp9v7NKt6yYm+v94gxS2QAU/gw
A4oO634dZFqCk67LQlIVe5U8mC6SfOVG/mFd+36zAXZqPfja1UieDJC2Oy0c92Oo
CZHp314KNFLIFkTeLnRFw19XNfvljlHnU8+Um8oErFPRi+1kIDw2tdXu99hcTkc/
xp+Fme7W6jLQ7RI8Z1DeuKNvNY8WiCoEeTVytj04bOmvyZtZAYaNd3gtIB3kVnHR
Wrd0hnL0kOuIzDnbQpEKAIsiQ/aT9Et5jxcmYFwAjWGmlE6QLN+EX7ALriPacU9l
7DUYwlqF5WTKNJm34TIYw65HusydbcGrsq4bKhdla7wICupVBrVZ4D+omklIH2uG
43KfjhuLEZwT/nboNlEAg9xYskkKlgaTDtuNiLj8/lu0Vs+R1Zvb+mp8o6WufyGb
+LxTWrVDRMBjjMOWQQIKJiOxON1SY004qQ3AgbGvMNQo4CipTHsgmVmKLta5Ct9z
ktp+LUYF7f3hlriOou1dC852uLr77oIYF9M1tnho7UcNMfU5ffMsIHdjyB7wu5IB
7axhHzcp36wvMITwBVvbKIQx7/t/eVI3ZeHa6AcVncYR2wG8fUYawqA+QOPiESNv
yfq2iTMDgx93SpBbFHPi2aqxcgo8oZdfi3Y9zslBNUwA0cfny5mJvImuDOsDZ+2b
qA2AsOSlsVARxP1iLQfXn6QJss2iHWBPdEe3itJuaU9e0GWhUG76WySun6mIoBNt
+jURDwl64o1Rhke01WpRhr4dLlVH7TmCdWgb5E0OEtivZ/ot/ub2A5fuLA57T+8f
PAcvtLe5g8NMLnf6pvKdvTLRGh5r8Gt4fRU4SLJSm9EDgJbfjt4KId6OUmhA3ODc
6yody5hFqvbBu30LUhq9pcD7ILq6W+QPTyQ0xXh0yqjIv5X4iOHiD4i7A47aznHU
YUpTZc5isCljmnZH0GLWfHOiXNNqGnSQcZ4RKg3WZ+6P5LiO9cvo3qofPVesOXCR
Xropwo1J6uwlmqqkWTJl1qQ5Tir8MpMea2XUYsGuvavYGYOegKZi7I5KGHOOKiSG
A1UlLP/ERD5lhcXGfcZB1RGx4VKLRjf/J9jen45eXW3Usm8aZ4zMRJoZlujYj3Qg
4j+uPV+pgJle+UsMST/OCiICVtn95fJoVrqScprwGvzUralSbvfVJht/OjqLK6I0
lJ/pDMtC6zTzUVvRoW+wFiQAOkfUrfD7diWggMqto4O08h+4juiDra7qCfacPRAF
k+Fttr7mTmYcOutPh5Jz3JrQpmWzCWsZq0qfYf0oTHuaIg5fuZbQvtNQeAH2k6rF
7jW1qzLZ3ky1dxM4SrTK5mRlVWRuaSBFg+Y+bhhxUS04fyf+XvXFWYyAKU8UKsWS
rfpDXGZa1fTYHTfTcKYDzo/b3fkFr3KIQI8/J5exwhmzbBbXPBbJ2l967L73y99C
96wsX5rQavgBhARGCkNQFfZejG1KDUUHgEYiypTu0rOzmNJO6LC6dIeGdilSqsxu
XL8KiXF/RxPjrkY+Y/u/ftod0elu2ywMFm85OIVdc2EjErZGfp8o+TU/4YSfEmNT
I3K1eibBg58j0Lr3wP7YTyvT+wGBG8o8TtqL6q+QmMztfRdwr9zkJXZ8yGZpkEv/
l2pKp8lvvEwvqH9qjEzELvJv+3cSPBrUWidEA84N2jS2SCijcEZ3iWKe0iRMLkt/
J1KLkl6wPJQygIQwDrzhNTN82PZ0sbrPVD0fwH3vKhvwZ/95DLwt+lZ4iMy78XRI
Inb1ikKlj+vZxe6vHY1RonXV8KM6bs1H9eGarFMwH1e+FU7C3Wgx63+eEWuVtU/H
vzFyJEZFxTuaywhmSz9Lr02Dp31VH7eDeMkvu5lKsIG+uYo9iZp0eCn6unP4PoV2
3VcG+8c8vaAAsL+3QDIrkcDadTjbqgQMx6T6/toIyeFQeKFeSzo7HedN7jeZM3LN
qqCqHNnTpR8QtSSY13sAsnVh5tRppHKw7/PyW88F0lpFXbtn1fUn+fpZ+dZ3/bfp
qMMFg3X8V56nKEhJmtY1WTwiDB/0m/qhgVajn1dpeypo9l3/NvKsEOHFj4HfPV6T
EeYu26Yqljeabm0Ah6a27r4B5VrUvre1i44umwlSOuaQ19wsmzh0ua6afILZcwgu
byiezqzPd5fkBAcV9uxB6fc9pEWv3cijLrrcPUxIaoyXip8b62ZWgngXkkh0OBHb
9veJp0nNH1A76GmMRu3uAVV1GOn0QjmnGWMnI3575r6wYO8ItGHITeDHjrXOrNBA
izx2FqsciFi8NWYE/sCtxUJDxhXUvX7et1E+XKIuBJshnKpfmI19xLtUi6gn8//s
AuNJzh/s6S+ZTwZ2rh/LGo6xc5916fCc/9TrNgBHk4OmuGaEcAZTc7wyzl+JsuAl
8VLUpcqD2Z5hXylMYuj7PpMQ89i8hXq01srDfe04G/oQGLDahUrDa/PQYcmJmxCm
yqkcvf8N8zWXF+w1czFImoX6ZOL/rojwAh/EqEAwoSUOMD5a+3Ll5XZPeX8ufOT3
ntRFzQC4SHfmIOB5VPJuQa95u34XU4mnEbxwcyAT5XHmvy2IJRnSGTWYyRP4iGf4
Hn3UQ7rIupRcdBqWOSAhOxSntNoT7jKjoYKacxos1nd9CjMb3CFBl7KGugZSlIv+
oFsqEG6Wa0prSKAVVHkF28jl2T/YqdXxnqGM9UkCzzJT+0BtcNZ71Mit270sKqE9
7fLPKpfxgu79z3xEi3XZRBaG9BuDr7enjGdtsJLXgR2tJDLN4WYrPGWbVIIoP05d
9l9eQdzCOjp9mrZyagX+m4la/cQkwrNVbKTfT6QT6ocFKH82oH/RCGVr1BBlfxr+
+HfaLHVHmAGbfYDZz+cbxt1Xg76ablRMmYEwB4Y/Fb1hOB0CBagO5JmgWkbd6R09
ot+fV37BQSMZ9JRr/8lzeW4tPB/3NzorQ2IDOTY1CrVZ/Cd5h1K7vMsQvaBLSI7V
fVQVImXojxv4uofeinf7g6BCIw/gejbsL80CgGUyXVe81SaCriIwPBO0KxqVHYh7
yDHJXObTJVEkgOjFHnRhNvIDy6SOHps9koP9z/Cu1k8DXldM+b94ksI8o7dfwVQY
7i8uxopPkUKNpPY65+DF2bjPTQeZCPQuZxGjyi3BC28gwx8SLuRPe+WtOipMdKi+
7Nox7O82v6imoJxvZa4U0XXSX4LYwUoImFvA0CwZjqwZsQJJX6HR3KhYUQGcOXRz
RzS7cVPOlvNJ+GIiPEZ1HdGuIkM+3Lr6Etj3LCW4XBqid9SOiebxNI8JW0RUoyy1
tVA/aoCDn/B99MYt/c9/rMn9LEaW86F5rBGRuehqDBKzhbHmdWP2Vidl+24xgQFa
fV9cnW0xaQ+ti5tLxRfx6rtgYq1dVsu78uxQ1rszP77KCNOBhpdKJbgcBwdw4jaB
NKvY3PR2JT9jH7C4WC8Y9mn6xtX7YuBQkB8NCjunXdRgJ/mlAhNz6f2AHbvsc+fF
5HgJtTIM891S601j/BSPyO1xwjtMvyClX2MhRi3/TKfTkAeHaTFkO6VwNAsLUmI7
366tpjv2sLKJXfRNBTTzmCi2UA9nHzfG8uELcWnJuJsAmLEoO5cxfW/9+XPLU3u3
neRrlEzd0CmKKxfj7GlW39Cp70OaZ9927X1RWZ9kU4uFuJysSmjiKDBqvJRIoMd5
DpHz3CYDSP5BU3QF2zu1MqmKQrudtvYbWpnMWHhA/mYl6LUqRs6Sct/fIQJdiL2k
da9ccwA4Gx7hX42w4XErZyyJIelCA3g2QfCnXZo33LTnoDFKrVvQjTE//RFyEVDr
TEvc2Mf8MTz1sEIP0LNnFOGRSpu4xjvs/PuR6SjAJPvqK2v0XTsUtF+odMRyD9+R
GzZWF6HrTM1E/CByJ8kpIAHdBqx72nT2pU9wJk9ZTg0QK7JIlQzgqQYPCd3TruP4
mzF8x+sqXJxHrJ8w3vHG2cFvm6kYB5WTaKaH9pITC5fxL45DQ0fZyi/tuNpVNzfy
+PjHrxNbMFzTdHjnycnucXwkrAljXUuSeVf8maomGy3WxxVSfDWIgqDpjTuwSSUF
7iyvAjtmisG5Y1uhc3KKfBxY0w/YA+dmi8bKp72MLswZDwfMRgxeaolcgOs7pq6A
tnvSNL3lFdQccBs/Nklsk+8ZRgV16+fCheT230JuGcYPcZA3gJKyzGDDapsSHHmy
rqiUvnq4bvGoDjoIw7gDZJ9G4QpT5i6YMqGkMyel2CFjHM528UxJ1Zly+VrfhOb5
XxvljqCpteBqiXWH+3Ew6CXzceZWQuCrS7r8ZmVcRYfLlDkN6Y46rnuXiWSUxyBt
Iel9h9Afna7WGjxOiACqthSDVQ44p4biq64SzUOeilrXF57Q7bLVRB7xPYvH/evI
zC9wALcg/yqhw3djdUtZN9zK6HUBG5DQv4EtmfcRBeFby4/2jxOMECKE3ef1qWrR
aP6mPB4WTj1MQAS+9api+b9V3lts8VK/krfF55jAYJTKeQWjhukSyw2plwRTZgDB
s2+QOXGdf0f2McYbkjUnbGbKuMbJ1oPKujX8B00zDQHe84t0vYnnfno2eAqY949F
uu6+iE1V83CvSGatUGVx804xfPetyzp7jQ61cvwlqSSRDbRil/nb69yWr8HFj7X7
+tm7AZJTzK6K/EXFUFCd0vijJ1Ptj37IW0CpX5jGA9/7FPRKeffaCgrjm3bXq3ql
4DoU1W4IRJPVZwPaPogUzyhFeNYBUIRqGFu+mnPpMMDSXufvG8PjIte9KR7yMVG8
XBINbdickbNYHurOUjcEWy4ixfV+tHMrjV+UbWt7d8XjXv03r2EejGRUOA4MTdqO
qygmuSV/5OJhXr29b2VYnPoRyC7XV5FQPfszpEiaukKjGAa6TW/5EGwBzTkGmWEp
IrP+3G7V3Nxv/q1CQnnNSrxMJnVALDFBDsHdWMAXIzCcxI5hIXMnrNZQ2VXZ0paw
n0bU0EwikJanSld8ArJdKwlN+JOBXZ+ea3PFNY25xxXOCfFBa4cHXkp7C32RnzZ9
06/vz+HeRbT17gTswI8DsQPuZe74MjNDALoyL0GgJCAF3R+kr/kKRddw/yPU3XIJ
JUAYlcs9Si1sXPN4/LklTkyR37lShmJjSQ1IE0YkUtX3o4o832/DHPzrjqb2PCte
oz71uqJ8m4sdaxEZ6BOwZDfeN8oUjAQBVPs+OB+ygUEtPiEhw1VuODfbJeVc43VH
vaTMVUwaJeb4Eh3B+lyJ87fXm8jaqemUiO2Tbuk0KpQ47gqmyyRhTrHTK5XaXVmd
I0esjfAW3rNiLxG0qHG4tw/Ebt/IEM/+1hRa3zLdptN1OhP1HIiRdTts8GTX1rql
2aY7X7EPTDxrBUFwhKdJieYo5IYbO3saPRd7fDI4XhxMiOI9e778GQLAeCAq+GWR
GaOKjUOSLNO3/rgzaNQ/jY/7qsE3Cj1OrwmqSYybr49++EmRZIbgiMKAY5YIoZNs
pNIl5zvyhM/61wZxIHfovpwx1bdFzPh/qyEG91Oq39pARPe+GBDT6f876RVuu+Z1
KrQx0WaF6vMnHYWsyILOuSq8oaNoMjGfVOuBZB2W9m5JbQD65NgEGVIAt6ztfGMq
syWd3GQ+ZZ+Vn9J11AyaAOVJ2hjyucLg6OtptzaZusI+5DAtrYOkyW3RMkFXtTA6
S7lCiDGhXaWnGoEn1Gm077Zw1a90guyGSGCK9/wVNRK69Q+/Na3unaidDKFlu+tD
zp7z+nGR7wvXdGiqpGjWAQdxCeIyrBBKKLKbpMH8K3BU/0BjTGpYgAS498O/Bm4h
PSxedP737Wk0kjMmBjwY4mDZHWQs13ZGxa83l9+Oh3yOQcumuFvIepUfgr6fEsTJ
MjnbpLjZQyaU1TqMVrpyf462ZHsZ8y4W9PtZbQtDOQgzL5vdCGRnrZC63g5AZQxb
rwXf4o4qRp2rW6ogP6BOQO8vZGo7h6plG0jL2YunCjwwUpJrcr+A/wtVOgGRmd+E
Om5vjeqn6neCfqR0JVWIxEYvwWxhpWW1gjci8yEkQAI8cZSL3m3SlE9Bn3sqR7Hx
l0Zc7uB7gsv6VQBloSnRwwpNKR6RUTEfqxhxFaqG3FXSYB9EYEqdRAlfajAjzOrZ
ESzIjp67cka1+DIeewaT0qY7RArMlAcB8pd5m1TrKJPcE4GRorQg7c5Xvf5IdBxO
lyTFQVWQeX53Xx8nvLfA1lgVefiD2lEkcsU8kociWPQaH0j4nJ0IpbspReEBz4Cu
C9K3drqY9qExQJCJ1fbYSMyKtolAE9SPeuYW5R6eippmPS86LALnIlSeCEo6vzUU
Bh9Nr7Kxj+r7tvP8naeFPCxCwtHqFp99SzKxNtfOtRdIMISHFy0b/XPMsgZBG2f2
rdhEJY04sKqs9RSpu+Hi3q/TTcEa5N1vjfUkwGJIgiBV4jotDIOJrWHpY6Z8PNwv
My6m79yh5Ag7ChycvT9PNv5n0PKwtz+bvmid3HIE7Ze9rWaCalIj1f+f0yThik9F
E+K6kEZALvxaz2tVbiHyHRYW0yX+zwWlRGzL7Q2mx1EcQBRkKNFVi1oR8+MhXxfa
aSs7zhTHwjsr4A1BRCM5mCHZIQAPgyDp8g+9+bd5c/FIK2FXm5EXOrjjCA2bvJgg
bo+i/jIK5EXwNiZLwo5Jql/IqDAjwqNXEl8q75dXiz6L0kP0fEykMB+U0owu36kq
0Qo5XmfBYpEXPVn7+BVsPfj61qKJLcKRcTb0YaeDEt5L6ksaPiCtuW7yzld4EeMV
NIMqkaaW5hLFYxkWQwRM4goVFGACb/d1SAeaMmnH3KUVdIQaVNW7FqHcX/e4sqQj
oP7PfR612QrppcvdWjCu19+gOwc4KYE9O+X6jo2UR1FNUcPvG67i6BNfWrG9oEEl
y4gxOKnkiVLIqB2a/JFy5nUPfnMeFeRFMStwJuNyY1VlJPOcPb4VqAzvGiuIhRRQ
5inkQX6/7xZDfAogvwHBF8qB6LQJzt4L0aEX909i2BRBxLi95G7BSbMpdXDggsbz
BU5DWxp2WzY9tZrnMtkyMlu+ZS23QQwweC6Hj4RQT+1mQKVF1XXVnRWDWpyO0Xzb
qiMQ7eGK9qkfBRexfL9PBNpL3HWeLKXc8nTvli28Oug0CWCjM7qE/c+PH2J5ROmD
6zNW4daB0yLHYt4RyezyGrwdnzeenoxU02c3GmhBl7ogFMGU+mUJnTB53GPjwZoK
4lSnrvpm+w7qnfNdTNn8F3OHB8+kQrozFQTOui/2tY3IJmOB/wH7xtroUMVREEea
DjY8laNxFvHrTTlIX8IWL4Zvet7nv+qJQbqdgAqBTBFiKXcGCaBKUypyuKerIVap
I7rrh1V7acYoOG1yc05dQ614Lq+tgKS71BtAN9cw8Ix5Pxc4ghU/TX0kg4EHUsxA
xXt926yQnfxQ7pudQvXQdXLHvGPSATQhI2Lm6Uqxu2As/QsFHWyoVRrvwrzYb7IR
rvu2lI7voyIfaQY5zzzTZd2jjN2Yq6G6BmoPeOnzBZmv0wSUEiLJa08zplJBl6rH
T+iE+9gh72yApvCGWjWeMWqiRNL/CdxmNUrserxn4GXkg3WqdBzeu8/y9NH+cR6x
je7g3Dj/lP7WkaLUL+LAcqhwWBmBvCa+pvzftRdtB8qECOLMHr93OqfoIA4NQ4+r
PpDryccHz/2FLKlVhAlZDqYat8mM6YqBwsvnmpPcx061IOrKt9hhqMFVsn5ldUav
GS1kALUXjlX1rRs55/UGsYqrcyYae1Co5tWWJsBVfxF70LcEdC7BYNqoOXWv371G
tU2xTM1HjRVvqzEOGU3kLo73b2V4288Hmeudho+f+E6aaY0OmrH7Oby/MgLzkUWo
WZ0jn0sUEfdLAR0XYHMEpgbdZXN6Vnv25FkoeOUz/r/cvYyNeuK2+gK0aAEjELFM
f6xAFO/jOK12v1kjoZENr7MN16tofATrGk0/tkJN9ARF0MGk4PpEq+nGhlVBn1iA
9T4o3EYsP+RJZRkQIw8rE/TEbaa6ZagZLH3CDJCaz0bCuB+SiNCJ+x78cgrPdFV7
nOwNV0I159t7X8PseIoCOHXxDcuQN8QMT2hbiboFMRxX4F6FBgyhSZuUh1ZmuziQ
8ukrlNv/MQpJSdQhbN8UYIarzJrrLHhxKoiXh2vJexOHu+bfTBZ2dBp1G7v7eSm1
q8PbCiyzCETRFZCpFcpoQDD+MeBAlg5MNpRaOM+B08lDFhtEfoonCgYHUi4i4a4j
WkkINLmzCZs8X6heQKzAWLYoaftkgeqj90MQ6omSBl+RCnb+DIb7tOuKeinRyXL+
Z6218pkrw1Kbuz5+FrY9meYrX3tXmH4Nt4/zsk/l0XLUE7WMLVe+kWlOiGqkS4nV
sKXEukeWwDboWalvgVj2ssxnp1seDd898QKnn/Lqa0LDpM6zWy6u+DYo9It8z8h3
C/95xeT46JVB06WHUksATXG1HeTFn47s16Ejtv9YAIoa/5DlZER4GcC1Y3JDCogk
zWuRRrHzoaN2EPI9cjkS8jKoY6Y1iP0vrawN9OAjIcywVzKE0T94zrXZ7/dJsdtZ
7fUuZQJQfT/ZpuQ6KKvrlSoza8olnHVRUMSAmH3YDNqImKjhG51t8WhJyVKookYI
l8jOKIR68mpBOfyJQ4h3xzkW6lGwO8au/JTjJ7Bz7Szf2DMHZRAY0UDqhfJpkIVS
j7G5KPeYEJq1T+We7v9mjEbKhRyyrGbAvH4HxtOqcxRPwYTg4/KXSs90cpmGg4uG
zTdqC0bkKLOn1Ytqi/Kgg6qVyLImkzREaUderMv5h4t0OqJUK3DfaHAPqMJjpK1+
Dk6hD1ZRoRjOP18+51Sgf56xdbjraidY0m6mb1pl8eFc/la0rzwjWSHHl1qjcQ++
wxFN5fEMK5p/u2pEQ9kEkETJnogi/2VBlP3JxyKVqlVqG/yCNLkJxGqKzW8XGZpg
e0H6za/qWYLLXMR0nHdymqpzKAeFT/4djHsx4oXIRIz6AWEGXidX+xNXdvpUvYPt
rMLhcsW6ChKxyH5GhCzgaGvwY2Sm0fHe8M+hZasDkI+vnvpvpHy0sOPLfSXbmqjc
pl/Zs6vBIEPgI9L0EofIrIBSgA0l7jtJjjK4KBErF4dbv68yTLAw9SDRiyK84mTL
1T7X7OTr7sfqGq/GTj4426khXE3JrUemUiE8yuo0ZSaBlDFhuzSVoVw3/DJmtaZ6
6m+amARYgSA57g7Hc6sacEvYlR3Um4qmGhsTFAvtspHmB5k3lfGCIYRsw5xDwz5g
40UkfrCdo9/e4ZPecmeQfSSAQ0J6KfzxIyIOf9jiyi/OjzuNjWLbu95j4UDh9NMu
gtvm/+aEolDziSu3bxxg/KjLHNcel+swTE8Seas3VacfbHCeg3teo3V4GiritZ7g
Y+UbU17i6TBPgDMzmbcmOI/kds615sK6WSxOTIUBBNJg5kyrU0EZGRdlNcsHOIrQ
tQAjCtR4krTGCE7PmfAlP1KWd/DmeOVsAq+xF1DRGJ16shRhfsBxAKqPt5INsnPF
VpjMtK3qwGPTxON0Dw7aVS9eIQgeFMMYdhO4d4snlC4J7nT2I6zQsqH280tish4d
olhcvZh+86BvjgYbvtM514qkufNZR8iLQnZo+5+iLxS0kDhheMkcKarbYyacOmuL
uN43O5LGWMdPtgBK+SBfKRYXyJVtocyPUtkxwg0zYLj5PqYZvCHB80q4Qhi8Fqq1
nQLKM+JY+O58rGInaiLHz4IGvWESaCb0/2OXgy2gUrtdJHOvY0yZAzHwZ9Cv8+je
JUxbU1n821rJbFcAtrV3zN0s8eDnJPxc7AWPyXL15HPk/0XZJi98GO8O/THz5zih
kDi3sOi4MjfvHMUq6J2iCUb775/xwWkzPgYNuLbK7Gf+tSfqDzz1MYwHHs/SNy6+
pk5H1KhxohX5v0ghXgDiCX/ZNyAM1ktdJO1B7BQ/oy+jsz+j7I+BQ5V4P00Q2ACB
bjMfQLGQwxMDDU8ZC96JtiJnwwdtW7bYTg85olazaHWdeqkaDh8PyAXgz3nv/T9D
S2JyoWuqT6j3f8HYPI8MGn6FUBpP3KC3bH5e+zj3uG1HYftAD+8nTLiEi9CbxEG4
+6sDVqJRyvh3Zpi6WlkkvNjYAmYGPQhCxEW20+FsQpQzBJXwJkT4H4PItRvxOcGH
6vqvlehdVP+IpaKjAm/2r5gt0q/is+FVfpm03htBQq2xvh1mt/ODlzDeGlj0ltdF
ZgIj2Fe5tcL5XKKHAgHK8SKMbc7yqQbLFG16bmSHjVdbsggOyD1mykGlxIOHlT50
plQ7wjFB269ProH8yWm1NsfPp9i1n6t3uukuHn5y6kvNrXSoWLINb4Cj79S7hTRi
to88xCCwPQZtdoXSI41nvh0sbbnkQsUaYGZmB5YRyGY6P3fYaIuxQZsWUDCzssCG
UajTH7bDbzeKlUnAk1bGIDwAMgckNAf3xl8jOhlCugzAP/bR4lIUFTrWuvACKJ3H
/j+RvWZ8+VYVeeDzK4tIEVdB4FGFDqtIDJt2HO6ZWSDiCITQjNQVYdDUFJpf4HXH
Xp5JJKPcv5rRKPf3WkUAvuUVi1u+6mqfjtLsCn9v5ZozCKxpFdWhkmdzz7Gpui0B
XIGG66wjJPJjNg945W9rG7KVxthzaf2lrJwEr8HQwdpEAWGBoM2VHkqgoEwG2PWh
yc1/gTlNfL9CfynhvGmb+w+R+SzShs7PpYiVz522P2NXW90aLpKtzukXbiHrI58o
PScQzHrAHQ/A+eq+GSGLYG2knxjnKnATBTZu0OeJHQjruDgcv5a6SJMwsD+c2fe0
zohGi2oVaTZm2xWxadOFclc+KUDcS8ZSJg1ZdkVNW11MlN0uIoWM7J87+Po9CsUA
cdO9DykPcgKgKlkeTa5QFH55kpihqJ/KsvSnaEjF3W/LL8wTMBbRt3pJ5zCaQAtT
gKi3Jn75rI5VMTRqay+LGsCLeDh40uy2f6L4tkKFbx5q4i/7FQCdrqjlHXZBiExm
/SCqOHyH/hirfqw9NvbiZKfKpMhpYE1WMhvuzrnmNcgTeabYe2NqF9qDww3djNmV
0HXwD0q51YopCE4r0JkdY7hf+w5KLgCJg8O0JveVPR46wkOiEHO7/BepNe76jj9M
vFv8NMEC+Gl3yanqsiwPNJ8FL8l7o0KH2bNk58tDUuGxBArkOuH/1g8atFYFUS6f
5gpWkW4y18tHsKq7dPogdNvkwG2fRBba4++KOVekYqUP6DF35F8wYjiIVdyw+oBR
QqlhmasGrJwdWVmczWj+eNDhd7x0j/zNlG1OPaQypPFHDZn6bi3yJP6QPQIs8hRW
rYm6h38souCXIvzD4CgfHwh1kHoRh5ZKu4LNuO8mslNYvt6ovk3chhsyODoSDnbq
PlzjLACcvBAEraCWZ4Sa8D5iUcVX8is73phLihuicuyFcy3iL6Q8AvoQ0UO1ajWb
G8NBZLhunMk8fgSsiv+3SS5igcBT/ijsmphFao+svcJcTX5Rb5CInoXehKDY+clV
dVLimz4GbS9GLO3eQQECaAD3XhPG8gr+ftTX3bHe2vgGge/i5/L9PNAeWkFY/UWF
H6cI3YvxKgK0Z4v1gyAvIIf+wHQ/UZgxcRBuPWHLNmncbN+6ShlkfMu17VBjcpO4
UtSkxn+4/2+3nMyHlUmJvkylZ+k2GeE8rASvcAxdn9uH++XPE32NHC1iTMh6EfFX
uYZ75gSwMb2TVVq22mIPgbVVo41Vv0bsldBBTZxeUYQ6d+WOceXPmemyRg2B6Zi3
H5HD1WB8b9HC0E7Z0cEpbG7kJtNzsLZyuqUjKd2iHjNK+oMrtdg9hxZQHnW2IC2I
S0/K2WRVfL0vh5zQzQFd4bkKZV8zkNiGq08Rw4m6KB0trvJNO9JIFQlDsFgh+VVQ
CSBftbczaf5vqTOnUHpQpKXITdsRJ56Gc/4glMzjxf3dz8EG7Zxvd+M4ieEwkMtY
g5Ik1zWiMbnnrr3mnw/YNts675QeFCHOwOP0OfFb69n9umdI/WubsH7fZWfbWAOw
VQw+hJiIuGHxNwZMNvZudPMFsxTQTksJ9YvzDonQmh7KWn3AraVs8wvZ9d4D94j0
6it1MrdtkQlIWjcrE1if/MI700jXNdtboBQO1Y2L18rl6S8gJiMFC8TZdxCAJAau
NbKZ9nISf848iBktvIJRdndU/5Hb6eNd5JR3YCmtWd71MgMgIKAKePUM2Jp7Cs31
evelKAM7N8CKwpDHp+fsJLpIPLgPnSO6mC1tIC2BGGnZXSpDVtOlX/tx5X7Ip5jN
WFNoRDRu2/rAFYUSxSMAaR/1WVmT/dgt7cGRW11gOS3QcN29jQPCLghhLk/L1K8N
UGLGtl8SBWzODkARRC9sc4knds0xqgQXza8cuKQ2Ez0o2eytYGup7re8TTb12Yho
OGw6cnBS0KpS4uMmJHrqm4FAarKWkBNu+vD9a4rlu5In1G9tn6nyUElhF4QmQsNZ
7hT4qkbLXfUmKcClyxkKjPU5FfFmHfoFKSJ6PDTx5Yid0uWigvEFWweN9cs56WC+
Tj2F6qtqX0w6nkVV3+yMpNpzc42BLetJ9cBrvXyWebE2qR1hj9xXaN1zCFVvyi11
zRCLkFEy+Cvtw6CnERWkcIuSog7mgQFzTjsJM0TY1Rw0S2X/JKh3hwHSn31W1lNR
mpCRdsSnOXiHpMb/3w36U4g7Exioh6aTKHwIYipBW2Qh9wKOTTe3j8c1cg8uwhBd
sooBhLZBgmbev/SfK/O+kkgkAop+ZD+OTsxuw5WTPY5GkTBEciTELnBzjh4pcs6k
LyqPNe4x71zivVpm7tl/csJnukQ4eI4DJLpOiJJdzqh1O8wcFV9riuC2zVyh27Vb
qjqGqpZJ0PXbg5X8++QF+SRP8Sim69XBaNVpyBb5m+LWXRcv/YQhHn1+jZhXuThZ
SKZ3phsxeZSezzXqXxcuK0gfhV0bpbYvvIzM3y6/YuRIBJS8OCdLmQ8nL2GQjXCS
aKtnwGiIXAZnMUYF2jENsUIu4kU/3VUK28BGyoXn8GbOKidBfrfnF4lXijswdn+1
W44Xtrml99wHXRCZx2K1dCo99vCzvPUcr2DLhUam/aFicMmSwuA4uGqf7NFW0nkp
8OfneZDP6H1W7H5vmQ9Qm245wbXUgLBUuVeoN6uG71ZE3QzANuUvmmHT7rleqa46
JYVtyNy1bfGdPF8sPbU2uehhyySLNSD8VtQs7s8gZdfXBG3Hg8hBM1SHrluiXECk
6oYc4/nKU0qx1E0DGn9TL2mwazSJh39F4xRxSgvBxmpIn3GZKVkgEo2lJRpBkw1k
7A3+K3pqzcpjOX34nJ+qgSWNSlEG96trX9Op8mZ6uR/LUjk8RCIKY2orxU2njWgx
pHHDA6KnxeRYt7NZJ+p7hMTKJRFxTZnpdFrC+4tjAk9sfzywHmXVIAOkGouBeE1s
6F/z274x3F7KltWNMlMtnXa1SOvMtIynfNg3R7+F5MrPP8NlIjhrFPfmcQ1S8Tx+
86Vv2zKk2CKC7eX7fqH/Vs56PH6+05FF55QvXdJy8ndoqiJCCeHZ0T96Y5IUtje7
iI8+ILCDm6ZP85QyhzlAA7ECzZiyszo17FFNYxLzOSzei7ltAIwu4gp2BaXSlV8l
bgM/t2ZdjH/adM1VyM0ygCk4u+oz7EoiN+ydCDj3y+z5eLTdqwaEvugwOYdzMifT
SHj8swovBptzD1QKH0zGsxlHZNqN4Pug67ty+7T0enEcbBShpZiyygpdFA9jYiU5
bSIusU+dUBzsLUCTutSA9Iel5ontaOR56NxyH9F+W4wPS5+RjYybD55Lsn51/Gv2
21FiEkYxZAaEIKMiKJw/9esYQFRXRjl6E2Mx79fb5Qz4hDDNNp9TDTGbA+K3YSxb
EvTK70QXz5rVi9V9iCgULI5T6yWm+WGRYNs9SYbFGB7m2kBc+ZkKDVg51BdUzL3H
2nJx4MWtd4igdkvGevJJyh+d971KU3tf6J5ey+eufBkzCq5/0Flmuvcl6fPJUjfZ
r42WYlFXs900CFAPEz1iiFJ2eJwZQM1O2C9+dbVxAcd4pgUPX2R7soSOoaqM+D9J
+nyFfsx7f+QUBU09C4KvlXqQLt/5O+nDk/4yAux9r2WN3YDSKNP/iuP8rAwHEOd4
T9WnK29V9zDwt4lcmj5WtP5KG6UwjgZmanCLj7MWDLJV2vm1E3mExx/WiSfKHYJp
hlcTukOO0Ueqcx3zZBXooi+keOCfJjrsbouTJNI0946xScnmUGSX2K9wzcs7NImB
I4Wfs0fsgUgNLboqcWZERP1HuhINiK0DW5NKCoWUsI7PxVNqiMDIA3OgWhTk51TK
KymS+p8xqrAVOyYqMYq/KB0GqB9JoALqBB/ApH5SEh88u9m14E8ABtM7Z2M90bXc
q5635MeA6e8JjiCASO1a6T9CRgmw2WNGY/eYj/Vx+qiOoK2KeeZtpBOmqOaXBRpQ
kNzipDoRodGPbV0x0a3RQvwNvciXs1xh0jtfo/5LqUkz2liOT0TRnqAXC+Ry5C8E
exOwiU9ZszyF3Sewcs60P1FAdVKJtX31q+9v95MMxDeT7XyKzFMxcoZPwHEcdqkn
qeT+lLA7RcLkd7LbdFQ5RVpEVYiF9Ba6KLFvzosxAhiXXl0HKRkGrwD06jc4n3TY
asrvXqsutLFMCUeUfYE7tmoeegYp1JMXDtVqgebtMBS+BumG5VxbxT0X+PeHiKkI
pZab5P0SMSqVgZLuzzSG9T0h1XrbR3pNR7fhVQekyBu8ufFWa4FTjXHvN9NSBZZ/
1wcFLUcWO9qPKQ7kZ4w9nvbiCrEBkSwgA7/6L0NwwYn2pW8h5UhNl29F+jVV4TV9
PkPqKtuGMTFORK8ijKrgKILnYBRT+OwV88+pnRJg9Un8xv9nhenlUfstWAr6NfTN
KgUlb25tqQ/zEWaCb58lSf3BwIEh2mLHH5CEtYsMTzkCjEOdI/JINPdpzhHlXgpN
yV4f5zsz2RkzfmTqQI1q4hauLN+6m+TEmpzevgEfyhvu6pWIp+vnVjpDjIgGpK64
uG5oorDxpoqmGvPrwMCRPwiakJUzAP325aUIw0+tFtUilGLuJwG4ngeWLRiOqtNt
YhHBIR+/2tsxkVU/16qBiiTmi0JXdIMMGXj8XVLfq7K1cVJdFyU1M9glZHs+6mvK
QJ0LPPgLlXLnQZ5jD2OXfDy5V05U24Ros7vHol/JCpHP3ZbIuLVeheg0sDhoDqJy
LTZeJ5o/5Vx9VNj1TPHV3V5OUA2dhMlGQaAE/c+433un39IM9surEumuECwxuYDE
lTZydvhtHqo2WPOpQlHOSnLsPxzY+yxxfSh0uNw65J0cTzV/XtnUt+Ds4eGIB6Xm
4kXEVQ4HK583/JYggdKQy2AyG7RO+5NuMZmWFkyDV5pzgnFVO5AXc5hhVqXIelwN
SFFGRCneOnmcwrZWSVosfwls90GSSk6rrvKRKlqoA5jxTLJpPGJvxE/6uVoXnykX
+vWQtsWZggIX8jSPJKmlbEQXpmV45J3T5v32yVAWc6VPYiuF/IyONNr47iuvxIjb
NKzCBfFHGt9h6E0YS1xr3OKO43vsThPLuRS02ASJ0Ttx7+IcCF10atIHgPqw4Elz
Vds097FZMMAWWcdbXXkthXa54eM3V16U3dA7yrZMNOCd4szJxSQaBLEMyt641oAG
jRy46fhpkDiAiG6eIyY9gw9uvpDikemDwuCT3KHhdDQhJgSEcJzdcK1UC2OrTnZX
A6aH8AG6kmutwelCziZezfe5MoUhbofxgOwW8oi7pj/+1B32MLA0mObp8jzx38IG
/MM6/4Lt7ZZ7Vckgi2rAQvW+CQfIMUNFLXHIvSe5rx7NObytw1dWo6wA+AsychqX
i8hYCT6YpBpsHk9Uyy0bj7NXvM0f2shBmwR4wZSUh1J5+c+WuvC/fAfqs3Udkouz
FpQlofPmMqt28JGK04PhRQsIJ89CFzbrIEyrpMbJn7QqPjJAE1DFpp5A6mQcHod5
DpsCDcJHOf3TxIYMHQr6B/CDCXfXRt1QiGB3kABFgzOefIghbP8E8Ij5u7h1lr7l
1ZaJ6HC1SZCjfxZiilNszyWmpI2zpyjkMf91rE/b0gi5ugbbsYd6qYBSbXBTbZzT
Oi1/3tEODgn0Yo3wTOvon5d6mSfJcuDSNKORsGAkFtXh7QXODlv3rX5y3oLKuS5I
liUo7UyV7Z9NvZypZ2kLETHEr77IVeru48Dw7JGBIjSC7173YR82gD8vZ5as7weh
1Z5i89B0ESMdUKgN0UX1fnqgK2xyh+on2pqLqWonBh27NantjpGJLOKpN7hOwGcz
NqHpjRGRqXVVeiPg+82hAAHxBGC7qj3oZWH/ceJeo5TQm/aH4oPteQhd+Jya2L4u
Q8VpmA2+4EUdYuyuxraJL4lGEaZyl4yLVNe566tAQY/2UmDcaUHw3z3A9vceCkAQ
PEbs6+SqkNiOWXBnd+CzYU0vNHtAz0nSQPgsjU19gDCmZuMLvQq7sYMJ07nEOKnP
FBlKCY3Jfks7MhmHqSWvqpl6sZ85FNu4T6A1xtm9DjhB8OUT9futaHB/qyuQ/11f
boxYg0WEBIln8SsadwVvbeh4IdC3cBqtN3kz661LDmV/n2hoMtD7ZGGM0C3lM9bX
xCt9/jp+DvB6C6yVnfzhXQL/+qDwZvfpoKCEe5mo4gMfnN+fHVZV9mGo4j7YwHer
JYQasIvSBh0MdBXadD6zneA86LZ9AlBv0Hk2fKl6ZzscLPrNh0KJyjp8umkCR+EH
fhZX/FCnlmXp8noOzhDsxvbN9XYfxYRr43nl7JxQKjQA2ftUBGgx5oOipyXZdr3t
dH8BtZ4HSptaNFX3PQKf+eJBlNthVa9qDAVPEq2VajlzkY3IXninL3mQELFn+9Vt
AqfreAUwQ9b2LGKhfWL7kh6UAe4+DHM58zhrxgpweEqb03gfaTWYC/q8i6NAB3QM
FqnIO6p3eelfkGf2Q9e5mP2wQWIVQRmOlFgCvaE/wbc1Reu2NKWWhjGh8n5E1RrA
0jsEi6855xgf7PcPP3pZQt7X2sTYH3rBzPXzpWTH7vhfcwkgC+XVZZ3o5mFIYb/6
3N6gVz1giAYPqUN7XWVkXbWAlJ95eusXA19BqRS03ePDWayF+HcC/rDIkL2wb2t0
24E53t7VI7ly2LySrYKRSuUPGW94GeZ65Ivf7T5vEscPQmylvJzpWzl4XJ2Spl46
E24Gxk47IkAVYqTsXuQS56o+Fev+0uL4oK6MmUqcOdrWpXq+2/AJp2bNWZfqx7VX
s/UH0IIhTkgi8Tzz23VJudvbT+okYAjs5a5X7Gnme43KW9Cdh43bYfKFQb01i2iT
yTqy9QOGmtQOw3+YRiGw4m1FWf4AGBNOR1SR8IuWTIPTZF1Po9VGC+XAh0lh3/nn
+8vbyQjdYV5lyy3rWxhsNYAVCzltSbsng9gzDb6x/l98+HMG7CKb7KKX0crzJnCj
fvEbhplqvGfRCtvneYhBUqDy/zJsuTUsL8ljibkQWoO3Wthgxi5X0adFhsI0iLML
Nu34ZNkZQhWJLH41PjNlJmyr00D+mzK2bLtFjPSnOWYoEcvThhFx9mwDTmqOcbft
P+B5rw5/dKQ/d/kND1thsf0PaCALSP3AAjXX4PG80m5WdLWAfOkkiUdXfBuxC+Bg
xE3I0IvjFHyV6E8j0A2eNpLt4z8Nt390hu4bfxuBUJVzy5+M2zGB60eIDaYubGlA
Emtrfe0HH1z8XkTfmrUBrW1tyC5UAhiQ3iaH2SBO9mMvzv6T6StmNrhugm6AF8UH
vNWyyiJZROMrG9b3lqNRjslQU/zXhMJaGBSoInGNPdQ4Nc5GgqU7Fg/BXXSkqPIm
Cw/6pVStNTQfTynUFHfEOwhn94Faq0ykztuD5hugZOGiKUbIAJHHOVAFoYGuGSpv
oBqXAejmzX0xNFd7JFpr+xlHjT8ojeqn25mQIMWuSu/+xB6Ifx30QN3WoewXwMah
di2Xu8hTEbYZGenpsk9bm7kkoCY4hGm871i+1GdEhwEYQ3MzSlW2BBpYoeCKn1mt
WvOpxx4WsLltFPi+wfz5XHeFqWxqRKj80vKjHLIwsc+A1U2JHh2kRNRPTSW7DVkX
JMuVgxR99vckAvVgSMJTQGwp1W3loVs4fxpj8csqJHAJwHqpVxYwIuy0MBQXHQJl
usdwjylwC3U7mOfyUnE0IIzvD5bczoZ587nrAm6cxGv7fMwhUAUBAN9Cvi1Mp1R5
CMOzqpsX/7cgcdorL37t0B4nN+puORjR29zeGq9eRCVKjDESsFFdk8Y7NFihSj4l
ScLtZgY2euuM/y2+Ar6Skn5P5c1ieQcZnKf4+oK5BuqCCBO78BxE6HVutgRUt7Z1
IFAU2FoFtF7x00+R8UWxW+nPrhOltoSZA7JQhxbPi4Hmazw+ndUx32C57UINn66A
KGvB4ziPHM8x9Y2R2oqqwpUM2OnJfMWwCxIEXCO4ej5wPsJ4rxDuB+YUgQFj/82k
dX8W/rSxKLK3x0JlpXrn+AxRUd9is8DwqT/pPCfd2z7+d7eLmTaA213rbNl/o8bf
nlcQBgdJgCexOycMWv3fA+CtZSZeEwvEs3628WLsOMbdWaMwpmgNwootG8n+HfDP
X5EGGKyTwolXuzHuKBJJGr1fpBMeG2AKPYnNPRK6L+OLWCWBgs51x6uGdBkbTt+z
fa3b6k2dl+Z6D/rMQizKOlJDrjtKdV7NFp53GZrruTcdi9/WBc2RPGHXpxw0KxPz
MBImme94MKKA+3WCefz1gVOG2FYMWzcNqj7p8frysQJNhyheO26BaapQ5PeEEHXZ
wE9NmTF0ObZsTg17HMOuGSkUoKM5tyOFH23cYkcv62eUCjxwIRIvbLu31eJjaMgK
cBvcfb3YoyaWnf09UCQri52hvBVDC/2pqNyS6tU0gwTbaKSPB6ISE6FytMTJRRly
1NfZoMgGgm1atrz5BN44qOYZ/kmBvXt+Mab3ubh4sYImHQhL9KsoekgfisKegHwV
yR9oMwABLHo0C+Br7pLfjTzn1fI2sVhzYKAWRLl2U/XrgS7DNB6c/ka6XDxlP9oa
iy6HylAMRMPXAivLLTMQ39pE/n48FQrrEDFPysYfglObbJPQRbwjoAZ879ab5THj
3EmhZ3339eiq3DE55UHVsnZiPArv72GuirLPGhPT0Cnzrn1x0amUG1eUPy1G99iL
hfE9IlEHTdZuwgaiJWK36lsUqO5woZK5Jy7MFE1GNzR3w1ZNiSgpa6dCWcdNZRIf
m23qPo8o9UB4DANjxpjkVr0XIyybf/GIolAck3/UGmViO4gRo/YK7J8Ijd5XmRyN
pXZXIHvIMOa/F0Uf5C4XvwGA9YFlrwrI9nnabwBcJZUGUmfDZ63ABAFpt7l4X3fC
1yyuxsDiJzTrBU617BMYRE1ZjRQ8I+dNI/RXRtSXixaAs6lTGxaVvWOQBHHtpGV6
WEoAKTk+q3XxSIjFaO0Prm36WsAhgpljF4vZy+8DBxkrDY31anzVtT0LTIctW2Ro
Rc9pAWECVy8Kw1+D/WmzndB249IkztWQ3AEpl9oWt4+fjp/9vSAiM4cAWEAyEDZt
hbpvBpo67Kdrq63SM2o5JGRuubR6Ldxv5zr36w/0fJ6fVBmiwYN603gk16XVePU8
JqnqoEDzCrh5/IYyLpkqDfcAL9F8yKFMx9jIWNU59HAWtwi/as16gYbEJkVZXG8l
ULtrz0vkx6QY5nKpDrByB1+NYrsIWvUhsVt6ZZw+bBP4fHPFZmzJIQqWivOWCDRr
FHRIWsx4gxfqjf2ziXBP0RnomTDdibJlALSWWdYVED3CVOp+Wg3PZaTLzpJQxXKQ
+1DdRKntpJZEldhohROXBf3aV65pWNsWADqGr+/Nu8GSdPl+6aXj+7cSr3HLwILi
6cF4FGe38TjNTWW6CPOGuaLqxkKe52u8dJoU04Z3ZP6n0io0wKt6JbrbDRcjhrXC
00ox+HNswkWdd5axJxDr8QCaBTBukL6f9oDEh/hB3tsvmuGsiDdAkx2jA85WHvx4
FWf/RUyuSxEVmCN1p7qrBIJjw6xw8jsOtyDyptbNEOUgjrcksDFGsKXSwrFv8lmc
HjLL/uyFU6xYmQHnZKrnim0bFkPrvzVzF7Hyw8G4leEzDjD8ghfIR9Mu2gJBm2Jt
rxV+LLvQAeMt7KIoMFlwKt/goHkvh3mE0hUxoVtjYlhPHOY9oydXpXhoEr3wIkH2
hLA3iyn75vrM263kM2GVN3kZlPp6w8iRSqzYs1/lNC/5m/m9LXqbpsbiQ4xVSoaM
rTYpGJVWUAzj0IhVqI+TuPVz7AONKgAKKyKX0ZUXriYaFJO5oOUdx4H1aceKl2cg
cmdFfLfCcBWGpqvaV0yxeeqs4H0OUBlvBxqpOSNB9fCDhtPcFYgAiseLJyqG8DxT
FWU2jhqcoOC4ZC7Xwd3CwvReGURzUdnDqxwB/5FXU648jub7NzsIGBR0InX49Fpp
9KsQ8XvT8yVWulNp9e/Yh9859nSnAsvmkVgV1otw/nthVWn5+RPbO7Cg+WypN/rf
8y1/veFsSjefNgZxuWW5Q5WAziTd7EyON7vl256rtuJIE3PRyeYbdwerCF3LMOEb
zORf/W2xNiuLBQRqDfqLn4551m6/qII7AkeLfq5LPYF/X7SFY7FiJZfWP+A6Jnjs
raTYmxTNrpFrcNTDLS96yOLA4pTKmFc15cOBO2zUa57XfV+/zdJZOInMnTfNKCZr
ZA9KRjNCnb5qlxi3JC9s1czLN17NUbZn1RCyKW/GfkpdRpMplsQz9gt+pJwPof7k
zgIiJ7stWrF4d/IGyQ2XZO+UxQ0gWt55WVfolu+ek+RdOLNlB86NqFTRRBFSnWpf
McpT/J7soE6evXZogG42XdDjCjLq3qWGkU/SGz24Ox4m46jeIGundfmlCJOv6ewM
xQFSom7QKU/xdeEqZ8T5O8CFp5nrm0R/4wc/EFIRz158t8c00672bt+DyTnnr1KV
ChsMoEk8hpLxdt5Q78yb6QKX1jSxzzB/THFr4oM7BxCUsIR57wMnTNbc7FnA/dCX
F0CKEH3QxyJn26fZrbQnZNvkCZAb0/lG+Youq0b6Eb1jWcf5cmH0dlwtPzkTR6nF
qnq2SuRbC8hcI+KKW0PJbcMwsjtgG6QPZ/1NlVJt6MjlanLMTqJWaPHtCWkxsMVO
vaufVsmGsDam0htIOmAdk0np1lqrU1NwAsiQ2R0saUMWi5Vj8GEueGYx6272cEEG
qvBQvWHd64jqTurw5rVHHVMqah2f7RWXFpDpiwknxJ0D18me3CjSdfLbmWn4RJJt
SZasfiKdVryMCWv1cfsR+otGhYa3AXzDKORpDFOsvCc7uZZAKom1iAtSeb5juRz2
VmWg7BO4KpPBaJRWGD883xqtZLonMYiBAL+eFkWywR1S2bexJHpXlJXsUSoRwj1C
7PBwU4Wa3nit/GGCE6/28raJxcheUISE4KS/vUXOY/YwxXwlJVfaPm6BgajZmaSq
VQTvZMop4cD7v7ODPe5lMerLpiq5bNIE1nfyrMGdvXjOxvF3YHL1Ici00I9x4Ysb
kLEgAXgvPPagUxeiJ6ol5phiwHKkq/r5ipyUxhEtu594pgKsNAn/Zm85t+ZzEU9p
7d53nfGDxdT376ZT9Qk6fqjTWPafmHVe7shlI8nnyZX6O1TGFFx1VLzO5qaEiNaB
Hw1o/JUMop4Q7Jg/wh1Xtw+0udYOlmJy7IvS3o9//DZqXieKaBqB6TfcpzGkCYOl
nQ7+Z/aVH/PXCRlTDD70wk+xu0GMz/CYbq6KHErku1avK93TdeybS+y10QX22Iv+
JIFl3zABVSjFe5usOMylSkYwVRP3WrTTV6keTizAfyNrrjPx9FjiDCBMFNjaRl2Y
i6wQ6guojYkqYiRAdj/48Y2dZ2NhzSDamcbTuRnJF3W8bR5r21r6sKxJXwBiSJKv
t6nN1kd6pCIjROgqkv5C7RsQs478nK48hzmn83y9rgeAhanHcJFMFMq/x/x90+Nr
sDol6DFTQu+tGP1UGYSHcAgkbVzNgOoorUg6nvtuMRimvirkSFGxFhVisnHiTqQl
fD9+HtRr40JWXBhYgKaWnzmZ/HabNeoJK0e7dBcj0l3I+4A/s1jK//eOxAFl59sb
mqugaWjL1rMD0MFdEJovqW0hqDHim32fP4/QnJvlnsE8Tav3lM5j6WqBj2xACoRd
vj4QCw/fj+d12adFly17d/4UlvnwYAzH5ylrc1Yyr8ryU4haR+oWGjJg5ayt+8C4
xkjF/OwQLQp2nwtQxszbHhsDSgfDdQ6XIt1v2DYG51oVeJu5DIB+TcW3f7LmBVIi
sXoKjDCqQMO1rpIWvGuae9VUAdi9O5zhJYeyp6eBUJlhyCMi2L4TztX1EXUBprrk
CteXHaD1lY0uS6nN6/leEJV7EJKdCzRO1nhq8mitwyRg5U0Ws53GjHwvMrVIRfnu
N7hT8h7tLzMrff87R5sSJYc/pS0P5YM7+/vAngIIxT9QWL2daYWoEJhuq+41oR8Q
hAnxnQ4W7heXq4yFnGqGzGA+Y6kpgVlYwag+haV6X+/2bhQ+1CE9DKpu574P1K1b
VItjXZ+O8/oYfFSmQ+0qgGA9KzFESq0JPCOb6QXxISg+dfOspAOUtRcMvNbsa5GN
3C25/MJPtfYD4q1QF0GmlrjS3WdNAnJUh734KNT8aUVLXCkW7/4N+0OQkhkscAZp
qia5zh/pzBSEeBY274jmvFv7d5gcq1XXhYFyw7mE/CgKR9Dj6mHIQ0cEcO0hLCkY
5Uyy3eunerfB325LwooqfUJdRJGFV3Gtfi6ddVHeGoakdCNJNjGtAX8jvNsvHm7Q
Apx5f51WSZo7pRFIh5ORvWuU3oKLFvPZa/juL8mo68Lr/+E+YcDj0hhf477Mrl/W
rl8xytRD313eucCu6/bq6DGWWuiMcXkLxU2ro+xJvfahcXdxWenmzEwhllEoYiyK
3aKtN4N6Ry0/G4i6OC31r6JtJGDEZcTnv+Q9Xb3P9fUCIvTjKW5+ReVFnEOLc7Sr
mHsj6jbV3HCR3QNQKZ8CJARg5Mzz2Pr8PR/z9h2ySeSz6XdfgeLfntdkkpV2XW07
JxxvwBScaQ3puX5b/gVZLbHXOFOQNDqLWEx7jKz0loZqxLojPLqZKptBN3tKXL5z
dzfyL5h4qVb+AlOOBV1pVr467v3y6cwY80MMEkotpUiwJxcIiiM+t9BXGZAJuht5
YyjFBIbk+dummsm4+/Prx7+YZ6Qe2/4HsYA6+w8vfcvEuKiEdgvxLtocs2F9k1Be
jGVb/YwwDXFJVUAxGUnGcOhq9FY+WwOdk7bvaMB3yYjPNfUcgnquHg31/b3GBgCY
xKZ4/9wL1ipjL27Sab1GmDkMMgKmPfhdJ4SekYEb4b40oDid3uB1o4BPYbivVKph
Z6bJTGPFf21Ohnl1mXAFchaSM8IRHnc29M7PooJ+NXi6jo4aVeXDfUlEX93NBrxY
44qYs9oQ+g2ozynUmSClxuSfa0IzeTsuC05Q9zt5x7sIgyiQ+yoI8D7K3oT1utEf
ctCGLV3MdZfXvVso6FypBlfAXiLEgQMGtHQJ4/iHSXSLsO6QOSy0WfVubUOpOGTP
Zc8mLK10x+vIh8MnwRlkARKeJwadhMvR7ZSZWAh+JNakD9ae+nXSMqbc6jVjl3tE
TNAxIuXA3pBAbLFvqPU5Hn72YZpH9UPeSJHY1uWmLNWJjpG6FAEbhJ+WXPKeHZWt
p0wXRHzbhwDHHzAZkMvtq0mZlE4eHsd/QG2XzDDVqpIuCrcipclW8gmXgjY412ZV
wMAjfIHJKfPZRs2/H9zd4zqWWk0oZ6JLxyMUbM1KfM51AoVCriRPQ3Cl0CM535Qt
wuDqvIZ+yJtoyLRpIQUUszBUh1T7Av55nTB5rpBKwVLRK+5mzHrf4rR/DclXWtC0
ZKp/BQRYk8XeJtdGpJ4HplUIqK8psXgbll5eDZAN6IdVcvzQlRbfIjeoWZZzLraW
Acrmt/YwnZzp9SLQPrDFFAqYhnO27gmSTBHPZhbG2LHzc73xb5Wwerjum5KJQqyK
9kTmrXQeP8aWJsWS8EWL45b+ZEfM1W6PZc/sh7lhYRxXAVDZ/2H2cTUo5a7RX5j7
qIikXvvsuFzbWnNqYev6l4P94OLXu8C2IoFbPmk4NcKW6Og6ENJicNn38V4gEo1k
dz5j6VOLRSDg5M0TTE4574gvd0xahCpsVdR/MgNqJnXk572LvcfJ1WoMccu49FtA
K6NQ56YIQu++YT14Uh3pE5Hx11xMnxsNhLkIWGdcrlPm0E58WCaonYWrnhmcu2/j
Ieqn/lFvkmEYMWpVMRxzPMqVKyFSb6w0D4kkWcivGdTAX9VNMSGlyJDMGpqzfv48
TKKeusns6Ntg6IbOZFOiEeKTbhTJiAx2gb3gwtBrBPfAQ2dHLV+luX+TfZDHhYzl
ccMEq24ZSjdrXzWi/TTfFxi3VbsS+JSMJP6GgEVCbOoLvqzw+fhAd+FlkNTDKdTh
cODV4f520jvenN1JmEzVvFiTkyolKQg/qcHVQjOJVo5SoTFWeN9gXFQ4Bhg9tDxg
mimqn4GvqEALwqIIZqD8q17yHliKoy+NPuO9Wz9wO7LsZiGgi1RoLJRF5roCoTwk
951Gi/ZIXFkhsf7Ht9RJEXyfYpO6ZSsnfEqem7AQAWVaY1JpSJfP2X/A0EXKiFNC
f02w4KByb63iEWj+4JbkYB2GcmaFV1weKhLYUzwhlc4nK2OSFDtb8zL7awyIuKEN
G7BrkQnEuFvNtkn8qSHfxe2SEep0KQV5VChFd6fvoMJ0A1ds7hZmbx7xuHajQ26D
T6G9EFMwys1IdZNQltgJwdoVONxvSvzQfIw4MwIp0c1xdlooTyxk1fxTNSOrqyW8
EAqBTXAxcHsqUoNCePvJ/EJgDlr9Va3+XLsbifTxs+M3TolvjvOSQVZXcfVTah7e
ft1mk3942hcJkeP/6UJF8due7M6DAH1km0No1I2fZUevjp3X+S38T9I0ao4uCDHE
B14hRaZEMN0WmU62xhHF15oDAYCKreH0tGzU5ipNDcVU/i0pFTjxoUdgrWiiOfxk
LLe4MkunQVnL6kPve/IwYaXQIQPugA4zxIU2KSqm4qgkiMAQKnMj3izuXjA+NbDc
FRYKbtbAIKZhBoRNbVmbsF+YqSoS4NJn2haeRiOHkaYa05gvqU7LNH3uHsWGThPH
k+967EYy/3QKFRN/RMmYzPmkE04HxFfNcQ3xTHDkucM+ayzKtGz5L3b6yzttXWxA
gadLxaE1rS/6H+EqJ2qkKLVQtK+hKn151awl9+f9EOfYcrCI/Em682YDbC0aBKAP
dQ4q7yjAi0qsfKjntP0SSJBYtqY1RLaXl3D2qxr4/sv2csa3oaRBnAgYN4pjE1A5
ZnBN/GMP5g/YIxJljGAuTEEAF8aQRta87q5VobWXYf9QGk1F9WdjfZlSx6mwASu1
qKFiOC2OXPH5QdLA64Ap+8LbF0yjysu55pS31n7aOk3cctGjIqMgwNyj3txx0WgJ
JipR2KlfchEcRpR4ZDMtlWWmeGU8PKXZk/8jZbePwVmlf0wAWo/tr7ypyHxzoq+I
8FpAL4Yd9QGdgHkR3Fq3pF6gDqI8e3yPRNo6PaCmAtFHppQJsBaFlKJ+Jaf9qiC8
zez8+1drw+VOLvpzP3IoBK3PSnj/LtGX6/deuVSXdeTvINT08NL2eaNbjLhknV8C
oXhQdnp2JwdqYcO6Y206IpQKGmIAcrDqGX5oQYE8yZXgLZreuJbjayTWX/3zCRHZ
woDln3NFszsFqRacnyWzZ3vPPM1c5Cy1pYISD3vdst9l/wgYRkh/zgsujowLYWMZ
XQW7Yf9EgavKhP2VN9H6zE6XI6RfPMTr/S9AIZF2xmIWdUOHIaDCAnRnAxIc4TCe
IrNdFLzQGEX3oHlME81Tw3ipCUJWvesO5M8pqSVJWZmirPRQEyixZbNyefYXwCkI
obHl5IAooC0u0tFqhkcXYkMV+Awpt1o9JeH1Br8eiJd7DB4LP3AeJEJvFdioGZTI
Ioju/OretM2Vf/4GOs5KMKkQZ2ItyJAbIfnFTMr/yZenqAXTnavKJvwnKKSr+HgR
o5OuCISldq/43ynbaCMMktY09l70YonZ6myzqA8HbXCnGX/aCiex5/SFGY7dmmKE
1ISqyfoTN57m01Kxw9lfmfUTAzQsVGhNj+I33GYk3pB8Bmb/9qbEo/WKiZ74nMAK
/BZLgtIzcv48Ut0Iklg/3hAvljqBfWLOJhVXnJIOugeBPOo3Sdui/f6Wkzt3YcYR
OjDYPkYJi+tYpnn/+rAJFHCknklQpGmIz8/6Sexue00+45Dac086J57ZmMk/e8i4
B9jphMGlPdFw8Ec7NdKeEhw2ROoQUV2+oB9Wr+3npEFFzUCGKY4czP4Usy3n86sA
3BM/mWQ7wVa1J9xWqB3Ijcu2VVh/LRb41Ad823MmUnU+iie0hizgoSQV+o4PCL/r
fIwM3+2UwQfjSMPqzOWX0dahcxtD1Amswzp3J2F0QgTeV9Qrvj9v1g6vMIsk01Mr
+SWrfxS1ptQ4fknZcbs1uSHYnA8mj+X+dOkLO+ij1WDh3gKTBmdyeAFFlS5Pfjmt
vXPj3L6z7DTzDBrotrjLSybxNr7qfIcuSFverndKAMqvQ9CxDUsO1OzpxkqOLrQs
sEy0dtosnRd4Hmh/i2bDjuWLgJFnkUGlBJGa55KH162hGcgjnwlh1TDRWbkf6czH
psV4FlgSx0hxvRoU5VcowiRjPOJxmhNRm50kC7rQ1XcvJkin/LgujZ0x7qHb1r4J
/4+qEQh8AO9e2TQ4VLQbgrIVgOms9eP2yciNAXj3JacMxrXcNi3Hut3I/lCCAevB
GqgKqcclU91MahlxE67z5O+heV0n77/KlJ8wCb4FAOH6sCqxm3tj4MxRyKX/mF8E
tbeztr34vI3xWEnbxJtJPEfNSpKaC12aBfip77Kg4r69W60oeyMPIuv/f6xWa+JY
FuRkjSmE9JCTrQ4iEpelm+a4FqUr/IZv/ve5zOs/bSLEljkXbEXlJAl2p5Cbh0PZ
G4TSfMPQS68bTIjl19oYf3g+A+06wBRf3jA24+GrXT2rsuWRjfVhxG/8BVXcZFQU
rwnVLcNnJDhyWtNABGZWhOLrMTTrePkhNirLnB5s9xrWZsjeZW6+gbRw2r88Yh3/
pxgt+rvjzo/vCFM2filyA2fd5xjRzPzbKRDX4yjLywz1ZPsBnSzod62TnoobDTyp
2U90Yni+MYnJVtEwAib1osGMB8fly7xE7oI8elC5jugaP+vmHwrNMw8UpjHmEzgj
3K3LtcEldN6bTSu7t7330bMbf4r3IoZ9QCcoXtXYo/M9CepClRYC8xljYvKcrmAa
kq18GPgPn33waKUyN0G+KEPVYShd7P5+xGFZ1WQd1+95xGcPhYkmtcSEOEaA+oks
ykaM7rN9zhfhzvGT/9epJyb3EInmqWXcuWfkmqBNHVqonrBxZ09A9rNw7TYDlkBc
rvoi/bMOVROO0FzwrJb2a2EPbE6BaW7PdmLa/J4cdLZiqA5EGeUm1DxEolTbVE19
+faM6OdiI/SPo70v96ohfH32nh4GGOWhNU7lgQt3jZeUR+frXxec+vnk54gGKKMd
vjfPYPCMNIeHj0Mlr6r9OSGcuqcoLMDUE6qKQdiQ7bbXm+4uUMW1LEKpsmCrxUPi
Bd/GbK/pIzU/OyQ8/LO5fXdf8xS/EyuBJpaD04Udb1bzfabT3DYedk19i3AIjY+E
SL4c9le+TiPIrpJ1a5dpkScZP3rptLmL+wdaoY3Yvb6WfsIP7DW5S97Y3UWoR9gy
VwcYzIGoUkDy7p//IND7unH19U49zZmzrM6tGMJCvyEt+LDxAkK0dv6QpX2j59EF
UgJ7rEvXMYlLueU9vxsdlTaHBHD+2lkilcrvF7j++qW7YIUNKHbDfBVajSOcTD9H
/yuCw1VVraXe+9MVreP8YIjXNVI7fx8/ltaZI7bUeBDx8cbrCOG+IRi7OGCvdDGI
oIg3F98NZQNRooX/gDPOFYuXY6FED1DSXb4DlROXC1Pjdt/jltrt6uyyYaKvF8Ah
bsYd9fIW1V1+q4dcjQo65VisrJBjnmAQQwcfPk2G40TSrlIQG+c7XfHIay2m0L/Y
bpPBoRlXIcpvj3ze54BEWEDA8mm3Gb4P84pNea1ELLY9xcXxX2X+iRE7lyGo+by9
rlgJPFLlEUrygWglQIlhkSYf2VEhCLKMekVE06XSaLGJA5DZmUbM4isJ9V9R9vEV
JO5BwJN5r2o+rZLef64EM5cB5S+6QagNUKGWSedIgviEF3bw7I/gsYZt9lvl4Xe0
ZqiiReB5QRU09sDxe8gD8PBDmWP5GlZnWmW6UL4mIBO7zPxsd5Pz1dXNA4bdl3BF
3RtSCvjtHdPU98/aH5JrhN0yODXhayfFGvZnyIHXSb2OApntmJM+mAgYknoeeYvc
HmDUauQTMdNPysb6s4cPVJbZzL5xRW6V9JAu/V+3QHD7Bz4RGfcfk6QTxiTmz+11
YciRS5+lH8EAw368Wan1I5XMFWtz74S4zxHEjxuhfvQxIbth2W34YVDM43rYfLCh
l3a5iR1PapTK3wtMHb/vB4hq33pJiDQ2Dn+Qgdbanm/NusaFJ04p/JM4932PIiwi
dAbK8iBhTZavWEJVRfNpA5FbSgG+iIZF3ZzTNaCbO/kp9GF2zUjDl2Zi4Tx5qvJF
OpEq43nXwhiL8iIYXCdWYK+3CeqYeCq3mQIKzhtuUgPxxxLbKeMTnkgd72SLoszg
ff7Pk0LK0zYycw8ZG3IWRPUeSVEj+VDlK24Yt2hE9eCiRmWvyFQv3/t6Q+7UPgaA
1THeJQTJCF+Gpy6N9pQzn+ab7y33sGdvfKnFUG1hs0sUKped2TzX4eawZX0OHBdG
yJJARSJameM1mFfkBh2etoANQ3twccmSP3rAQpt9knFlsICpGrchadIdLIHX4nWi
tmts5ZjX9PBsjtmyhZX5jNAXTFISBRnq9wADgy7ZQiXZKH5PfE0rJ8b+7w+dTAgx
o7Hl96KRHVz7gMQuFh7WUk/Zliq8h/RvNG/PSPIcXCj0J+KXJIyFDpk1FyYkRa0T
yeVtKcRau+c9G0h1gJtqXgW0XDl1l0Tn0cOC05qksIY4mp9yDwhsLa1/cM6r556n
nSUHuDo0jfy1lZ2vLKGsJVJlmbD9+/nKeZqeUbGnTIx+4icJ5HCCFwvSad+j3sc0
z058oBwRPy/XraGUvD6w4zuaUy8Z2o9uXNEzg/3kEnR5KD4DwkHvN2auUOVgxKey
TFjPlehro3T8mQ6C0mLqxuwMsRC4vS7qqnxKyYoMA8V+mBzRZGPPecS9x3e0u4Tg
njr7tcqTZn08AmE4Al3MhqfRMlEjhip9fBtqnAqdr7Qqp0375N1dkM2QHLbD1qlq
U0W3uhRpqS66Z7WOu6ZJSfIHK8KJakJhwvHlAVbihP7SZzTBC9DKv/Bx8A4Seenl
+2tzMH2tWJ01DSexmakr21uozfF2+aNlyRV6npe9rhL84m+aDc3vVb7e90WCxxV1
opD0L5UA9C+ZuthnnhxQ/0rf2pX5r7Q+RZBNVvoCoMFeSCtbHAjTP6cKAMYcGRI4
jWXGQa+vJjsHofb9ZzH0YLN2NIIdbtspSU0cjeP0Pxla2Ypudf69aOF/jZkCni46
T3StbLpZBKZJD7pS65WoD1Ogo+HmGwKqdBYrvq44sH8TQ9jOD9F/naCWOvzhyxrd
YKcAPt359HgRI2q3W7KXxgoVGj1PYmE9odRsLS6uNSv5m5pqzDFWzol9kgy/LlKL
F+5BjMvFQBJ+4IX2vGjSK+jAEsAIQqomMKCmx4q2Bz6Z0xpzMC2XcIgubHG0zBZd
UViAygG4I7b15dEXs41AvvnkyVyv1frVob218+/afl3FWiptR1SuUQOjOvBcq2BK
UqFltxm+wOLzNDAGgm9+9zbEJ2NOlFDOeT+8x0lc2O3FLVhFIwXdVLF0O89/Z7mL
6VvssBVHY7qsHyoHJR2zw784eF3RccN+IOLyh/drfLPwKn9i+hnKzzuAziSeGzGi
w02b59U5p+ns1hnfVQcKZ+QjoS74PZ9ajVMueDC8LF8cvEyPSP4gAT/uNlsTWt9h
JuYuO/DO6Jb8g5oio3sqOQ4m6X+vLav3vFNz9J81iZWYgSmhgLN8BdgyMUXsqVwr
GcJwScjO45HLR+kALNbArLVDIrcf9DytpswqS7aa+Ok6uuoMf3LcaFf9zYaRGuks
PTws2moS3F1YIF2ZtzbJoL5G2G1m9aVjUoyykwo3GtLX9SrBqvCe+BOsWdgh2udr
+HPUI0Q4hLKzRuraaEg7gQLUo8M9kbuDHVxyO3wS1HQ0pImABpbJnqWgIrDi5x1x
KHcUXRwGG3pFyEwFrJHwIhnO7WjmAs8k3hqvOEg/Xt39BVJX1VTC5/GdBLT3NU6x
MY0F4PtzybFWpzGfsKlbUSI4YWxKpot4ephmaBnlQqLGrinlEOLMR3Omep8e3+Yv
j+PNDs9JU/3y70ZCMADAIyi8u/6iE+8iqlHOJpv25vsaOBJ0aE5DtBHhynHE5gms
XtwWYtov/fd+2PC2re+rBr8W1SQCmUtYYQz9lHjotuzRUWin2bLo2M7wcZS8C0b2
oK/ih32OdxJL+rSBDOF9u0l92crqR47dMm+8zJ4R61pbCGbTj4yolwR4Csn1hmDm
kcBKxoQ841K5Bw+Vx5WsETrKi+PHp8Ql5qXg8fh71MyfywSTObGGdsawM5cVsvNy
uHdaNaVpysy+cYuuKuQPmxk10VTdupjVnsu+mV1e15riaWwYk5XOqefI3jssfQwu
+eVkQPeDrdSKeNJaXDLn5nhNIc+4IrDt6l5QaISxgTX4trkgXRbesfuef9QZGXJ2
InR6CMRPVa+SB8vmuwKuvm9E7XFMea7fEmAcoFtow4rXx52GNXq6lN7XQ6dAtZZS
0RqtOOkB9uWpxwKkjejtb2HahjdKelFeM1rUmlT1kembddc9GXbm0RmyjfZrIyzc
W+HMK7kPo3mG/cBb/C4dm/jKGlwUhUZ1WlTKDVrsaDCU4NNjrLaO9zGAFMP7uTJk
mAx2jWza9LQuyttl72I8RStzEMDMmdcuCp8zSDm0CVr27rrbQYy8RP+AQa+S3lh2
ZwAuKx+i1aer/vZVryz5sUwuNYMTJBAuOABvbN68t4q7oh8E4y1bEu/6bRqdpXjD
/O3T0l9fo8fejR6PedtS644N3GrUFAHRuLaDpa4TAGz2lm/1N+ROJoH8YMXv7SEX
pbwChzHuOLVZp0a8dSFkHkvo9VB1+Zz0JMiYBTukFVc9miBLXFF0qgcJejnui5tW
k4Zje1eLkcXzGS0J5DXG6tiDeecnIYpM7ozezyuz08nEYJ0y0rpXnmSsF8cbZHhn
iyR/9iZy/Qk43jNbubRQvgoYKDG4ovEFQIZCo250xs6D1If3kwCfoEo22+ZzmEy1
6brDpbmmvm267M67jRvh+7C+u0xDl2v9SGCq/StioNBC0zQZT4pzloFZESIgEOCN
PMQd8rqKmoqrhyI5kMcVsG8ABZhYF2p/GDp3phUET2rYCCmhVH0krr0LCBMX0vIa
EOepKHN/KkLz9uMjZoY2MtUoBNTurzI5BRL6fIbJOtJJj+SMfpEFoIh5VpVsqjtZ
CcoaERo4bbtvg4aAXzyNYIqN7FQPNaqv7clwcLmvxCtOIhxLK5QhX3Y75DuNPJJT
znU0eZm1RyiHpx5gEB628Z/2vikcrdsxkxtug7J1A4hGEUwvIbwSvWCaRCwNZ/cd
ikBlLR+KVz/f1wbl7R3PKtqmRilwQouWZnnn8hz1EKfuvDR2h4ZGvA2OWVtEvLFC
HyjW6QFhijpP7J+VcHFKtF+VT1GEiVcZGd/EtYJppZLOZVru9ozg0dKpnxG/kRVw
uheugpaNKj5X8IZZ8JDALlXp+ts3zdTPKB5o1RM0dOlJtmuZ8z99MVN7884tY71w
9lHY+6bYb1OVxPUQxccETq54PX10kS6vCyYo+QKZxTwSS+Q4DucTxYKa8oZ0AU6W
k2Fyq2xNb7f4T6zhJFIkU6WUCgL32BCRSt3lKK/x/0bAbmRrK6HtyNOM3tFkkCx3
tgrTMc2DCQnjeAY9nCiJBeSzOYYbUniOivH8e7aog4UMghmciALCrvcu6Jz37KB7
zFPCngYQRpUREWrNzlJK3AS6WLa8kHNG/vu293V40i84hba26MBqJYIXNS5V6AYa
r5mKLQd2Ms2y+zEjrjRHO8ncgNTqN4b21EhLW96skQNQymjNHp0QG+IH0OFxOrDj
TilqD5u1TXnHOETDNXB0yVagy7WPYOBFIO7EszwPKiT0Z7zjKSo5nvtC6U6bxSlW
6yxenBCDyRhYQQE8Htjr2x8OsblLKzYK2XfxYI1fJD5NXWAC9MZyXdqW4P10yeeD
zPynOZkBp0Cl6xl1Ia8LKu6ynugNf4MbspShkZO17ZVC3SgAvwDcrvadLumcl8Oc
y2WsTTk5NGWKzmLApC4YLsOkgMCjNEoYaQ1XnBKZ+b+InobCpGonbGkRjmYC2NUH
meQm68uiX2lwP3x2wto/nO6EqP53AOtOnLPs99cw2r+zcJz4pQ6omMa4UtHbBfok
Z/+hP0kYsqQ90gEmCHw3u4xduCg5rJXbez0lrbDy2S/y1u0IGNfXKXU2kHqDL06y
fmXZ3YXXSfXtB86ZQHLusU+2IL26qz6JgKahSe0y44PQeyqKczJM73op5SEmI1Lo
3zxZR3qmWp19eAoRvrA1KqYh2YibEVbDqPPRbV/MWgvGTHvcDvkIBmcZC8Ivfg5x
qZfVO3ZpcYik/g8GU4uo2cEuhPVA90KgK5ahgDMXCV+Uc7jm6vdHBvVsBIm54oR1
7jQWEslRoz7H5mRKWqyQcw2VWqfOqMvE/hj2C0fkhHG93lspc6drnkeVDnMc+SSP
3yqDhtpOYlZpPgqrxn+R1ke90iPTcZSPAnj9dP66RDECvfiuNtxd0qOZNbGNdbN6
gwq5q7lgR57FN1uyrdHdLMQ0X6WUi7rmMQ6mkwPWPT5SKBDC80SyluKLsDCkhGNA
f6ZBVg8/8mzo2SXk+4LImA+OD26/SiF9i/ildxlY/6LgdkHD9HK481Zh62fWG+kh
Sl9bbMsvdV+oXLo8ILzMAdWGKVjINVR2gq/tNiWKFGuarDB+gxPnsWbLxwH3FTrP
LsF8xlEIvm+eC1u6hmkeDoWkG7myWh2r4ZdZqrEaKYqBawD+8NUFTtkNBK9h21D2
NcvNjeyc05F7InxrhtwgLlZXvuoqZn0187ffnuwZhDCfV4mZravbnkaVQIRWeh3+
P8iwYAW68li94te5Hy6g3I5IU6WpL2viql48eKUC6cEDIjno4Ao7nCi/JEeVGd7L
qlLl767qyBV6oQgiSDOKD9k1WIYXEZnkINQSgpKYRzFKOwlq35TrpJVcU6917l60
2j7TeLWWqum89VT+YNZCBCYwPeQjY+lTO3C2vLPdnQFAt6J5aT2IELg6XAhBkTtO
8HJxVMqiTq6Ls7SsyEOekvq8yobPOPWHS2hPLbTTu8KSHcsKeSA0Ar93QHO25qji
jx6L8zpFnIo9Rhk2THR/EkYnITcuQEbClT0rweIsYF7YfpyVEayVIQ/TmyZpu4jH
U3m2cS++q/RSlM77skN0vV1GVCaJIuJ9UkkKUepNAB+fUDaDQWF+JcMTHFjvjTiX
coSRTHbqwkZchtoEMpwU8iqkE7dWLQY45gzpBSTWC/D/nh9C3T8blsBfRSpiaDhe
ytPE3KI3xjTczmi7NDsQ0yupPICWeIFAo63iZ9slhIt2XkeqO9KL+iIFsBcg0QNW
7/Tc7/XWXfSs2Bd7X48hgpHR3Yehj+4k7BnHDQ79f/xaXDp9lBRJkKrZmjWr4kR3
vgI09hm1mWwqO9xe7YzHzyy2SSvR2am+0Frh7UHnY92npli3jn6yvNu7+Ybo2AlA
3NBqsCrf71P/56qQPu6FEP4jd8JYN0E9bzhM+QpE7t4YsT1DcUswi3wkqhJuxlfF
FCn54uM4qj7/iEb4bETUuYaGhg5EVm0jL6Su/kDqgbUvZo1oJrGFH5DBeiEnD0fj
YvH21UMbLZwnb948fpgO8Hjyg/yqUzEOxNLRwtEzLyhTac+c60v56L+IXNRNNd8C
CK4FzF90f7L+HukWRDRCoq6j4To5lT4shWwn6qH6pcivf3xXr5cdLNV4ghv3uoL1
e8FXgpOWkG9fsZLib2yuq1c7pmT9FMmE2tPAIDoMALl7TDD+tTS0KBZ9Vi7/qQvf
djMzUThjRzokRRevCdcRAhjILRnR32E3fjAtgS3CsHuXH5sE6GPwAd9iVodJSOod
Yxjn6gX5iYx4nCz7j1MMmUhoc1L69d8B8tp87yUz8NTCifvNYs6k7gpBQdAi+ocn
i/9s03jaOEkNWbd9Rncfg+0F2en5Qd2MKf4aaUo0PBjIqiv1+IWhQ15NKCkinzb/
viD8+InoA78tE+TzfjgISO7Yx+cUOr1DM5re3J+1NPQHEAQPayTDJdKK2UpojHRs
FicRdtb5r7sZpcz5RTS9bbnAc+U+YtLB+ILi2jxkXdU5QYNqpRg49z+mzrJJsmlX
UVNYslEjSGmAYG5jD4e0Beg/CDw81tyjZkf500w5ydOO/QtmuarOFvoqpv+bo9kH
OaEZ9nMsZapAJBchlhsfzTZPtzMa7loCqOICdRrt0FX93DTAQVq2PLSOMBT0XWSB
pioSNnRsj7ZDPg+nAFmXeswTcRGHddKQY/sXNmUVXRE+rh6Hhc2KeCLLe2clEycB
7NK/ux8QB+iKI6Bn1ddOjyrmQbLYa3TLmU3nqjY9wKrZSFmX6X8jEhchqHD59FXK
DKmDBfDYoVAOS+9qG0c07cpfYhBNomAShOLSmQHEnGx7fPwaYe6DR7oL7+P/GY09
qESftZxMj/hNu4nMc3hFRyhv+WODbfqRS2eg6jZK226DgCg0e1Thq96l4Tka2EZR
6YtAyQLIKdjUhhnFQsStIQlW4A0B0dz7E5WSJRV7wBx8bjjmF4CrepACyzyTXJKB
M+c2td1WQO+MyH7/tCGyj6I3vHv9St3tKNWM6KiUhtIrCSSBXalFgS4VTlqjsLGG
uJ1otKbw6sLLEeXNMySQMlcFYY2XoxLuR+nP66k5NEObN3p6tbJLwXrxh8HRnmEL
vIxP5d8B6gYO4wDijZuvKBnA2S6eLeso16J5H8FHnN5ICCAYkHOnz4usm4h2MU/j
nkaz07zJLzo7rU37IzCTC/MgpXIONrGuch2VRFwbMQ3aWB77A82CT9Qg8Be/qDE2
oROc2SBIx7m7UgdFTRu7466UNEuxP/2h3wJp2ds6hKCVkr7GomVTqtJhnk9pGGJO
PDe9FBeQvGxhUMZaMigPJbhcPWf6Tb5GM3MruPTl5WZyWP/owCMsNTb1JB/QsYHi
eTkRRFvGdowKZFoq8bXF6NPRsEMNSQ+/+2wWatBKXIolhFptzHYm3RrEINMZkVHo
RD32CCFdyvt2KRsy6jLrLTO2+m9zQLqv48Yk3zs6xkhDwwj2FSGUplD+XLy7ma6D
6uE2WMcFbbW7JVE2kTeCX614yZj7ALpEpOU0nv+sNTXk058gMQKkjEXEIiPqddii
TrBwaag5DpyJGudtep7G23QXyfQtTc61TqZ0LDh+yyIL7xUvdZoz1xAonhFnYwDe
I5uAzdNH4kZkw9UhbhYQKKz+YgKoBZ3jDWRVQQjsQTUDbZe/SMGiiwRuZyXNIdID
`pragma protect end_protected
