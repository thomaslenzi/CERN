// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:07 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kSbnxk5rJ9kRphrgmpjkF9QaLtUS2iW9RJQrUA3qCquk4TXx0WB4+cxP+Z3bwwV/
MohbKCDpPlI8OlvNYQwmK2xBOWYgNrNOJ3vgVH1ufPcxSAlwksOAUh1b+Vz0MjAJ
GwIQ0FAmzKEOfHdkWXI7gYefAqFVQSO/0Huvj1xltBw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 181168)
0Fi+hOrvq7rxk6cUZaxpp5+pZEBcHZ4oWi5yhcfM+crUkHKts2zLqal2hUtPok2h
w5cwIsBIm0ss/aDsXG+OOchnwlonYuoOJ5Pna/yA5//sbUfnUdmubA8kYfJ6dUPk
hZQK1ZcIwJ7glI0k9kL4U0rK3yuhXkn/a88+boDv2OA2JhNzytPIbELLiRB1+P9d
oTnBr54QUW2V0EZRr0PAJdY/AE0n4IQVKkb9Hvi0ilSfAxBn56EZJi7OGzGBB+hz
pUqF4Ly8+n914J74ZwuDgy2fDUCd70oFlRwlWOcqm9ZE35+ibzb8jtnoMBKloYr1
kZc24e5pGc4TXcQhsjXPQ1n799W8fDc/nXRvTefD/oP0//Km7qLgDGpXF8OeB1f2
4j93I0KqP7XYcQL3lf5BYecRqhKSKgHkrbU65s2c6YV+3/Vt6s1QNj/yaJVFTJoi
AkfzS/4MbVsl/RzmtYPpSDqTtKJY8/hWuO0YGMzwShOM7Vb1lN3AGU021uBq/2R6
EGnuvVoSdmub57JMc6Dtr5TwjGrz1fbfTwE5nq8eI+zSB/8JEYHabJzkLi/MDNpR
GSxpkrbVYx+fxWqDAzV+upm8asLCCfJWMKVa7tNnmxMHs8sg2MhAYeFVvJ4EdjeZ
IQ8TShLhX4F6dbVuwQNB8pSM57JREzvZb9OVqs2Rx81ssmbV+FI4qDd3T6gjEkuv
Wlnf1JmOvPmanUv/K9lp6Npw3d5qMXR5YmVYqSzL/s29o5jVrSBpNxiqnXGXJGyc
Ta5GU/9QMQfThABfTX3REr++JYa65W/JR7UqMCuac67oPwVzKIOXpYRIhWWngA2P
a/xyFevPQjh+4z5Kt2nQSDb+rdJ8Fw0ukw1OdeQerh+Q73pwEkT3lARgkFeOOvYE
xh25W4txDxxW3PCSW09lDTWUFHSw8UtoLrsB6XM9SLhZ5ib8bpmB2pFlO0zLdHOC
llIYFTJigJ8KQIhLR9t5VYZXs0EK+V1CxuvaMkm485HqQWX8CG6S1Bo9yZTWbIAR
jW061/04A8yiG2QAYKMhPIrbPFoGa6FwwIPcCuH8Z9GXZmk0/FJBvRKoEc3dDNSK
oYxqrzY0rU8mmwkGmtBE3b7m697snv616LC7LbLZGdALW1FIy+EzhQ87/7kfCG0J
HE4DEAimYafGGhY5FNn5cdjtF1BIHkt1DomV1pFzpfwqrHxKkaGY8JSjzkOkSo7h
tPGNxcbX/l91K2WAYK4vHKUlSYOBsRDUyzHRZKHv7RbkkJBNY4i7ln1JelyLUG3g
L4lnz8go/cnrJK8GE2fI/eNXc29PjMfyNdTpbojdNm+ne3t0D2ilTI4LXlJnLFYD
5WCfrGgsRjakXq63m1LuWOoMaYz5Pg9A/hc9UanYoAdQmuTdgaGuuY0j0h8tgHim
+LaL/9AU6LtVAiBhNSxkb0h7PANiMCY9dV6F99soJfwt+fH7ouMG/8ono9u0/sKv
8MrQvPiOGrWemZwPetRF8kUfWN45XfgmV5XXqB4m1hwx21FyZ08Xpo19rar9FOXX
DQlX2qWiQ75I96/zPIw0STihY3ADGgJWAY12bbWIY5lfH0i598dzUB/GiAY+zYcE
htM+bDK/qYza4kvvzH2HMsEio9l7Gs4npAmqQLYfTziF2s/Aek8NZN9bonkyg9UO
lXQd/rF46bdb0hh1d1R9W8mOwOX+9BBd9YA/NQdfJ7zWQCT/ldxHYYgZpn1qVUNT
jQg6HEBufG1udvYsf+DPC3nwkg4Uv80+YGtxnM1JGSQUivMLkAWRy0m3DOSZQ3S7
fMx7EY39uUVTlx1VBH1VYhkYqQ156EjXw/G0WS5nteIjBkz8mF5r8P68q8DTuHuo
bb3BWu+ZRPrmJx+lFq6KSTD4aaBNW9cdBDw/ol16cfF2u2qUq6K+e7acHlfe35aY
PbKd9BqrzvIE9RazCIMl35sZ9AAQJgrBjyy0n5EOU+yOu6eQ91udR0N+zpa9rAJ1
iU36U5Gf7ZvRyGawu6NSlPYvRG6RJNqE7BZo/hrySIb/5a75UzcTBXvC1VX2yZc+
HTUYxNp4L61tmZ0AdheXSjWQHr4c/DFGgTEZmmYvh23E0PCYsqLEcGbw2KNzs+J2
RBUog1+/hWqMI2y9dCNRrJZlZ+GVBA+nootQJs+xBOHwCvVmhIUl4Cpst/VSFEGu
E0+FkuM9/CZNu43hu1ug40gbZRmVQp4PwdEpEtbEX7A5WIThyX6p8LC+i1LsCHCi
t7Coj5CXcPryDlv0T/NqTnsdcQ+ygELquHCTz4ZuaF7Kk4r1u4uQ+c6Nchd4425V
dPhrq5KWh++KXO8Np5IqJAVVwlXoCIaNdE7EFPtO/03H6/dR2NXnU46rTgC/6FQW
Juco3ZJ1Af+8BMF4FXtw2uVlBrt9zadKjmFONCTAAxJcGZz4RyCuwoMxrM1K92eY
ZTDX2qM6er392sZMwPeWJBp4RNd4yTSq/c1PgQ/9ShOC5S5u3IYiBDPilX5KvGVE
mbmFGX4kxe7ttJ/DdF0D1B2r2c9SIvIGoV3ganKnrXq0Ah1AhLegyzxiGTXSTpGM
L27lCnq/3QuwN5NKLPMGtwtpHYQKIRxyav/5wpMhKaCz6MsqB+m8uAbztntXZ725
XGFn/cPavuZan1Msiqw1n5+4kPLpCdd+/UirHnpMhQTOlNioDXZRpBmC/Tmke6Jw
V+a1+sX+s3AWlVvHjayGe7J+eCpxqQPSuNb0oLwYOl8jqKC2xDVPdKcwXx5uGjOo
3luFJdo3jziSeOUY+ha/xbALgWkIlB4Kk9ISM0fdfZJzk1zt6aFZILP5/EY9wGrm
eoObTxVUbFWdTJfDWIZZnO82J2hdU8/oN5tYS4L5hHieEyKUL8Bllocz4W6m1qEp
r7CXkWyc5vTnEHvjNszAIckUCnvI4E7oxU6p2SwzK95nplHCqoodf9Xe6AdCmiv7
MvUrErusB2f8PfUgQ++Iuwit5ILrqwHr3wBTW11zPno/YUcrWJLzPxrsgQ9Ju/N/
/NKWXuJlnaS2QDYgXkC+e6hBwFzuE/m4R+qbKn3CpQJO8siFR78W/mKsYc+0evTU
JEUfGaf/lZpeDb4tN5DMPUJvr3ESZthhJG96xJxsoeKZkt7q5GRoDl9J10mhhQFk
meQrH4mdKTiQ1lZrOrTtbrn4OecvoQrJw8rmNMyp3dEDjJsr9T/uEQ314SBkwtej
xbvkvw/Qw30iVMw0KPQ3E3d9OwPflq/FcUBMkJs8LUiBEIYPATBU3MuBE24rISk2
dIXveIiHyeHB4vOI93z+AwlxOk88H8oiKFT/Cr1c2eSY+5LiZFeXBDYJL3nWev0z
f/CK4rDDFbPC5qqEr5NZQsN1RrSiJPKpVdoS/io7aGSn0lD9js2HuqrV0rnrZOm/
9l3JOwvLNn+2j7fagKIL5v43uDxgHqAPKbcuODSOJfIzTXqs9rG7CQomwEKSuY63
DrIV2TgCnYm6Dh/yFwa0fV+/QWNtxv08bHDwMS/VuwL6kE2jYIGDfqJDiBnUIwiN
x5ETYxr7Y37HEV871A60Y6QkY7e2q0Fn7XJlOcA2ETx9QRNQ6LHA1E+cP24xSvtS
mShsP7JmUOjmY1Zm4Y4bphMdEYcaAEqBLmy3eFwSZ5WDTvLuNrnGpH+rF3w8RPRp
Ze2YhIKxh107EA7Q3AFj4BDMtDK81wI8Gi6P2iigP85ekIOUDTiQQdF1gW3wJYkB
uyk8NBGb/TllSWv4Zg4NLBC+2lToXhBi526weTXTqCI8SqmOGrkzy1aVn0+QYTE1
tjm8iGyE8BZQis3XzwJiHsP5c/lAHDL8UdoGkRGNfZJcUu4LbXubUHTHW4asIGgg
2u6VHgA2eWURodk0RnLydJGYF7GSYBxvKdJiArcG/zfaIUHo/9iqkuq05kiV/uyJ
uI5qHA2SF4jwYsicMtwnCHM0JKSGYMOkZdLZLG+C0wCXEovvAagrPII50WZ4/GOG
hL/5J7kNl6+azgpbWtGtVGuKORAvcKwCkPAMUKD5C3ml1Z5gX4n18fM6p1CdQisp
wWRBlTjxKBVAX8nVXp5fiogxXJ8VuMh8BdPq5L3NrUyufUZefk33thQCJO4wiPHx
8mCTX/8VRevNS5vlkND6HN24BmlvtDWRfiBzi+1pUITxzY7LHQ2Rye2ldtCO2JU2
zKiQriO7Rot9uZd0AGw5FUtC3i6no8OeMGBqkP/ikIV3YdWPB/BM6gAR0nUssaI4
GSMUShvCBiTu9xVn/cPHvjVjPh27MnJprrgFN1y9NG0hU3L8t5pshAV7wMS88Cpx
RjbVBld4Rl9JbGPmOEhK1ferOUP5o8CIQzZa3fCOBs75yFGc4jEyZPID5WlEwYCl
1+QXiZiq4KJoAZHrLQjS7z7m0ZXi2OKiFu6TNl/jEIphEfAeuEit9uamq0Xryn0+
3LpM7LNoDDgPkCe6+TsMoHUNA3fIVRHGw5VkxKHlqmCAFIhdT5TDEUtGVev7uY6I
I92J0U09uBLzTbHMpuq0LYJFie51ewCLqON8a8/qxSV85fHwe673i8pSJwBPs50Z
rbDUV44DVNx77tuAJSmqtMeaWWey+Ay3kwfh3c1/tc78SnQyIX4gQvpez21v30L3
Ogje/kQ1GdllxzFwe5tCvbb7GI+cV0wAV1xXRsutwatFGPssIJp9dW4QmBRSJuet
GduO77oAYd4HjgQcs1QoXTnoSqK3xYL1sBMDNZLR0U95YR1ggd7mNsR5UJ1IujLS
q9RzRx/0o+oYokgfk6TASP8mGmR895Z08+EXCuV4mHY8a+uxlxS1g/mfP1JOa35S
0rToJrvlc89Oxqec8fAub+A2HxtjrgNOdjEoonAAqqZ99mNpjIDqygxOEDRQ6Zkk
o6Fi1gu6EhBxCAggkj513zN/TREM9xxXWqAmbvQQecsBw2qvsltnfnea+wvUqqgU
S6AEMx/JXr0qqifUnEYLjXkxAohhYwey97NppO4iPYxXcNRgj9+anRMuWse/+O6K
PK6DVTQodcsR9E7ngUZI62KVqVJyrS25KDmoyo5riQWaNF3HPvir9LvvuJPrqg3Q
OrV96HcNipLwZt5OdT5dqnlhq/dfhE5xm492N5144rC/K+1vdCWx5Up7FrWc//G/
ItiEPpjcx2WNSxKc/9ZVaExeyDTjh/dLsq6jF3Sd7KMhBIvvEzgT2aolCmEwUDKM
uM1Mp/dFFpdKscNIPVIuwMy4J7IQtKvE5C2BLdGK8mzDYU1tteBgF7sdaIv2f9ua
UZ700e2t9eqPRhhFyhtI+kQ/rGWsgHTcSXrzHBeV/Wq8KjjdwzrBSrcjwo2Db+MT
94FacWGWmM9Q4IW/LIjUNIVC8/ywtULPmwsNPjl4/oVHxDgvprRvcN1FRo3aEXym
8forHQMlU0Uvh5JXpXFISMOGIrCEFJxsw6oT4YA2+Zro0oFuSg36/4UQz7vSO78F
J7MVds9RXLg0OYTSGIWGucURKCQeGFE6nftFXOT8v/nShgH712h9G9uB1br7Jl9K
HF/xjdXibUCqrrxhyGJfrbsfZFro9ReSBDmQiZxYZPupP03eBHyMgbGFWwxVrE+O
INFf19EbmLxVHg5xQzmVH7YqMjevu5p8+yjGzSR4fOV5Z2vbyJTqH7ZJDOP8WGRY
9NXzFIMwLqoh6S27TQQbbDzYQjW14CrHggJNlnEQ5p+C7TPT/5p+SQiPNwojOsFZ
qe442oGjmlcXz0rZeJeNTlRYxgyLqtUqMWIUhHBcrU+EhDDC3bexIyXk73ClT4Uw
vGwJbmTMGLbMGV5eFMePNruTUuE6b705v4bvh2WkUrP2novFYZXVFRVXpwWuBTE+
piHfnPo7r6H5926EgvOSg5mo6GKPdMRMUhthNM6m6ETCRbUwAD6wQs0YnuFjBhD0
36iJVxrqyVxO9JskKVcGpOmYXknIa85RfLw0N5kZSzXznqRirB9M08qzf3FqnQjG
PelYEU1mQFXr1Ogj+Ht9DM0enLMu6x+zNH7IcOEP4GaASuwEDoTZECOku6+vd82c
WZT0mGp6xnjL5dEJBG8DTA/k3H4TBqm0sHW0lr8gAd9ggDmEseN7XFJ1LqBijnw5
8vF2KrHbshcgMvlzkldkBy+0hvu65hdOzmGUWdVubtEicQOjAN/pekfdfnEGdfMR
FgA+DzyX4HcZ23hjXoDiwWlYiKeshSSVFT9WqBaAaKHxSX/LjxbhfCPHeLp2pE19
c10W9jx7fLycgDMvthunj9E2jZiCj4ukd6w3JF5lhluL+Ir2WDYgFMJ2uCeh7HOT
qZkvjv1IHH3XdKG6q9Pzn6sqplSST5Zn0Mr/erZ8/N2ssiyCJDqTW0sIRcNjgycT
hM6bqvXEp3msB3IraFy5pkt3S25/O6VzA8q8nZVz9szjdN+96ntfuWs8bYwpFjA/
ad5piNv+81q9JpnE8eT8egwTUNqBtvL+A0rnl28j/b224Hd28aQxGt6fKBW9oi/X
YmKIaCsW+qhMATGd/FFuYOdo1kiGSXGfkirmO2OzSgwe51kk8DLgWSAR6TACcZTM
+ufJxOJ8N+8NViHN1kvHNAewp0Cdjwu/z2vraCFDvyrqiZZjzZ5as6DGLXZckHg9
SQ+kOstHuwebXkNqtd4g0F5bZvdz8CIK0+ReevOJVton7EIX/ErXq922c1ImZSJj
x3F00xDzY571/H/lYsnWHxBIhC8gFGqqPvK3uNaMfoBkgf+UkfqpM3g1o+l0O1Pz
Wid95yF6cqoIya/ow7zCPmAmsFdBpQsxULbWAHziG80vAVacdK6glfRtJ1spvHdi
cVA9iSKre3NkCRSHQdvIAB90X04yX+BJta3HMF90BQGGE6wzuvOABjsaXFJz4LzW
Xfnz3hv1pFYWMFMz5/2x5KTiftQkFjitlFR7jgovHUjC/aebmMGKEcvtsZ5SxMg4
l0UL+qTOZqHRceyegc4k3QCm9axavTbUMkAooO6JIKzmmeIa8Gkj/K0O+GOknvtw
jPheoXwUHyXC3GVwXfk1TK/1USLjJFxuDc16Z6waApD0cjxRYaY8itrXiCQBwFqj
t3H5F6Qx8mjzu81M6qv2AEfZZyfKQsLkeqz9K0ZfuHxgNFl6k1o5ZLnuM1RCQlCo
UvQGwyllGQCfM7U4u4r/876m9Hq75TbM73P8GIBgkoo4k3YuineVBz2XZDZo7kO4
6/GJOhsscWiRpuZiyAVXEl8jC+EaxjChvVTGM6SsARdM6ixsuK+yxRmFr7wAsXHv
a/Red31blEuZUFJZEf8DizGpsY3GV2MgplgRCXQCD6fFwjYYKvQDcm1qQQWWl6bo
eUwejS3/UT+YICx/ZmCU8ZtpReG9NHD16js1PS85o/4/lcr43rbx/ZiJdS8RDLGb
QsZBdyNJGSUsDoDEOhgb49AN7GYPybUvxf23Zp765qvvIwMySxfTSX8LaMMo/5ZF
cxPWBewijZeow7p4WhYOPdKtQjuVJxeba0TYxuY7HRrLE2Tupj+MgE5IfFJmB1pn
PXxain4dHOzteOxGPVCfmdNibmQMIG9KI8xSAEDji25Fk8gglhATdYLS0roC7VX1
tUDbAoKF/690PU238p0Shm2y0eV6xZ9nuMRPg/x5iqPEjr3uzeUROLR5IDU6NTQN
Z+QRWWYuK/rRKOvuqf3rTFDJSJR664kJl6q3kTB0HXGDlBZVmM+AEAOm8TjjSvT/
fE/QXXrds0HqhNuhnPT+xDUTiDaQGjhEklhBiT+pHyDYJHcFZQW9ztFH7uhk5xbc
ZmRuZf4RwRKpU78ZpdSkZQBe6Fo5n6usV2JuzOEyJmAQD83CT3Z7mxR3J4YzvrwG
JCBuC6ehSrU7Z5xacX8SjNDxOVpToxl2OgL9a6/g8M7obwRq3keLVBUFawUXC4Xs
+mCNpZ9q1ijPC4uTZBdTZAyJDn+79ZNxb8IgZXiBMpMgn1CkBjickIgsR6bX92oD
r1IzYtjDB2S304J/LLFT0lqoGVrqPMQLps7V7D4sCKGyjbTYOi4frkW3TJcfbhLn
gCyFdJKLgCUaDbrwHRAX46TLMUTU1SlWi1tQ5I/mvZpmMqloDon5qr273fEpxHuc
jSTJDokg5sDIdsY42sl2kxSLuRG6gPfATZ8yV96BHbRkW/iG24q01NwHbAqtJUlI
Q2xqxkuFabyZzmNt1LMrckJnhaOwCstWeNNBEnZcNYKHKLIZakEvUZoYtq0JNQlz
KdW7bGXiyTKVPE9KhzzL1oq3mmbfH4m/fk2ErQuvJmM35RvnNc4DfpAILFiZw35C
sbP+idEs+9v3wdzRZWn1nDV6baG5qeGneUOcee/yCJfHmkVVOQKZLeasv/ZZlV5a
zjpfwQgRcVpU3qx+3r0aw2B4fHI0jk75wQBfCpwz0FownE1Urz7Gsii+0IhMoEAa
cSvngEyN9jYTt9etr0bxt+x0axfcF/HsP9d3pw7z8zfDeMMclqPWG9eN5SZlYmRi
t1ZaOdHrSgih7QrnoEJ8setG+zlYr+EQNhaKWEvlsBAy5AbJ6BsNNxLREi/RoUBk
Vd/dQUXItU6f8vslxDyu0s3H31X4iiDNDtyYjB88VbUh/ug7TIMca+XmD3juCeoi
qo/IORCPbqdxEHkscYVjVwJdGxDiSX58OtsYaMyaKyRb7NUGpyJFUF8f49wK77bQ
Qwj9ve7ps9ovRsmGCFrO4Zkp0mCb6YXFvgd6L0S4KGwBqiep8ahhxLqnvUohGRA9
yCQvRjhRcHVHldUwQqedbAJ738r6ZtBpkJ51zHlqhdKM7ymAPO1GGsTvSnQxBNfg
LlHFTqOzUTID5C9KywDrljjRIWagyK0D6bs8Q3qzAQB/Y/xv7T8hlrJxUg16Orrv
/UMCVurX777JakkwpSm9fNsxEWeEmtfXeOnwswwzaFBvpysw3Oy+JkiuKUQ5jKwh
p+4n2gPEiNc2ap2lspGzEylWqR1prl/XP6MgnAX+MUQ6UpjnyNBmRNv5yd45Iq6+
GrT5NsSWYvyHMtYr/Z9xIC/rN+ru5z9e35D3kVYsuXv054RXYwBCnJ+MRC8fP7Gt
1e3AHZCb5b8G1hJZurNcvXyVPLwJSi+7QansQ7GBxWEAcU9YVFGadaBDSsZmcHTV
J7YU0APedDFb/SEPaSu1z7qzfNqZzFYSWwokAABUhWKo1i7yZl1M8YKgsSWjmLqU
VMDMfZxWnYcWhPLf5lNzjtCgbktAWMwZxCPfM6yUSpvTeClBvcb+eSqqdaAD2eUu
lPTsenxU2qfFmmu1z6if8LN8bCaSUroYhm4QMH/ncwyvk2ISwi8NcerloKHGFGgd
R9Q1KIhAnDbTbxTqBdcujVe3b0W45i3bVJ21HhDVBTHsXO9FCNKu3GZqKFqneDBr
9wlabUfidqcdFZ9mHwpb63NJFt68ZPcnaRAl5x8o477/nPIR8o7l52Whiy8931bS
gkgSJcLqfXq2/AS/dRHQN8QQEQOavKCcZsLVnlBKmKpf1RXADgYCKfztnSR2IvOr
WqBKh54M9nPdjvXEyYIw8eaxinZeV+JpovaYfhD4jLbE2Q7D1QwN0TuhRRbj6aM5
28IxyxDAQo4kC1d797sggTdGGPhSZBUIgHgKD1ZJTrqCEUWFmQN/hfi7W0WDldQC
beEe2pRBsa/NrndL/346fXKlE3MHa4PtoLr6oR6tStldVbj9iUzIVgEgPA8xCZbR
Ysre/C0d/jfuO3y5QM9o/LwnEmsZBL4d5sK0WgBzgvufhPsPp/N/NzyjPuXgJHk0
sl2jLWLn1GrKxijzd9fMT3VSN4UBOoy4GFz/ftsCshNMQgQEpkoNsZeYJ2rHKzQ6
bFLqJbV68BV75BvtiMYyDoL0AB//v9Nn9+tm31tuLr+f+kTr+za8jr/+i1Ik/mYZ
dTIrEgX9EAJYpdh/BYLARQgGoB+Nz3KeA1UTzHb5j3zcvlTCqBbP/qMb2t6aLFdX
HCxv5Zsee1OrPNtJNJ7c8PQr9gFJJp6HulT3eFBD6arukOR4y0EhN/NVRAxFObF/
VlfJpNUxL6kRhwBctIrkDXyj9jlAXzBOrpLuelp6N1nlEtklt38W8tK0c/3JMQt/
KNWTX1+QclqkTJaU+SZ1OKA8RaxUiqyQwgsK3WTrJUJ/f4GcpF8bopUTgxSBXIOU
2nnF69Cp5VNNRpishH5MC304YsMco9NjvjmH24LeshUqaE5pK4N7TzVV1Qwox2UO
L8UQIn+A3hzrnmIO+1QXUERZkQdXW9OJ36W1H1SB0HxK20Wd/yWrMKmZCiAWW/G+
v7q8V3/GFArMYAqC/LK/v2Dw0iE++UIG+dZOv6qEz5c9C8ZyazQKjjY79OGL2QyS
Jd3ZfHG8ujPrQ4FdKqherKSk/h25bIpnvpCOI33aCgLn3dVJuqKTBNGWQ8XaD4B4
udK5uGnXAA9W2Ebid+19nhJVdeq4WAB447t++cJHJZBL7if+ICPfB2yiVTl4fOiC
+f4QnlHc9Emikh30Q8bGf8Q/pGScDQngapDoEIF1RjsuBz729R1quLFM/4byHdPb
OVbqEY2cwacv3AqrIDVy9PL/NP94/6P16NPEnyzIW+eO+EXgdKiJyR8yN+KvbaFY
gRJhGqKcdFOlwvpMHsBm4AFAHJpmaVF9AMnngIGiofJkZr6oKaZmjUjc3EiQu9LL
OU2A0TCFbzmcJRZtAykho9a0VfdfwQ32dP+iDwA1F0OUDNERmuwHuZIC0Lb9FmbY
E8MIFgAq4BJSeGw2J1RSsJKQzQmeW+TBQWbNvjIpxCwJJWZCWgngNKv1jJlrWuyN
61YJjJW1k+mDa35/7h/N1jjitWpf4JjHv0qYY5EhrcO8BicjdkQ3aAMu32Zqz88R
6e/qAF7SVHj35hLRWcs+r8eCscZJ2jsLxFNpqFIfdrtB4b2KiKKxpgTnUIdS5qDd
wvtLi4X+0ZR9AMPgNNYutO9M4zONicZrtb2I58AQKM9xe64kqo6nkd88YPM3sr52
jUMhBJd7ddP9nJn8O4wnknzY4mZpdtIAxpBNiJqZsgvHbPkqz8fCkwiCamIHabYV
SGQqNBWdQ8tjAMXXd+6uiaoEpRN5+L0ghOHn8qM9bnT1ygD3nRIMrYnsAf48Tn/w
7TpzTYz/+LJWnp0qwTVycseC4S6Ath/Lbzxhl/kr6ioEgAsF/eCflQwyKSD4Y0/2
yVPcbMAF9Jd07Q+uGCrnLY3fqxHc68uoP3G20kfKlHdFr/lqz/kq8v5jiTQHID2L
/Q/jlBAliRHYxLwySoxy4adJelH5vdJ4z9+AwyusJjxBlttMtyN0AievsQBxED+2
E0601oAqdb2XKkOX7/zKULJEJHDSphAVIJGwGdwBtf7V1r/zCKIp9lKkGdJ8l6fI
3qUPAPtboE+0S0Q5++r4uyKJl/RPvpZONj6a9NFcSrzV41oBvX9mvTF/WkCIdT0Y
83ep6uCRmtVNcStCz9GafnfaRH4eQdzsuFw5iqndaALj3idGNXf+0n/Qqy+UOQs4
26UhC7zaJYmDV8K9P82C8t5UZ53IUzDMz+WauEY06iqGAjRdeWMe9t/dKC8cgnyr
OLYheV02t25jCHlYrlkItkuq6rq6CvmBL6kOsGEXb0f35MwycRkLET97sGp25Z5l
9bBUq2WpmsoiBgRRJQ6Ee8lHXXndcpeYYcLmFiLzhDPhohuKAgdbHFAC1ffLmP9a
Ex6iHDsrIUk6o0p5KTfu2MEOAm9+eiVPEWU6CGVU5x/sBOu550Ze8HUormjX/lkf
Pi2W1SI6fI8En4VVGn+NpGHfC3u10nlBPHoj0Xfp6O2ai5fQuHnICA76p6v9gd8u
1k1yVbTw5ZOQvRoueUZRFKlae5uEqbumbgFJ8zMa7AtJWem58QBxRhro/f0xnSEp
iLhPbrjCts8Wwj85y/jChy7JtychXrkALWVSBrm9xDnGxrown03xSPCrM/tJUAvk
g4Lbg9djQytamypKpuSZ0gwoOfMuEVXbIOCw3DS26MvwPqHikF3PGtEsymEOFTp4
jXGHd7kkUFXUl0pCNomwMKZ6LSdhIfYU77lxnHGeWgyv0DWrDdb/CS0NQvUClM+6
FQ6HN1KQtHabtu88BfN73mfN49ClaN39TWNO4s51RJOVu4N+mIXaimzb9iazGxcZ
g7jNAszotozaF60hRlzlvTWx1HckM+GWtSk1fySfWxO2HWIViy1Vc5yBHOE65X8a
+TM8mE2N9RLFxYU/ejZS8ErttwSWIg6vZWLytkjYJod6DaqXpBXG6/loEJq4x/hb
gEUdouCDkzb9QxvR1FwDWjxSI5GSBLxpox2KxBTjQdyXhPbtdMS+V95WvVKqFZ/X
AVo1TH6WnrpY3e8IlcOfzBdUC2mfzUYHZVYzuJJy/wmcNoB+ZAK9vkI/hRCoZXpt
DaPqh1v3MY7TLZWO09L5OhGtKW/ccX/L4bcJvEH07LdlFXzMZIBX+EHISvuEKFIu
2T9neNbbdspI0uRCWLl1BWm8Emd3kFL0IvxRUsuEEzdbXMiEw21IJgmg24JaFdiC
VBDnJjce+jvxAbZkARAWI8yMZVrDtLSsc7FgJn7E/CYJeRgr27cMbkGjupIxE+cz
bxklyEfvxU1AgKSn6hWKSXPsVRQ2LUzc5NUS3OgCpN2jnpzbNZbtwT8nqTGb6qnC
9d91GwInI5XxWZ57L2QRs0E4yNWxkXNdRiCo2195qogAd8LSKJkItMm7F9KKRQOF
JHs5P7kOFydMv5GXM7ZTZFZy/DnryGFIP+BGG6o7Jyee6kqnj5T9/3iANRiRFQGE
3NPWPXCNWXuS3hQShtMaC+zJtNiYXph24tynxEE+VVwD/MxNakWmQw3OuLQTCH7/
a9SMCkomIdIyMhwm7mh6Tf6HeElUSHZWJ8CnQYzUvQHe0XKNO4m4d/50a3idV6KX
OW8Zb9qc7KE77sr9OFde8ARTkM35m6CVZRA/1xM8TXUKurdIcl1rtrFnPJLBiK9F
Qolp3GMx0nhpH7c14Yw0tk//w4ihukmt4odjJdvtgXG++BwcB9ccpbwFt//i+rPd
S5soAiSFdZ/hvvzzHpuWg/jSK4UPQdjfQ16GnRAnNTktsHkGPwOz0/Rru9XO3SYZ
UZycDXA2qnkrRTmBMp76PFGw9ifrGFqxjZtMed9Ax/yQ+DrSLzsfY8n+YhAYKaRz
L3uySFUvnWwxcOUZ5MiPFSbFxatL8nEb6OHx1xbVk147J/rV12TEbMH08MNFPY4t
mYp3V9QZTE7cFtWEtv7v2yBOwyghUBDyAjqUu4AT52EoFSKIhEQ5aZenqFNnMon3
1Cj2jkbTnmy9NCAv91x/i+pwgWibmF79Ne11JbzcInGHEXPOxMisCdiBmR1a+A6D
HlxpGb8eUBvWz2mqEWMqbfnV2k/BQ2RkwJ2P6PUs2HTYKpg1WuBMzF90F1ZJEChx
0kqBnLG23jj42b474wGM/qy+dMPjnD0qhytZWvK3YZdg8zb0p23kVUvruaN/ENiK
dbq31TJN45vJSm2/s46FyA+f1F3iV0pUKCD8kY8P786r83KaHq30jiHohdkfmfF5
B+ntkjzI0Kd0EN+IzGEGmAE6LahNKH3AT9IeYPUpP6WJ4wkSwK2WFV1LxyVMrl9L
SP5/l1rVV3tKrm2I6zBGAOXEsrJLlLPUhKfxfhfXfYiyHNRPgb1AP0kwfDe17so/
Mw/r4vntVydd0e6INgTvdwaENXZsX2P9pq18fRAboxRteiJASfuyCMS6c1m6BBEv
6CEaEm6nnlTyA8mIf4ooHgTSyOOmw442uRsUHErIfeqOSQrpLRy1oLpJOoCin11u
Pmf83mMu6npYP14vLPobUzFLtX6QqR3PeD08jQ2YejK3mkgJtbXysO1X7/B0PsjU
ISDZXEuud3hNSawc9rQ8uiU0p483xc63ymjziy9tI56G9c/9wPSiS3wpAenl0x+b
nHwh7Cf7l8Y7BwBWanDwSh9HvzNS52SP2XDKIBZ0UeUi4wfNOZZXJR0+TMB9llVI
WFAQ1iuPPRpejWnX53OV8hi7thA+o78+OPtWF1ef6x8vWnd8tSICQXKjYMhUwU/w
qI7eiI/+DAcP3T7dR6jjjL/uR1z8iVbn3ro7w5kmX/PPPgGq/Yg4zwS4t0Xry7yK
CSlLvQjv38eiFa2xZAddRfytdUfRprmr6/beGhKEy/tVAXWFW+MzXp/iY9DS35qJ
c1QN5NKzHaTnFkhLj2wOkCORBVufg1KTmjIDcDv3GkrSb47S2l8f34WPVovHXSeL
M0AFMkVqs134g5nfrexsaXFgtAaKS2ueLv0RrVOCJdF7biFDwo6gFGriAssGMLvc
B+kS4jT1BOPXMxbK/PlEVeJIbaoe+Yk56J/qNaqq6tTPaF8TNZqRDeHd9tJ6JkbE
Caf9xYrbKHl0U5N7mFhWgy6aC5p3pJ3twt4fVMn1qKRNhK9y2eQ0s9gM0m9BnOQc
7TFbeHjNT5GMG+57CX7zVOQT0vdPGH0IY+URX3sNMgefl5aN9f8wosYU/tva4cLx
CGlatWZOoD2txkJE37HBTTkF5vNRjDGStxi0czP/QtkC42AAoYipT3N7Snp20vnD
WtS9ntWNR7oJiPqG9ZRjfSZ98Z+gSSkg4Yr8om+xeavaYeqsImUyfKY0j4FhoIzN
19EnPVCfetQFHN0LqoODhjVJUeN3UvfUXfGSsXYaYL8e7LA1OAI3wl48n04ToBtJ
26fBEvgpbiZt1VDSDjjwHvSzJQ/l6+pjdrRP2pZr2Jm7qgJnY3/NzXLn6ZqLb661
qAUvzkzVs1n9lpg91D2pCnIYJAlkO+s2KETRhvjWsCyOQ653LD+AnLKeo523GTYe
FgTlnlWJKJ6UidDif5b2DTmCTl7tqnRLyGYGItsKuQ6OsA3SuCDOkSpfh+6Yypdn
EkXj6lwY+wszdFpImjkR8mSSU7XDj1qOlZqlbSlLrijUdZ+7jsILeygP30r9PWfU
KEqp6ydjSnQU9gTlIcf7xOeXU7hx3z7j3AuCUjx17wUpFTuUsKo8qrgQGXvNkWbV
JuGcmHBKqn/M2zhiH8lCVxVeHLUsy4y7eAf0V0GQhCYcEcrGhjug7W4Qxy73fNt3
2snEsn+Kc8obJtmrKvAUbEOOF8/WGXcKsaBQqOFFIvmcSqdqUuo8/XOZctn/K5om
zEB+ab6S5riQFy/6qAvEdWPf6KJx5BZT0rQywhdFrRr7/End0gVxm/kLo1niblpv
nupxfO1D9RABnCbUO9u221PpCk/mxufVwXo1aCK6gj+mDDJprQa/GlWO8uC8YvDi
FHy73puGUCoH22xHpfL75I3mxeh0OUdospf2EUOy19IYpWA49Oooxkt04dm9WFvQ
L/81/FkdcJr/e0HJq4mi/7jD/qRgpoad3Z/kpy7fl/eJx4odxc+/uz/vPaYw7F/W
UatltmDrZLa/m2D8Uj+R6/wSOxjKyfYzU/hJCeh6jtydguXOItIY4jBsQTQtM/GB
vhsUUit+cXONkmKuZaOYzSLvsBkarHspemPVgoj2kh9I0OcywiDn/rpe+mBr4eR+
6dxslIbYNoi+Vo0XflMx8haRkiF4WquzyFGi8RFXqXXQrkuGTcQOu6Cz0UkXRtP/
yQFCr5qe1AaYq8ZIuEPY1DXx6nw4DaK946UTQXQZ6Milrgp2t5ST9HiNMkQzyXK5
sud13P7NDbMk167rmS4d7FtlA4Jfb+hChw/bhwIWi5bXGYBEV1cM4fYtgWQ8oJMI
sYPtm/jXFw0hNFHQU/R/G7Y2ax+XV80c1UC07PhUryqlCQYljj69yKaotcc9x9XN
mGJJ7GfXZg/3mjfjf95TmIVgAnN2fGPAuVKYoF7HnBRMNhrCF/kKutc88UwGCpuM
blKGj+TULbwLIM/xpsOO9WZc+81ANG8YgjdwlhZQtqrPBC2SC3r4Bl01CGX+RQ+s
V2hK1DaWMS+DDrzqCIx+xetlZBeza5iYiJylCKQLQ3UMZRkdaT9JXdzkXF/SWq1k
ERoR39UeD+jsad1WMwAv6zyG+//HZ92arizm7ZEt7ERl44Mc9MSPBFtv8ze9otfg
uyZqtLVgVsN9X2s/28XaVlJkid2MfqmcD7xR5DQzTqIUttn9/W8hdxvzwvae8tay
f4Zd1UTZaAy9ywKOQ9MYgmM+Bz+IebVK+M79CjHiD8O1aDzdv/oypC4oVIbB0OcF
K++JIS4NpWBCtg/Um2nCbbjpDi1H+IWgotguvbAYKxc+1zgJ40q5Rt/HwsmKI6LV
AdW+pHp/lm/3kF0PwdtrCvbnooW7fSbZTDEMDFB/OSFxQPn34Nqir+CyYAjJEswO
vViQValCPCjBBXytVWeuh8aZBlepwUUbDsZxJU2TgKEzGOkKeyXjJQdU0I7z58XQ
k+gS4Wyac0ygbAmWTjWBnPjIyY3XqswX85bCX5cNXqORbKLoLoPhjn1wkUo9f/GM
wicaRuurLNv3i6dMgrOag66vRnjuk5yDSGPbM+zNK8faNJlyB6nahDSFTd1ftSsy
/bZGK4aGzwJhzmqHB7a5cCf862cvbcXgRNc6sv7v51V1+OLO9UhbGwxbjlyg2rGE
opacWuIMY/wiEJY/qaWy7GMWJXXA3bihyvSNC8Pd0u3E8Y/PehSt2iGMgKspOmgA
lKJAwKPqRtvzJGPLRHzaCbmu4+ai8lQHR6E+E1uY7Jk2CSQrNQn3USGri2joDlc+
jau0dPMUPHHk+3nA2fLfBlA4gcDV8YN5BVwqTuMLVqOaoLkGWgH3Fpolt84sTCpY
Kh8RkzoHMbf1/F14LyDBR/gIocyVzQn/KkJw/PqRFL4hTNs3L5xcZt9MYcG1ohdy
EyZkmRMHsSy0N8XrZiPZtDHwf7uEzD89SmLKokrAQB9ZQGTpbUDJd/xCxKQxi4Zx
llM1oZQaRuPdtHnGWsoEW/j7jN0di9NuD8GSxJMB41kkiFopogB4qZQA8F5+YQz1
C6TPCJ/C7a5eTijCw2ny07YanzI6w8TpW5oE8KFqwlv6O2u1pn0Fwc+jp7KjPqUi
4DzBrX9icxtpUxOQftb4e60lY3C8cjolnb/4PBEhiXbq7SSqXdPFBPCNaWBF/VAd
7zdDnsm6z2gRx41XJf9yu6DTksxOkWU/TZNjOwHUOlyQEzvcVofMymANZti3N4OM
iWOESLypv0QPEBZFy1sC630X0ixSTwljKPqqS8vulPUgK4V1i4egg0PZyDfwDOCq
dl9DWRpvWEC3tgNqmIoVH21bZcpA8sls3COjm0iyfur+H+q8r6HP2xHO5ewZC33R
JboBvmnK/ma/eFn7MQ22+1GTMn9GIxmc228kDHdMt42/osmNeogbXD333GEOAY0/
EBmzunIs/oUbTpZPwMRsLj5wvd68OsQD3x7+rN4yPD7wcIyr0ObpyahcRs2CUdfZ
Ai5aNFyuJ0Q5Yz2MSg9W1uUiIPDvd5U9K2RTA+p708VVodJOnRTf5nEJ0c0kxNi4
4lTTuQBxGMyVoSQpOFFJebM36iSiFgL+15NL2phcj50/Ccr+GfZ0SNCRYJ5ElGOo
Vo1NyGr8+/favv1q7oO2XqlZJTwAoCl3L6VhktYFRIz+EhMar5iiexHjlpqJGIpD
hO1gVflR/BLSJU4nsQvR1wc3/9dhLnBgyFfHpGHRcDU7VE3zW0/yc00bvBNiZ+gW
54oRyJjBqXAq1ft9paowuMatGZOLiQmn53B+qGtuz1mcaUfzT9kXS6PjwKuTqven
MgVQZwoZPZhEqvmTU+G/vKU0fs6ak3p63NTzQKJkQB7FR4pM5q2YU/BiZYPLelbm
5yFGvAEEwLrEPncuXJvdoAAGnsPSMgjsHZD2QmxI+k8y85uHZZMGxtHU6FcQGW7t
5XLPQAdIRYOxVl3B16MG+5dGV9lVjB58peQqmomi/fSMhEEbgZb7jj53n59/msqE
4OEIT+KwylxLTi1uUwmfokahV8thm/3k84hZANcoACtdPHj4lu6qPaeawfM1bGYJ
CL/yqpQkxyFoZ6fe4cdPqVwAkS+Ig9qZzu3fZumXljm7Ma83zM8OpkTOYBi7z2Du
ABs0wIsEjsKziCYMfA6p6sn6M/J5XJGB5xDst7UtKHJLIvzkyaiCHSQYZE9/RlDw
/c+d12tPPmE1fcrfWAbN/DNERuGU0SV7STT/kfyp2zOI3f4YTYgrWuX5QvwmlbmE
c70YoLRBpd/CjbH7rQkShoMg7VNP5BTK9Nsq6lq0ix3afMmsT+qAe87utdU6YG1G
DPn2pkKqNK4J8k0FQiHIASkeeXSIUlMiXMfJSjHo1nlUXWrmcLOfANxo+cgLTar0
vwLv9qo6wR8SA2p3dzDrvr9ziVpfxKEon6jgQUszJ6wanVXhCWXqAo0cFylYZRu7
LG1RAgDhHXM9AEEt0KzwZTCpYWGkIQtwaWf2CVvvyY8L6SS5cmk5kbjQRiq0wY0N
8Ea1Yq7pQev9tUAKayl9vtHrapZwitABj1c/R66c0+B+pMHBhMEPyDWPfHh0aN5O
hjAzQk1OxHILBHkITGJwJYX6Eho3iRCdVJg+du/Bc5tk/ZFR3bTJyj/37RjnLSHi
v3CYLd64njpafKQtJwcClk7QkoF92ehdqbhBsfISRA+MlWxRjcxRwpTS1U7LaIqD
5gsHDipZ2PX7aQhUNfxrGWj5Kv4rUCUlAO2/DPeBRzOjkCE4fYADRn3xZhjSfYa1
+BF/yb2GDEriPz71srITo8cHO+WTcrKkoUoZhwUZ2wI1xuhiAloLnFxqgbcVbBf1
9TuLt/tRGqfmMD8paS/l3rmEDLd3qOpcpycsPRVTljSZ7sNSwgjNHluFI5aoaZ16
df5bNTPvpKpmbxtoOj7SOnmsjqP2CsKq0Gt/7rmhj6+ZfkgFyTGvnDdbJapUvrza
4fK6zR8MdM3VVLpL1Q3V6Y0xP7Ip8ckOVsid4W7zfRC98A4CNmuO4t8Wd9nj+jXF
aCEZ/Q94HsaVktOpq7CPODxRAGwsVfNGpALq/f+W8eByI7fQrWX1HBLApy7jEfpp
BnrPD3FBJqyh30oTYxQ/7596BN+/IcHEG2+5rJ2f7wURGd+AdlvSVzgfCh41fM7J
005BXC4nMoKIq95icijUCREHQhqMqr3eE/GLGJc+xQ1xp5KMYLEhE7iYE0wU8m9r
i7cY3oGH5eCN9LgUSvWMO/Gfsp5MaW59JzrjaVHTNAmLzhHPYwdcrV+xsyKWXh7W
PbK4DlFGFPlY12jnID1gOMjmIded5BI/gI+bDRYhTX30neFvHYE5F6f9X7wRz2Qk
zgqW8CNL+OSY3yl5e7rRY0qIYUW54LhgBG6jheCxIQWcE8H+E03pJQCsKHEVceAn
CPOtnMdLPRpThlc/E6QzKIbs11Muws6NZnTKjUT4TUmrCNr0FaUB3EUbS9KpjQ/z
7bZ7EngLZ3WfuGv8wqJ5VzM9KASN5eZf59apd11P1krkNw69KA+c1GRcR4Q+bzh/
gqso0CjyrG6qwwrsYZvJ/gqWl9++Y8LQXNkV88lYpV0cDtRYThJG2c34gMY8Au5t
kam6n44GW/6zmKi4z9UFMwD0xHUtqhNg2B0jFyQkUXpgv6y/+ubABBPpVJkcnY7w
HizpHSKvaJYFFBc5Stjj0d2wNxnuT+tuimd+CLD9DK7SvV9jeoyG2c/H5FbKwa53
JxQrF2ZIYi383wLskAgYJ3eyonwKHHPWdqIwyCvVBn8w7UM6or/557khQI6Due2S
9W1ti+t6co0ZzV1bgthCJs8tuwZMND/sd7/PIAUejq3kTE2R67VzY7p/ldPwuU1B
jZTusaPpFhLamCfjsrza4ddLhpx2p/dOdLcSDhGcqVzQeEHc5hd4oWLsA5lEZt2f
1+hdwvPT/NuQ0xMFoqWw37Iy/KPqtvs29y6I3oMxDqPSy5qSASLWn7O5fWo8zQ/K
Ghax/LzeVW+MJ6jJE8CARvAsjoy9CDgPveZ5OWhpsZatch07Pi4u5vg9cg/gNYjI
L7xLIA5gmakvMxvliwuS949WW1lGcH5+BrV1Or3Ee6VWio9ozTVF0rAhAtpalCJa
p3hhrQWut3N5IFQxcubp6cPyfwrM8Bdanu8Ss39sDeIO9IgtzMogTY/jhPdexBQu
pw36fI42tAT9DTuAuOnHAg61LpSnllN2rWovVFScGypIMkGKZXvBkPEQdFZPOQwq
yS50q71FuKhJ2DDrV8KLV5+WfaeJrnzXwD8YKag2TFFIVlfgCKFBsn0cpFsHzF13
EBGh/4Lnwt+UlL1bbo7sRKzB1jkZRh3ZZP0AisgVxf63lsAOFYewryHac4JIvhDr
YaHc1mLK4MQI2k/bBMXVsfDku9J6URtOs0eZiTEgcfaj4DaDlP9z9EFJd0ZFD7qx
uEvGk4+ouOyOYwlA7prFejbZdsgf7BiBqMzjNSGd4KZsmXd32RZJG2qZPWqRTB3N
3TV361xrFKLlZ7Foiy9Wn1PwhNIEeGbkg8zkOq+ESYJ89H9o5ivBisv9QgenQgJH
XOZFgIu/6asqzMjMEvsGpw+IS3G5wBk41CkBJW60MJpjvTGUJCyNyYmHSHAfDM6q
1mzeb0YeCcoQGcQlgokv5nBPqfosoEoYUeSUECblJN9TP0P8LDhD0auaZavftlyA
6mPY66wfciC1Q+1+6r5CPsg0xJZMhCA77WIPOSXpSQItQMIX1cZ6QwQQPaOZVJ4B
sdhrkcyMpIsO++WYV9Ea6qOBS2GgMlZuC+Wl+ABcafxhPVcggtuxGsGp3xjArBUu
lILvM89BKVixaQa6lJQgofWlIVJsKReKEYfRFtPEXJnx5cnmph8K3WeDi4Q5i1h+
3vPYMqukASqNPFKiDzkLlC9mm2KpyyTzD0gpBNE//TEFU3S1M5MEI6HAmS9PaAFb
vlQcJRlufHAabgT6dWCj4n0fJNf49Q05QN3k1HrJuR5eKFuO+JFCI/JmY0A+4ebG
vERW4iM/dtwRUwNh++11IRUJMAG3JJ5/foEq3cEgigfhI/h7yeaChcbaVM7VnMO+
UjpkEdlfMWrddjpp2ti5GZ65lSGOWkukDw2LbtkgSXmccJuCLEtXv6SjutFHdvyi
IAAXcgwwU84ndNI1p7HlKs9rhvfdH6ibVeR8pzS6c/ewhQ9ehZVfQHhVs2XDoKzX
R29spdN1dVL05vWjA9TAWvNA+RzjdnJPbhpTGbvNmucbUtbrmw9Naz1Y5RlF/+gZ
6CqDhmwhGsqF9OuOXc9lroRYK91crIKZ/VnhunLhw9QxbtcYpOa6r+BAFC7CAEjM
N/lTPatFoSVnnXAkGLEU0zmGAisCw7im+jtnWP3KLOUo9xi+Q4Ih5+Ez8iOrvFL/
uTNROWJFrYUN9kPupCX6JjyEvUFWoLRNQO99NlBhETJPDCOnO1kMU26gpk0oVcqR
Capm356g3hS8ymk3H8WQcryxAJ9GH3yaYvL+UeuLLFxuu16Rizf2YOUBJ8dUvzao
HTakc+mQIiSX0usyhbZ5ulAG1aTD0DGTAY0yvEkjHm9t3d6HBLxe9PDVyk1CGwgZ
DvykXT0zC775CQSR1ba8qlFTH5NSiSCbYPdFVbyx8x1IKC1go6dKRNF/rEklXFCB
nY3FqB6qB7BPOR61p0tuQF7e4lMltxKo4X/3Po3/l5n+MIttsRFiOt8fbb6Pvb8a
jwbEkGXh2GB7BsuiXF0aneuyDtqDVs6wqkX+HgTeR/hCussoL//6kf5eJH6dRHmQ
anB/Mwt7JNWbU7BqdRoebPBGPtALzrh5LyBNhWN/UMI2dzXzS0SmmGxKcxb5rFme
2aL9xmk53fM3G82vPkYQixtF8YfZ5uce+JJYd4SlPk4CuOnrJZiCLIVlsjYkKGFh
iMmHzy6J1lmues0GRzgMnSvUpZopwyMT5EGXMWq7fuaxG5DrC7M1P8PAKu1FPt6A
B2L/Lfp0tSqpX5bESQbPSYzY3ry2M7gdCMgnKScQdETTcrEBJUPvEYF2mRIhwCHS
DhvkUtJxufvXHYzefFo3PKvDgDPSzaOWd3qr7t/tAPDFohq9OQBbkGwZBb+pPiy+
nCHbYGW/71umiuDopho7vA100dG/5eNZmcjMYUyyL1hZZohwlZORIY6mQKAyWukx
QhpvWMOq/TEtlTOWB14qTwyr9oqU4ddFyEYZEG6MdWpCfbPGMUdqzTXoeiT5QzjN
Y/6ZCOT3/woYeTiJVhMxaOUiE0S/4k6x+Pxq23EV2fygCWx342Yop0Qcf4EuxbkJ
0oGvBclxzHgHENTHgZSANIXBOSnVuMNZEx3rLscBAcULZUy4pfkKZSMSgVxX2alP
/GCYcbXokvhNQM5bCCGLdBEs6ZlKy8mQaFr+Vr68V5OCGaNfKye/nfGgL75AsM6b
2AvjctKdTMx6TOYxeRCx31l4Gd+Yi3OFB1DQE2TaICfas4gBT/Ieci9BlxIcm0hD
/j22pK7ZLbzQ0qeDZ02GDl1pTpqNNO4EEC2/Uf6Ptl+PhDpf33dZ2odPDfa/IFYV
4ylnKcTyAInRzB9DUWALwx2lfihph9BvqCOtKc5Ds6nGfZQM8BwH5JKG8wWs4tjK
o9SmJ7Zlx7FMdRqdxTL318c778+iL704w5CtBklAHkv1Tr9OhJOHH2/mRmVRRadi
2h90nN2hq8XiqR7HYEcGDbBVmuYKbUujbR5bamoa0KdAsxafzfubCCnLq01BLHG6
WcxlUHY/xoztQF/SwVZ6kTrciW4/0qrBryzgtmkA7RiPKU4pxjn8RxltWiujipq4
6NVfDZkjvR23TeLnJFLf96EvIXzjXRxGOh0N/dvFIPtdnu51nyxRQktxrYgDSQ3B
SfITgbX6uy7MIzyi+F0tDpbvr2Qu4IIZw6fkblI0xkB3dLbnjULXnBTalTZ7nTKb
3ynsa8x7D85pG4MGzgjONXs2bgLDfOtoXU8FC9CbyDOSG+n4tTy3b4/B9E6Ks3RY
pstTNbbPMr8WuGoCLE2ZIr+GHM6uYAivDKFVP0oH3swGfr3NQPhVC88nH3JDOdzT
8S4zqCeV+xmK4ZSijfgEdJcH3Svtb0t0bCuq0ZdgYRgzskq8lzdJBTt0Ddmz7GYr
hZAOB5JRQN35FKtuZszZL0oSeVaJ+5bEtbZo8+mpGJEmAmGVC3Qu7ev+lKrO3Hgz
l0fMJQs4ervPgpm+xUOvdlRAv/zS/DfYnE+unETeHltFHPmhKgVlYkOw0Js+ePOZ
0RvV50OwJAWJbPkfPEvTPc1NZXf/JqMH3frUjxU5nmM8kluxmzG3XUMmhDjrNp42
142AK9xjq16kH0GCldbGi3bshmmaWzeKegtCXI1CdotaV+hCAfpVs5SUIXpHNpeD
wUvyWha0pVr448Fofc01bgKNCUNpWPo5Or2i0hSki7xZGD3N+Obp4U1aXMDpaWhC
/0vTvOt70uCBAdxTSJ71Sws54aHOX9aKkQ+zF1Sa0LKA6IP01UrC948nujE44HNb
TaTHq8xK7ZFt2mXX8CxyHLmv68sEImfESTTAwOFSdvdiHgr6RMly5cdDlKRmohp8
2+RtwS/1BYcVyVTWqz4Ap14Hbg/WzqhhUA9MQtahjznmfFwsl5Ju3aQ81unvZsy5
mIVdx+bwvdoztxfED3LTaPJeNo5hg0+qhaq14peMcb4GHtzUGhI5mQVtXuyOYEt+
feUJ1hFQIe2noMKDKs7ZYoiwhe1jr52082IyJVntG3Rm3eBvHTfeHjUKRAi79QeS
u/Ip7RlOWWos8tmSBTMS+ce5hb6n3S0XaedRey7RjzMjMSRRjKXJiRSfdNjPM0O0
2kEr3dukKnKoOcjHRl+KC2vnWmks2g7e0DtvYqO4PkMXV3/il9Ol3N1FwVz0HFhf
53kWKn94U/Zeh64/frsPWGhNMRC7LL9EiOUl3C6ns0rrdxiFtAEOmW8KHFMMSwbC
EMSrXZwH+jng8HwQtFh/epA2bt3p8l0fwzcACXgOjPSmlC1U366Y+g1pGySYMPaL
UtlVIYbyR9H2WVN9668RO8mAhn94ZrOv+1jtsiPKDsa3Yb5NNQhzwqGA1FCa5Ek0
MnExFqVmAj9yKjE8vJe31qe23XNXNC0oCbOp/pFiPqepvBG15cG4uWcSo9dsvED+
NpQG1fKxfxiFfsZdJeVR5eMUd7hY9AwdczWsX2QEcTbE0MFclzVv0L/kxUmBMU+p
JuQf0EjaInrRS34DAFLTELGH0QJ5icVa9h+eafye86H6ih965ipkrFRxQTTby6KX
4Zb0LH1O7O2fbAbobfqBhkbaRauYmqWu4kexuHMk1/BukQlMWM0y290rRmz3L+0X
D9C1K/eMIoPHMEFbVQk6bI/e3Ld/37s3V/YyhrlyLmD2tVH2AuyCYr4Wwja2yORg
TRH3wQXxm3K+AXoZfIhfRbgBSHzHDPe1uQzkPsxK2k5/8cUSrS38SPi63rIT5ZPh
w3WE/s6W9lizEuYIk3aiA/z+A7Px48vSVFdoNlC15fz2k/TMNugaXA7elaPG0/nz
l8PPJB6Gc2V3hK3FByQknvtGYeofaTF9AgmgkzzQ++AAPf6gqv8NOtmLqaRPXtcP
03CmUPHdwi4w9Uo6WSk0q/8MUfdX3Z3Dr3EKTizETEp0ViVxkaUXZQkq8jodcJ3W
eOnXw2sIzQ7ulT/4PaDHbik7bGH65EztrA15SUf6rhail7hdcsWfrTUWfjpXb0OB
2sxhuyIVYMLhqXlE+zHk4q6TCePpBTTJzw9w/g7cz1/hOIOqAuG7Oz+wuPQiNrLJ
l6NHkaFKeCVrnrCIU9MKqWRnCatrPFHsb/hRTkFWmWt8OJlZzsmBoSKu8Pju+Uuq
8vrCtd2fAPocYDi/eIZ4cMF+Pnut0r4zCK8KL0OZnYGMViuasB1VAEU8P7aJSxdc
+Vx+aaiRcrz3UKrsaf3XtAxaDpTotRFCA2MrmqnoLeh+8a3QNdGLVgW3AJ7TYxDV
SoQGxSTu1OJBbhnn57bn1fSakQGRDuZ4uWX/jqFwtbrgFCKGCc+Q77UXRbgZxm0+
7CEYvUY8Y+Sb0I4QpxAB1Ck21b4MCG1KPcSO7UkG82bJ2YPhMUuPTIhOBCeVBgAg
67EJc+zHWJaSQM3+WLc+P1cnZTSndk52mqkRI9PGE16jvTGNmtm+bQqDKIVOK/Aq
4Ed3whkqKfNDqNhl8NPT3/iHGzlRH8vB6X4BOMcoIspgcaS/HWTlIUF9PV12lTMH
i6tcGfji3b8KOfTkjaQypIQcNQEaO/o3Yj52LbqCCcf/0QGXJl7bRYoEQ8eOwNOJ
6gSkfmuQgioDihpzHTXooK8rKHSB2fM33Ip5y7fburtwd17+gZ+00PdqSBGGeZzV
E6jSSq+xaVKXROOb+Dqj/+AziWb5cBZqxkpqCX/GI0aWBvPpCDcnjveogocHpYP4
Rs601VWVZexFGou6x4724QyhBLy0+5IytlxUkkqkegTvMN71qBBzQbEHENFOCQJ/
pIiHpQ60GUBf7bbsFhXvffBtS25s9C1V6SB74PAvduhXHg/wYDGIdbJc4kGjMaZs
pZez4V1NbrCs1ySoIecSZMeezXZZ75EcGhI9zBQNvHp6HkZ8HZV1ohTem2KA/oxW
9DbE+wGlXMi3wES53tR4t3Bh0Kg1ypdyAaF+IreKoltCRTVeg3xweUaXs+Yq10zt
qiwdm7xQ5JJW8Fo/zYBt8/ZNHkFyIo5RATrLiZ2xDgRzm+EQfE5FwmgAdDqIFAqy
tXMFxh65iBocIYJn94qrgcRaehR2A6Mn9n4TgyVxCF6Z8dEjib8rMy584/nROUF9
DK9m5KKFgJiIxSShELIfe07/JKOEHI88WpWqzghWKDoCtYFVbLT9Es6GVPuk8sHg
FpruJvpfi9aBAUyfIc9SOzFynSQv4W28rTqjI6EF5666whF2Pj6ZByFNxKcRExYs
JvJoLymIRyaN3kBFsefj5xI0kj17w1euuhtHihlDY/VH7TGahcnZsehmR83J+wBr
UhmbLr3dLYjKKHehr7oYWVgZNSrxGzJENNpBazRF5+aRMa4oOwJFIdU07IQrN219
BMU+ipxgvnLsdAK5pWO0MYhiJiikcDrjCXQuaIFEILsiYe45z25qJj/8cZ6F+864
RMdA36OmUK/PIysu1wgk93jC+gImJjcA2bpPuVM5ryHalfJSg5AJ4NMj16TAhBj7
W5ZJOV9jkaemqwNgWyBre+d8hXuRh/T+DdklSBCuH/Y7+jlMi/O3BlX1gyP8Yuw1
9F4ciA0RcZf6aUzbznOxoxS1Btvik50E/oWn4R+fj19LCdzpoHo23z/DpZA9dioA
rhTo2gWaNI9ZoYDcmHsYa0z17z2DvzvwFe31p37dKbqdNbARry6kDucDG4mgJkp+
vUcXBJUnfnUrPq9GxETa8iB9mK6I4/ruluHbquOF/vplGvipqADjPK0mkaNIoZ5t
FRDPlmDxaCDbU+Qq2LA08V/UJqEWk8ZcfWZbMW8/fXF3NV24E8lXJmmalPYCx/ZV
D6aItSH2hduyC8HDwBxFarcdfur/K2OhEwmL5P25z1sPfGtT8xYMtVWBPpISwXLV
ZYEwuWfeJV4ETT7XbtTPYvZLUZ+I9me/SUEmSYQF2VpifGtHf7/XSS427d3TzLr0
NWeyX3/wBnIUj4kzcj7ykbDR7/5S5b9EBi5b5KUCGvKn33rINbvhmu22TkllKV+w
SbUlBEjfYzuXjFMcDUZxOS+RjS7DIFVwy0xcdd6xw1Ddi7T+ruqg2Xz4807bIyXh
g3VnXhHPoep4Bq2KlR0uIIBwSrVxgOhj4RO04E74zM7x3CF+Tq+/6XumKOvSG0cy
SFEqv9L6jyza14gWSFYJzURVxI2Nu5ZB4vZabVL80aMBfkNDBU7Ljob43UVDNX2z
sjAfNVFp7sdecl2kTk2y498D5edDZ+hnjWb48xyHOjQr4GPm3dkQt1hDuIDA42qx
zbGfo+fMFGBP70HU+1jX8JJ2Eg3Ck2GebVnNeLZPvSTSH3njb0MX/7nJieTlYFkS
2u1TSF+vkPG0jq2dZC2G9BoIPziPGHzEtfkVnQBtLEh2Z4lGRwKzrGPVSE8B935o
yzpC7Zm0nhB8Gh+HHjeT0HfuV5CI9JrSTxR/XHmX2R3q2QBtytoyjpR3NjVtmOld
F+Gbq/0fNSD8Qrm6CBhiKmDRfBp93twBN9UDSUNrAZif+vvIVsQx8P3I374gGtqe
mcSdGV6lhdyMQG4ECu5r9n4DtRI/ivciiVOPWn9R4zph5sCFwOWSiFyCyzUew/0I
IDNNEWkOtSEzImiHZhiaZUTX31cCEWqjJZh6QxlwOE0sc37UHx6IUOUP7tdoPlB+
ATsEAkuflf9Y/rbv+RzsUxSwubG+4L0VcvQxumyM1u2byC1A2Lm7g+n+GRFUaHtA
fIYOTksJwZgtYJnaHd/CcrQDs4+/9CSIC8jRGDsKDMEZc3Dnu2zZLqTHUti3awRv
DKu99noNnccxiKMx/NFSgLk7lrfIc+h13m3BQOg84RETBueRPv0PSi9jtrtQHMFE
2DbYwEfqIdgv0IjFpKH5xGMldxEE6IxFlEcdCc3Y/NkEG9pRYzY8OB56/9KgvyN5
AHStrCxEgfU41qWZrnmIMudlWmZvArstdIolFqxNrAIqf9gt9w421+c4/GH1pN13
hu3lzGKxQFtDaksfDV5PyCfP7UGMsWfdpTFwolcvCQYAtdGSmvLTdSqZbKYrCNeR
vj1Es4Zq3+4YOi1gzp00TbVtEStCBYBel9yFtNN3JFMOnRO4GhGrLf53eh3RFb/E
UOWvEhhz9rnQVsZYmFFeSYOg1tYOfPN3kgAgJbF537+Qo/oywGLEQu4ZplHOtAij
9t6qWkyNpCXW/rC3xR9QDfNlHxBv13RJgCFAy5A7EDuTqCBB+O+rD+0ppGc+N/2B
1zZ1cNkuBtJcdLss10yT/PhPG/hd1llF5E1GkQZeSzhQa5RfjGZwtTLhekHcVcCc
BjwH1G+Siz8U9anaA755VZb70gkyv0cZZ3LVOqtzDLBcpK2M7ejWz0qVmBm+oNmN
Or6eyMw+awsLfkP3E3wrG2QiDlxCITNaxwRlgFhP2p9YSuAcI7HsL8A+ThMa9oxA
lELomfzJpWAEZYDRcW6mFVToN9iwgvYkQAZHrzRRtZQ9EEsHmIbN4/KZBX3KMRq8
4CHcV5dhSXDKPFHOdHFV7kiPW90Iiq8+46/fh7HFGJf4hjuVJi3xRMUMZuyAtwJc
lc+r/RovzR9w2S0alhrNi0yRgPUJLSbFLSrPLg/nZJX3AHg/hGh7rU3RTwxNCoiY
U31XjSAUHF26epR6Rg1y3oemGLnVKnfwGaIbDZ8nSRFKGflnSyK2iWA19ENcu4CB
UhBDWatASQflGuBSur6cWZU5SBeAMULiFZj7HRdxvdrPfB3WyNBD+vZ+vKWcR9up
C6Fqg6bzzY/YSnYsVCOKulfcsvNm5BIAaDicaOj6AXtASkrxUem/Ohm4wTRgNa8a
HBzeFt6QvGDkV7mhITVzxylrWHxP4iKHCWpVskJRTdz/2E4aLCMgc6xo4KgfLrda
bBQocSnAdy+a1/cti/Xs7XtGtTZcDyKD5V3h9aAU5DvoW/RCS/bbtYWfBb46o7ns
mxzBeJvXi8ETbgkAqjRm6zxxR3NhcWbBMegkZgQcpHaq+WeU7FzROjpQCYEogOrg
j1EFCYPwhy3/V1CLyiuHiaOnsjPgkHYy5MLK2Seg/p7R8zXvSQik4GOBDhADnSMF
Y75bI6CWcGx4rBTOD5U11aV+LruksJM7+tStxqAzAV/HQ5OC03fwkiLZlI9qRrop
YgvtUhVKWXtQLKPqGUHHNm3i4tr7kHN0NhplJlvEE/L5smAWikdo5BWVEoC0NJ71
wWKsfUtGI1S14CBoBQvb80hViU6zhWHiUIqTKBhlrc0u/mVsT/z0WlzIFaWrheaN
NtPnekl4aeEAcK21vfs+bIG+Qz52wU6QdoVSvJGKbGgdRgCINaeIbWR8cUjjzA47
5EJ+fbrj57b6sVjjvmb4+uJYUt33mH5G/5unHegJl2pHt/zBbJ9AFljILGrHNGHk
7tx9AXHuo0HZ0rHjeN/NhJVmMUpVzHZahIbCLqLoTmUZPU7Pg0s4fYRwk2o7iPIZ
NSnZbEaSyIngh5XaWiiA+WZaF75Bm9y9JZKaqz6YPrl4rzq6rxOovj8uAT4hVB/3
tU7G7c2JCZimIaW/UFSaPUzq1Ur8S7v7iYDoVXMuWxELdiMs1Hwn4/grn46SGFwC
YNqaWrn0B7PzfOO6ZuLlF/3h+yifxXy5Z65R1/LjFeCJwru/vHqwX/NPKJtJYNI9
zzEVki2CojmIlBihQZ82wnEdXoFrihdQL/GxqbLo4e/muFj1whla5u8/BvYMca1c
yfiw0CbiotI1kctIx7n3UpkSxF+tW0Lz1pREgKjQ8p8Jno+U7gEuNKxSKOSOmFou
Jt2G/AYDngUoK2iSh4RPW/JjZKERwaq91K9EjWW3BheRtpRVEoGP4MbE3HdOqGx/
Gj1yCr4cDMsJ3AS8culu0cAfurBeIGrtcDIqISTVeyqVRKiAd+MSpzim97tgBaAI
OR4ZIVMi9/w+BhZlPu+BbiKHb+knwyWUSgnNptnOTNJLEfOMEwWh0lCfLw0oUUcJ
1rgbrQ8WjaXEswoJ5732UJQyWbM9cT0uFCYDEP6kgKIfLlbAQfrIVOUjTAStsJvr
uSJNfliVNExc0zT+7kiYayRfFV/MQbKSIychHdaSff8iECi3eMTVtaHXjVT5cY7Y
CkPqbMwg0YnDMVIaorojleC5FZoYYn4Y97zAlLV7XYvGMffUhJGnNQzzc2HVlTjy
6D5/3TQ5vnQ8o3nrW7QJYlmQvDuPH5em/rJOnnvip+j+7IGODajV6mWBYnv5viMw
PmS1dglXtHg8v/hQjg4N53R5PZZJRfQQC3uopvOzRkjVZIg4MXx9l59NiidEYT5g
GUlNjkNELZjy2QBtLvPee0gAgsKG5yIhrJpGAW8FL2xdejelMEBmqvm5b+m88pQ9
5KpmlcVMHr7wFcmb1s6xYxJuUUYjB9B0aMTT5DqOsIEwfN6jFoPAYU3+6UcBbYw8
yRm1qzuc0UM0prkvQJVmIKScWqfqyzc7lgOpO7pwVc5h2OsKsrIGW+12lb1vGG1n
djhZiTIdr+TdErReGw29L7gbWvAjqCSCfHO9YVJY0onPSkRX3/bElpkVknWA9fkA
nfANF8/8AYx7xe8IluEkOlgSLOWX9NCJUFGuGtsSYRGNYqbYWaAPWDvEkTY2ODa1
9BevQRzphwpEr2I327Wz7/baC+w/3UqrcJHBZKHTkrDuigAGQp/Ng9oTtCnVEtYa
CpMMTaguRbAyye7api1V2aHRMA/biSOINapV40R0JMdHQy4uO4Fst/2J3sJuQNi0
zgE2rIqDmMB8pHalXaua3iClIsqLN2s18eMCGgBflLOwXJD4LfEW5Poy1iP8NZm+
S6It82rj1tOEhpkIHgHPKYekcjHJb470Gf9ygyzruyL75jMYhMP5ekyClhXbrEek
wo8vjE4Mhc3YWRlFDUUMjT1P5Ed0dB1jW0Y/U6qMEW2qYrhCHAl5q4poXflHQjDm
54uxKrC73+YN4wiDYUUjuFwCUTyRgC3AlR7T5E49RhRJ13g8AuvKPj+lY3f8FRkr
zCTZDSu1Bi0PpPZxZLud2nsJ82WbmBIyysdqST0G6uPvmXbrGUWebC5eS/f5kmE1
uNmLrQAs+J+CIP8zy+1I15OalhEVTtbd2CFJmW55AI5wFPv6pz0n88UDyeduyMEH
B0xxIBDFtFVnaTjHTpk/z6va+7p2TLQ8Md0aZB6ydPy/Sce3Q0Oj3uzqkcnb0kxd
Drx/CXvEZoxg12UnnOBFgUghFdT5BZSarJfDKSUwDdXGxQpMjRId2j5IpDqa9zXR
Ibv7DFM+JoMUYHn3mbLRlqFzrs+D+OcU5s6CmsPFPDBYNFA5TjzxbUpnbvJiY48U
+yeq2unIoP5PU9TGF5dkSx4vutBcJBb/N5pwAZq1Y05GWbi5En7+hMfXWn1RGUdw
/1htS6XnVS3mo3xMRISE0JgwXpWNq7GfTjiPLwawez8+x1VFJGlQKqQ0agHImYzJ
5Bf7YosOD9iMDH6vs6zDXVNLdSGbDfGNUcblKvGlqBS0WgyJMj2DV/APUwf4/VH0
uMA//cxMB7TGzwxw8sfDTqkthFKJ/AXd4nupzmmgJpTQ1oesxKE0QeuZ4+KfSOGM
y29eJSQABgEJElnZVSj6FfS625lshYKV0gfbXoNj+cM568BMkalJTwU6q9r2G5DW
SztFTsnF2On59xVGSt8ZPwW3K/Va0/KfUtqqGf+NFmogac9vK6wZAO4XK3RTACkR
gzWULAlB9ryTwThQBpqgqAYFLWodqYAY/UlEteU8jJBtpB+j/QsJbZ7g9WS+YkT4
HnmSI4Wc8cQEY0LeW2NQ7M5phNwpDfhgdevFdQPwvXv0awK98WZILYNW5U7zQi94
OrBhqykl4QzfqSBGKhfu4k5RPlxn7csH4f+MFXMTBViZRxrgY2LcD9HK0RZNScsR
ub8cMSYx212kZo9Zz50h5yBYyHctowvCtRFwbqpszZyWmS9FjvWXORzp/3FHcOOL
Jx203heUObJf1utf/AZESpH0cLgR26a9ILKUp6tnVjPHsC/XPnIzi0e0/k9IjY9U
Ru9d7MqIM9aQg/QcUNgZO9YnVwmR+ABEBTH0iuuH1Piq9H/yRFOFCMYmIWtaWEvc
nzVf0GVtAH/AKAFRxlMXp/a3IeLQpUrmDHvvShiqjkj9+OzBnwXCVR3VgpGlrH2p
TFi2nD5KwQsO1O/GyAkvWtCYoY6eH40Vh/iYN9/12GMLHccFtJrTY9/vfT8RRUjR
RY2hqYzkvtyhzxMgS8/ry2DoZ18sY5JBnSnAKPr4k3Cin00ulkSC/0jp4iksD9xd
xhd1uXeCYXMhIuwMCnVYnCmFNlZ3ivlrN9GCcvWghCaaGyo1T/H33P9TUx6Wh6oX
VVDov7YY0dyIjLjyzOyRIKWm2ilb3G8UHfboweeDKLSehUM8Z41C5Mi+QqGY7svr
tmxbsmM27Ivw61k8qQgymn3fMxxRaK3sYTlLwIlJcgbU4/BZez9/tIDZ3QsExxDY
R9r4ZmcGEbA90CJUjp4NfP2fciDosqrv5eN6rKS2OAVMi93xwebqMxLay3B5Rt2a
43NNjyrgUKzKihyiVXAVdyA5+fThjefnVu2R7VFxikKmvTcmZfXaX2g5ZfzjF6b/
+h6WZR7OV9ypJLAhPG+cTgWZc3hZk8J7USI4WQTxUYkl5jN4/ofCM+cMi7D76lWx
hYX9Byd9zkf2AzKW75gue/b85pmNeA6m3TQheRUSndWD6ktLVkKbdV6mKpBE7j3C
/cOh4ekKKRiEDov42fvoufOifaRilKVm7x70KTIAUtYpNPI8HjXhIol2ggd+lctB
Crn2nVBJcNAdl4QV39r1kf2CzI6dqeF9Z3hAkW0l+ce30ONwk7+PclIgVXumXSQy
DGo0VRVfiq8Oz73y33DJQ4TUR3jfapWSxdD7oBdSO1CszJddLFfPxfCYIFHrXWSl
Hrc0p9XycZbq7RzTEAMZiUWmH0NiL/l1E7kNlY3MFkq1Z5YIAFj/vCzFIrviFU2p
bNoXBesGfuX1N4san9JYEHzbnM4TZNm2IWyPbaohOkmu59myVMcsc0WPwKhNvI46
TtsT9q1Qpjljo1UO/HD/MwFQjQHqon27gBv5RVuQFEpFs7wjKoT7Jr3UDOCgfERG
0Strig4ZFIQttSGoIjIPmKAAoK5DGfZj1MxVAFa/LRD0dR7TjNVPayU2RUGMsY5a
WXZ499zRLkRaDupQe1tpy0cpA5/bM+4vISF8zidApi4wu1ROSVnlR4JyT4PXWPyW
zlb8kwYgr4HHNr998/qNQ/7l98bkuhb9qxuFIGWSBOkqDuFeI6WH/ywzdAJbYj/G
9nDrzxLByx89cpe259yZZ8EB3H3OzQGbtdjARfx4I1daZUs+WMGeFn3RP12rzgAL
Mu9UCI96BsCvwE+LHgt2e9CN+vGdnjFaD+iOZzdCTiwIbYMabdSBhyHzJLzjPn5a
uBTvRAuzFYzLPkQVDZHVzFQYymtQDsj5nruidoZIrU+l/c6TZfiaNim+8rLPYi5z
NpaMfEtZNYqGUkkZtICXYBYuQBbuCcgZ9tRhkYG0HF8wu8doUTAjk0/YUinXi48p
cfoHDhGJzRGpeQTUSToEK1n7xjsAUjSy9NTjX5zne7Ar05Vhu+0QI/ZvctMPFBrp
Pt89oWvv1nV5FLEU+nr/RH/tJfdMR6pGfXGDjJAXAQBua6lY0jO4N5hrBj5IrS/R
9Y+OkD/aUD3THw+0WZ3F46wwuZHhKNsdkcF1qyhOXBvyRifeOTCm2cuuFdMVtCt9
RiVQCFIOUnogA0ZgTIiCm/sI2G1yoi1IFAJ3/cMh/xz7KEhwAaaxDXwThh+c9mNQ
b1Wk/NGqBiTz9FEvjbqxGgWwerKdevY35pZTo2hdzMd8ORBriyM/d5NGAUvlH0dX
Wpku9pCvPWlkAq+XFw2JLihnjvf/ef+r9z5skkigTUkqZrrRJyB1apA0YKPyGvFJ
bP4Mm5vE1pN7xefh6tzqm5nnXbZWexu0tvOaYV9grV/wWgEcjiuEmvXdcFPiNSu3
45x04Y2ctZjW2+YUfIZfbnLSXnG+eHBPQlH4w42dT1Oi8PlkGOTSflRHSVysYWpZ
io84cRCTefv/kmSnKeViurlgXHxiZOORWdeVbryqkH2C4nl5Xd3KxAh5QqEUP7pv
GqMAnTGeMsheaUFiXRHCVmzkI1lOcrUCryKiVCOGnIQ+x8MAnC2Gd0W5wO7a6bDw
x90xzfbPgd9qZrxrY9dJzKkBuZpcx0EalAtT/5CbwKTLu6xE+rAkL7BAhznONNlG
ewoRLGTk2EOqmUKOg5uDHfk4K79K4fsqp/jqd7yZywwZxHDzLrpAUqkzJFg0PWWJ
2Kjs/X5JfhV92jEB4qr16umpdYsgyZ7XMkcK2ZA9hFZs0e60wlHO21++ixgKNASh
eJYD71FowVasHMFrxGlZlVtKsV4LDihe1MU5M65rXhA1mLyRLrp65FLkVzJMpzlB
B1GfeWwEdJghHf23rLDdKvbT1c7ehE5KKy/n96DE6UTENncoVNs/d+4N4YrUMDeH
BJ3PqEF3ihS0SOt9aOCJ4n4Xq2Tjr/6Z8pObs0zhKom1k/Ou1iMc+qIuJtTUGuuS
Ar1HAWcwCFUVtNmYgwOLD27tkzMYXNIgbFn/EkxxkxC+Yf7mZpSdliqcddSYGoz4
S/7UPfEKLamg2oPF7AwiA4IC24Ye+IK63WbUwlxHhBReTtB0w9DH423pW8mrLvwO
EoRurdNFzGWzZkItJuboP7WVQbj1e2GZcKnRxynHOxlTZGXffHO2MIbGq2Z5Lfvg
ESqvBn5G/54QHlbE5uX55KZt9rWptazH5W5++wpghBYTu+DiJNJkaIJc1IQV6r5j
9FKsnO3TKGUmWt1pDLXI0606cSFqCHSXEikfsjel1u3e1wOU7PuekLrObWPcAws4
VrfKseV2Fd4GDwllo7gn1TZ+CJAKS8Y9EeIOOZKsllwdL1MM5Szc3ePr+zApgidS
ylwBYgOcYsBK0MqpmJNQDpMzoTBJXmV4WqKqZdrPAACU8afFu/wm6kJ9macxrJPr
ImS88OzC0JF8eeEQlkLi4LyhyB6L6+/llleV2/UAyPAphuheodlgmN4lNa5t5jWb
bEbjSU6Y4A8JUeTFZn5HoRJl8fTZnY86sI6lNwk/ZRoCGAM5f1fr2arvqQyQDSwD
KcinWMrET9oGu0pDrJsvVNCgmKnRUzuFjrh2+lElqthNDlmFWT1MNSYOLcNCxXV2
0d+lUiT8arfdRKE1BBG+v2GowzZddk4tVzc2+AJxXS+Cth5NVo+Vz+941QsTeXrZ
w6JdLo+ymm3gdXY1ldKr3ja0nUBzXaVwJhtdqTvB6UhR2t5NY18wQjNaVJnSDUCM
NBw8lNSTlHPByuyA0vMiLFdHPRNNneVRDrvOEKeU/0QBySL/cF/58C3yBEdo0PyW
TjNouGgmCPMAT9Ym/qABgI4xHnbytWKyiP11WUW7LoOtSwonjz+PMowfsCbCgjLi
ALyXD2V9lVQgOWXy3JJ4m2uj8HyTsg7K9jqcBLi/83JQuJTErlxAiWa9ezfdNYpK
J4iURwuVGzNT11iKbuLRybciOlZ7tePmlXBrXRDqmAMTO/ROj3ML5yZZlDixYh0q
y4640FCMaImhd1KNcriF+GV27bk7rOuVUBqidZ2TvTsZ04QoFK3hMLTi5jZdCa0e
k8C/CUZtpgdlhgyHAiNu2titfsWtWT0/IjOH5F9Y862yV4Be7Dd07e39okTTT3r0
J1lJw41G5RociTQngyin35K5Q70aZ0JZkWIQVgCrSE1EYeHNe+9IjFZTEXbGeg0d
Sc6zZjn0LqJzQwxtihTBmcgq7nA1v0KrkXR/Z70YrRsHwpysNYld1AL3h7ONvdF5
laNQ439vUt0NR5aOSAHwG4MTspxTFdVc812rFi70Hlgc6bhfIXmN7DC5Hq+lCDCV
CRpFV6KS6pB7CxKWhQpcRyVoOUgSZfzDth0hfoIe+H/fMoeOzSIXMKuz8CyOkWEB
trrImO2wHyUsc4mh07ujQEnQflH9dx5ltMETPJQEVtrqjvAP7rWfSt71yCzctW6W
ACd/k3dU4vRmRj1OHKL9m8yqYbMMSGYc6WKgSLnnZoLCBfeEqnz+yzcAXmXhQroe
9Xt1jUShKTHVwP/iwFkIo/aHNzLwbGaI0237OgbFCRbBSjWDnzZe9nCBHEj4LAPz
C4oZklDpPZRBLneq2TdWkiiy/NmfViRwGK2D3ZeIgX874dOOxWoaPyelG3xYZFuG
+dG9Z3mFMuyENn62ZrwYKZwTqIkOiA0RoOvObkYwxugmiCZr9kFCPJD/tD/kScbn
H/ICzlwZ4BI4oC/uBUJME115XQL1RC1WwMq8FraHmZNUIDZyCySzsYU9p2p+qh2O
8Ot1CQsMyMRAFvRsnI0I2ardwKWs4k3DCgAy9tL5ZZPtT+YQsPY6hAu9H2h+WY1P
UJldhcnnJT0WUvPbaOwIfHMJ5mY0gMyFsEVnEFBGd7FFx24faPYylyI4kpIEI6Cx
GJb8nNHHOUPadUtCO0elY/Gd/7U0/wBSvFjnKrLc7EIOa3p159PDxW3tAfErBNJG
tsMnQ2PGoIW8joQfzjlhAYMgqbEn4fS3vB/TXG9HFHO86ob1GvQ7g6bQhjYRm3Zm
fzVprTKCNRbRP83+7z1UnmMj0lSG3vqHn+OadVwQdg1tmpnAp4AwEQUuLDX0yYx+
r2Azz3KDgWZ9S8oYJbAsm8cN9becRsvIHye/5nx4mmthrHPZfNaAG/aMdVMynCf4
PvvF5yX/3lgDTO3rWpuoXykwRQMMyc3abpayn1UyZJAzM9h5oh/BdugzPdo9zrGo
xSa3Wcao4DZUw56dHAqTChyGk/fAY4hXknNgrGJIf0LMzCr4kxiSzVOqx+XFv3Fb
T6hHr0/ISsfKPYmMVLmihuuqIe7wW+7Pd17bp/ToXSIdA6vi2FyKB+IZEdvZgUhE
ixjPE9HYYoj7N23oolYji4s8ZI6Q89oT3MPTlcMenDobeFXUkGiZ0NKgliEeGLzf
XRnKQdGSi2RZtGJoeoBzxJ9tpify0v9yRo9dm/9ekPJX/X3vusveugQJ1ZfkyW3N
V7ZaB8DkObimtYnEn7axK2Acox2gwEMpNQ5MrRLj6kx0+RHEIbhd1fiSsmVOk3I3
1hAlsrC++vFCUzyp/r3XEiFkkdO4wqRUkTQGWp8EI7pgaN+FKj8IefPkwk8gvRik
UcCdTz4M3bGTeJEoeEH+nFr/NZIcPZUCnhvBQV4a6ZFcpMLAAGUnS1H7ms4a2VRn
GKPleR18pvRkQrSDYnNcTYBb1bCri2yN2+3SlD96ETTlmp4yfn3vXPM4S4ypnhsc
B9TP/aUPSZ+2rPaLwqqnVPWtXI12dvQEvuP847wk2dYkG//QrUznrUd3nqVf98kt
3xCA/47MeIAbqPDkPXRX3oxjLdUhRfPaAXS4jm0rvJ/sAjqB/HBrp4NkDK6/e2Ct
EIMY5AuGnW6CuVdUHfzwyDfNtoOk14kID1T08YfpXawWTL4wI/JOAWZpscWSnWDX
BbzJ5WxbAqTDizJWOpZPANH5dEkH2JYAT19Eed62bANMqRrjnle+dH1rYxSp5uIU
B77d5qs9SsTPhkTWAvuVc+A7/wOZBY4c+mvA7wjiT1OXlC2lDf5D+hbeNK5M9867
ws//BL/YAgHMMS4HB/saTpb8izdEQy+wAEWsJH9bBxPJuBTmjSSvmq76VQEEdUPm
hPOmuKIdYeCYUC287YRsvkXSVLagkg5Ynw5Gq8Me67sdiKL7R+jhU5rt5xQ7U89v
fOK3uo1yZUmql7DDTXKYPPdK7jUomuSKmorjM+jXQLfD4B6e2bew2rIuo06aCOYB
KvUIPDVK9tquleBDk5Q7QAJu//Oh7XTKPXQqczKhnzEqB1lHXy/Hix91p61bG74a
qsql3EK60G/imd96O4KKxgWObnpu6f+ALHBXkanuFEscqn3NmlzCOessnMCf6npx
u46U8g5+FXgIuy4B2toQvwGe7Rp6+k/ET8hZgrj+kHMcX2hsq8sMz2LpUU3SGU6b
ngp6kw/yPYvSsv2DSaAPWLY2NMCUfpHWJUCRhW/zm0AnYUUpYjD0cHhY/nviHdzU
omN24oSOS0xoZ6RxCycJl1fV2MRY7iVY/jYCfl5Zw/l8DLyEGmpB3WvtEuRFVjVV
HLxbr6kU39BNRKBfcBrMSMFSysl4YNvoypmi0MIR8c5fX2NC25nrTKSf8clyZM+3
Gw589I8tnwxcwtVlPjLpq/F8VMLT4BalrimgOa/nZWitQntgJP+9yCt2I/BtGSec
MKpjumPz7UUA/FJPvvGJ9lETlfT8Anz3iI46qSjjm7g7VOsub7qk+zlL3KtVQlC9
BjlAPeGy/jaGkqxVLmsjJBlBJ3yRknBcRbNp0ZYSeub0+V9BnZC0k9iEezez3nd+
bzC6LYnWIkUqjCHZ0AcyXmwsexE9grw6UwJVvrsEU9VDX7Pc3CHoFLJU/5e6hkzv
wgW9jpO/KPp0qgvIpqTJbPqMcPoaJt3wVNe7jDIy65kLB6bjQo/FJ089Iz6LeB6r
jmfVuEEhUgX+JrZUgDEGrIZotmvSsJIv18F7FBBYEKlErugSYna10y9jd62HWC0P
5Wt7+xlt+h6B0xvzY9n2+XV/l6aJE04bzI+YHoMh09SIF4JQfrLFFJPwG9bBStW2
zY8lDoWFkSwdGnKfuKkCaO+bEMAAH+bRq02j46mb6AskT4IABI5mEPsXrxdnSFYY
8IYukGwiMFk2AP1oufBnOsblSs9zCZGj+dgFRbkKEcYNK9Yf8CXxrrd6S+HmgTY6
H224XGCrD11HZPyMoaQg5M9eCeSNgFZt70ln5mXNmDBEs4S3UI9JBEVEBq9D1kOf
oYl3MmtOCWpDR0Wuf3MKVG+i61NoW3ys3TDygPSlYFifinkjlg4gP/VM5BK7O6Fh
E/VwfTelF8W2+yzpk+XqVpgOlFaXHas8T8iRht2QNkKzjbrM94U9ggF7Dqjd/2/2
Lp/dFwnQH95BDLFNT3fulcU5LyyyBYTTyFbuaJdiU92J9E1xfw+jCL0IYldAG7LN
Y831XksECxoGNAUZWGgG/CkIqMQB+JfwL6f8r4sFIShAORqeQ/d9NctiPsjzPg3b
skVb82iTiinNzdoIauLeJMum1ZcB4FMA6wSyttD5CyymWm2B/Sik+wSSDQyN9eOb
wIMLiTFGB7ravngpxaQxou+Fh1crnQpbiQx0V2zpiDurttmI3RFD1zqYmTW41ILI
Z/A4VeTmoTHuIzufXCBa5AD3i6d80QQlDD4waDwORE+/IRMptDluSJpUDr46jztA
5bcy7BLyzYQNR8InNMwoyfFENZjTbS/6QZy1pi8mmAC/nmYi/4RiDjrI9KRkqPJi
Gvdl4Tzc+KXyMxvFtF4gcn/IT6lffI+dO4QjjhdDTIj4uKakRXYF7We/JSVqZ9Uv
Ow3/usNRj1xOW+Wg06PzuB7yTLaIIB5p0VqB5ZrPS4H+3Y4HpLT5zjRvbQbYZ4Vk
k4QsfPICx0ygF77WD2sD7jCtY2wR4rY1LsO3NjQPsKy8kV7xflEbge2Htt69qzY3
eURurXHtluSOj/HCtqsC2+vMZUJsFma82rqemOlkryJtj5bjP01aZnrv++t7558P
7P25UgUWQ7ciUHqO10KT9Iz8oV5U1sIxxZumdLYjDCAYbhA2wZjiC/hTY8JEWMhu
ymGRyHs0/IQbO8mFDlABcN+riguKBiwbOdKI2cv61wYPH6ADofhsCTHSXZ9GNhl6
+7aVzFyjhSNOmf35gFqnlP5E/OvJw3ZSlgpdEAuNvlcmNvdW2wR6Jww8G8LxrQVL
leLllxLguKLSMqutxdYrX3aXaRTwamufqOscafCWysIk7pvNlgEzeluURKSa7BBf
VW//Ca3QqhcWT/Cp3GDqqr9j7b8cTpkCOubAopjptR4QacIDidhc3jknpnE4VEGz
umJkBX74eEnc+wcbay1Jaus15aUSVjFVrX00aIISEhdNm+PHsE3FMMROATGJPDLB
DxENIyMCIZRyFgNAnKKFTjnAr2ieb75AtENHC4GoGV5kJxQak7/TDSDQBkSZ+VGK
jEXUL7I768Hiwsp3Xkn0KKtbusbsaX+nQ4gQ/22y5yo1esg7v1TbjgyyYn4aTs69
2Dc6euzisXp/A9Sz5AV6FOGPV2nSBBOm9Wqw1qXy6trIZkON0TYIjgtY5NPZ5K8z
RhTETD2Ogm8PXIsA/SsIb+dhqQwpVq7N/rklhh4aMnb0Ez3hvIakBbom4xibcmDw
IQwDoNaEhcVFsUDPuwSqf8dkWGffx+l5zlj9I7Ck4yJOF9JSDqPDE4bGd/qHZxdB
5TyYXuk2xlbqsbtiN84bw+yeC/izg6XnE0n/kjYhoZrOeDd5MKWLSKNkCc3LPa4s
FmKCtLp1cmLaK49TrFhcSIvBEymc5U4znssWx2dYlSYUDbfA1UpJ9NZ4uJSC6CVN
/3tF+JHYa9ZigM9Cp8RvPQObXpKHTlJW2hvUNVYKxl7Kuo9wDmIaGzXVQ08zEhXS
8XdUW37rMC40hBcHSvnf5dz6CjNRSzu3GT1Rod45mx//4+hZzOT1HaV29F2JvXhl
uORLMB+PkbEZtw1T5jiHOTGsREeWHxHNA9eVgzxGeMCQ5eeF9uacvK/I3AEbPgnu
PNV1bBixqSxo55dfVrW2NUOdPhB4GyM6rKWDtlkq6Qohaca3Z70yIr450z8L4hNQ
yF2SpSag3u/T06n9kU2G1f+JaR7VPDtmlJvocTfn8vLHPydQvngVeqlMl/dXciQI
EqUqRlQe6feh5dF3Wn0iN8OLTqxHbUEoLDUYICIZHDREUusFjEXTpLFUNxWQNrPQ
fjEsXo1hUgU3Pd9v2ior6+UH80Y46wEmSiPTwRYBiV6V6gdWzSb82i1weK3MLCiU
h48/GHCK4tOVtISl8JdLoL/APr6r5AmqtyL4qb0tjSAgrdJzyoJ6P2f2FyMKbUA3
XbUQGGhiqeDOF3kItuywKDxpe65/ozrTl14i/m9PGAzPCUXCP2yDegdPa9ejNfKO
z0+ihQjvce3hQFCI89TPwYEIvShMNxt6BozJnfof85kHNu6tlg1cxFX0r2qxLUNf
zfPuiv7gTLcdlaCk5dCv3c8waRyjbUwc2Dp7zNu3yxuB6/ZFHEsp+GO2Lb0vzxhP
iWjXglzZK4Feliz5pz/U/apCTPk3drl4IRWGUy18Vu2VRB7rqsToyQezH8zU19oT
ilng4AYa0VU2V42OJ+LTDguHMuIaeRDX+mLGXgZki8GORM26VCp5twMtjw1sjMoK
+O8zE0yla3Il1oXKlY+iYoT1Bo9moTNX4MHsfTibbTIUM5OXqY0oKRZayDf6ZBYT
o2XPRnkgUcVmqNjNREGBKFT9PepOXkjs3tX5UYeV8YAUcnRcyKLJ4HZTEOXchyEO
ohXwWCxvYcYKH3Dw4o6JjwkV0BL/ygwAifNS7E7Wmj1s0L14J3FRXvUcIye1GTzS
QeIgkdF73qp6XI+VOmOkAsaMzL5x1mbqRAGruUENm9QpGYLVm+5reLMW6YUjv/K7
h3CH8aKWRbvroyqO3vBxnSbAPIerfPvNdB90o5AfuzpYMa1mqIGU63Oj3Pb1teei
7TsV533NQZ2Co0FIEXUSoveHtTeQKi42VmDexda5y4GFfubejP3mtDDKYGhkIbOm
tjcCVytHJCyp+zeDHy373ZLO3saxGmdeC5Qvs/4FhZRoHPgsGEvXCeD0ASrbiano
9QplDg7qm0gshaz5NEmD7uF3NDlXXL+4ugQJ7z/zngZOmf6Qrn9bgHIghh/dbajK
DXyfld7F3Cj35lXcJDAtMKOCMV5LjeXL4I+j6QxeraGh29r71CHshH9yA7XWne1e
iWx/fcdBhwJyuM37D1SbZCvGfbeEx58X9X+1Nx7KbqTbFyfRqrg0fBu1mSOSxka8
zj0Jt9hroMSHLQtCEvtjqmOzQusJKJw7G3+J+oqONdM8tdYcwQ5UC0A8Bv8+lr85
xnfOWkaL34Q8zNyUK3dxjLQemRK9LPaUeW5ZLsw0jaYuRmti+HP9KmY33kEzl/8g
W3GOhnLOZ0EZ0XUpHRLEwn7Ltpv3xYR91RYuVs9Z/UlQshoCgyF/v9kWv6cUnQF9
zHqAzRT8KzD/wsKh/AQIMksRxG6l0XroUkJt2RrpLefvgnHfEE9WxouabBkDuK8Y
8ZTFI5ekdu8PYo4TE6MMyo7vWtEMqwk0MIiw73VF9knz1txKPdYaGx2sm8yEB3It
AhvI8roDbZN5O0NOC39dOZnZ5NHinJvfLnroa6NQmWebYolQi11OY7WVTuC9q0iw
btd01N5fH91aht5r4qDCjhOsptqieodQ4fh0em+DWm4mL0FiIngRQnOJJh1jy+tZ
1SHCKd9iselJKs70zmTye31e1Sa8FHLBL9zmr8H9RhkycqA0Yh9DMFKF+XEkHZwx
uBpGAmx20bV83Bk6AswRGaizW//iHi4pbgyytvR5ukPrWA2B1+Cg28kJEDBjgode
dMBgI8aRNgRrcuQnzjxS0Yno+Kj+pHtN40zU6Zk3aGpgqTRpvf5b5wV/KsdBf1PB
hIZRwHYmiD3P/qiCInf12eJEacpnvHPAsaLpCuHqK3a01Y5UYoVsuN6L5GNtEMoS
jENbyHo3gg/A97ELt2j4NuofZfvXSkVxrSWOx1AqDlm5SilVpCrc9F+dgYk2QNoe
a1quQC0pQdW2m0iAfda3i/eAPUxFmJ8tweWQsXGl4f+/Uqq1tIjruhDwBlsjSlZh
/0dMshltT7DjD9XYiN/yA3bGwVMptp3J4gQdZTN/4RC0t1Qq5ZDTx6JG3baYmgqi
JCqMC7wZhusm6w7NlJpvXQytnn+J5GSR1tHi7Ly9/XLTWgyNAJFtL1xkW0Szhylh
666aStCHI6EuT6xOM+diysOn8Kldk5TaDW/hPqe9BoNVloM34uCZC9nbDYds2XZv
hPuUp5BxCS7joqjbPfzR2M2QV/TY+E0/d8duynupdCvdg9QfrqCAAoRiS4hGD2gI
DqcHNgyI6EyIbMGTHtYW28TAnpQ0HBo9hfzxUm51iFZT4kyOe+AoGU0gKjy9qjFG
XmZt4W2il9O0e+BvxIVLF6toL/gwYnXkcfzoslYRLfbo4wlrfs96hq0iw4SQDdg7
zbrfYC1GtecGntpVjaERF5O8pSsONGngT+8Zq1SlGYpZB1yVCnIYolHPA/IktRFL
VTiHYdNkDh3DrGY4Q4OuZ+xxWW8mSOxGn+aprCGHvJ5SsuGqDYTCoJJ563VmMm9x
MT9gTXgAXCgYfh1G5ahJKksKRQwXCK8EUI4vDzXKiuiV+3KnwSVmWbrZDqJL2ZmP
NJATSOGu5SOsubrHUfoVrw9KcivqnHtqNsY0xz3id0IX9ZNoxvKLy1LB37EicDmc
MHKLV7s8lsyqnBLzYrDcWTK+8+nuseP/rkIFXDoEbj6H7L1P7s2IwE7n4SZhBVad
LOC6HZLExpqNcLS5lnsWBA2ptLxY7GnXaFWWCZqd4Fq28npYgyd1fFheezzJURzw
6ZnLJzaDUOGmkKW7ykPJwfSezlgrvPpQbxs+3oqUOeiHeLuecR+dQ2b/rmsz49D7
w7z0vGarvT7N5rLfFxpPNXXvs0LteF4s2lEMlququOYqN4zYJVOZqF8fBFC8Azbw
Fbq5pZVSTO8mkRdZOlNF9SUYiQ0dBZHF9vYgnBQ4SCr5Jzw9SArA19TI2A8J7mME
vtq55PCTkkBSFgDELFN3LFplSpcw/7j+I4INdHFcrbZQkJyitNWPfRvz/vRYGD14
CxQ/oWnPvETlpgkYjhWR+lDdiOk93UHAuaSp2fB14ajFQRh1UOIYvVeJu/lYkwpR
QOGKiLSKpWit6/EQMpJvi07z9QKqV2FGFvl8AlSw8myzei8E/ncW8RpFaxiPo8cV
RZh2gETzJ4FWy7C0mrueJjoTbJlBvVpA8vuIzWst90PlJBF5TGCZlHWH0GVN4qUf
FQqShObevnF5wlwR2aaaXF6+k8zKFTICBjDgQ282LV6mhnkrRyX1bNuWPz+EAoQZ
vHTzFmdgrpmVExwTLHlTUey2skzdujE2TmwIxs/1qHpoYSmFbhmR2TkJPjol9SGL
9dVlKm7R4j1LSusLfHcU0mzV5UMwTU5BznQPfL/+ndQ1iS53udfKuIuBm22jmLPb
WdHnDrFELRCR5oj1QlIKJ8yI/bPXoY2HA4KXTKqp/tqX0iP9X+VpYXz8Y7OOmz7o
m1y6qTZ5PEXfPxblpp4IR1Yq08PtRx0nNwUaWZmbQyyy8qXoOGQWpb9iut6Cytwt
XT2notOdLAKfaDCfPxJAR7OnPJkFTEfKDtvGSDrA1z+OsvCqTWtYZyXnRIk8w6kP
ZxQXab/jEVctYckUPaq+p8GAruXkk3TMjtV7ZtyzzYbvwMMBWUBs7Z22kgJtw23b
iGJ4VA9tG9aI6yduwamrKnDXdd25mN2l+kyV0g+UZuKTuBapEOR5lGsoTKbKm82t
QVsWPMoy8yYqSsswq3Wp4iR6barAco4FwUrwzkTlIqlEGXtGtV4RlnuAKxDNHfGh
slEKRgUIVc2EgN9g5BSjonTHe+QuO3xyo/wKg8T6rmKlqnbzTKekXWLKsbt7IdGk
nxMIC3L2Tv7kE3p7o6lYPBFe5gumHd2sPZw9dTowMK7fprbqc2QI+3GV2uxBwX5m
1sc2OKE6ansPKP+sPfbCPM6BsXBcinquO6ekdUyYU3Anxyzc8OgOasWzuhsU2Urs
LOub7B+IAgEOHnQU7ZlRzWx0dsIFvg95vKsqt8mPPxfcV5XC1Jif4mi3wdOHQTCk
OJtFD1rg1jHva5BGLjBxsvO+H93tur3EAAnMAk7l8coooUpatz8jdXexE/cCIsqP
36ZdLieoeXuBWN+resRw5FxJlSsYlNLtY1TW/XR/WehBxAoS6yWcLkNyGcgxOeMR
NQGU13Qp4oYFTNAXxt/U+QllODkY+OTyhwgBFHoG+RJR+JnBwYreHeCT0YzNrgr1
FMNkmUcou4QnTlSfDZUOVP6buxTUeGN2k87CfdRD56ZkeB+A1nRYvIElAQIJO0Fj
R8lEn982TXx2AX/1309+fJhwxsbyhz5qHqmzSzinW4qvCwp+E80U3FYxH9QZW/wC
HXMwdSWfQ1yoadXagEanqHnGRuV/eF/NfeY8P79ugvQJHfykPoiVR58NiUdCvCHq
RGI8zWTsbR7JjuAvl1Ie1Jya1pZPCZjOXskXMx5POPb7odjMGssSr/PmM7MvG0Aw
CGPrYuaxKn1nRwG+HoN604uUNa/7rA3IICcZeavXFBTL4Vr7c/5g3yn3z0PtCWhP
pj3bsQ37TVGJakW6cNhH68zQT+VG8mw62DUtD7DiNYLQiuOxEO4nktt9MBe++Puy
533fikq6v0oKkku2Y5UvK2ZXiM1RHBcIbNNCfaR0E0cwAuqL+jHG2gCN16xcgH+r
zNe6Hjhv+npSvWDyZcOzOzZW2EgUqk971cJQWv1SamGhpk08lr2oUbKHHAJMZIM2
yfqJuj8rNYkbIh3Ddfu0lJo59HoaQ4lOTkhqSePaduASSgACZFuZ6OiVWb0KyvNh
/TVAUsR2oDkyr9PHlg1DzBk6T1tcLf6z1uxKTHZALZs5SRDGEU/rVg8HI6lLj5Mv
mFyHkcxDz4j5RfsWReO6ZiOdc8SGbs92ezGGMsxSIBxs6LTB0FmFwLdv/r5n5ZED
ZYjw+/ZKXQTGFDOLMm5QJ8U5FVQ9l23ZjRMVdfopBMcrwSSCHb04sG8/z8tAGtmY
4yaiCyMc9daZI68oHOofMAWF9rthubkMCWU2nx6PthGHh+A/lfqfMDaNO9Z7nlW5
XUQZCql6KA8ferw/CdvmJfHWE6pf7cFAam1dnypDRaC6erF3wwM6GtbDTOs5mc0J
L4g58gzSU7rDR75CXPwl+oNURjxrbcvsq7Us7SZ9Qp4zI1Dgh9BaiYXiiOIkZ94Y
DdaFxav/8ibbDytpZBpytkHb019fn6DVqeOl86c0oRF/K5PC/59EU9YuCkPBP+8m
UemEPB/jRpRfAm4vL4qo4efJtRgpbx042ZH52U/lA861vjPSzEklsaoUfI4awLxq
mfuVuqJFiFFKp5BvxXUzuA+2AdpsrlydHNeMtL94QtL1U2XFVHl/B/ExuibfQRuv
voCpNfowdMB/2+3fHAoBtuWT3rvE25wFnrLUR/cx9gkYh2U4C6a8gcxP506nIfEl
QLOdZjRuQaOm5Pr2usP2EXx8/1cg/pvoFoHPmIYBd1oiwb+g1/YdKGidCguymXi+
djNnDjXx0WBUfdb5wsfxfw1ocscnRsrpyN5lU7kWKrQGueqogMX5xw/cC6tfYWV+
xel/n2S+ivgKBvFKRKJS5x9Ota4axV1yGiEsRh+ljrUuwxNau1mn81Rx2qpvGVc5
ME8i2c/DvGQgpiVmkLUIXbaFoQhHe5SqYKuHgw3fhy7M4GqqqLFwFtma6X8sViFu
yM2iCzDMy8MDCKj6A9Ewcx63+TeqXhHz1H5pYgpAW0dChhW9s9KrhRUySAFew3tF
7MOsNVnMY8k8UzSiaPnWBe6800LW6j+T+ph5XNn97y+TtD0FSh5YmZ3f2ScxJ/Ey
+Y/ZfLzWITTDRw5QwpI4wqEsZ0E6HqWGhjf9rOERAhM3+lLH//4PHnGtUbkDQgRI
L1RWF2Fc3bQVYLSVbj+eRVmr+wWS2NZZjCQBW+wjbCMONy44EosxvsseyGCbhdyD
yoF980MisPdJazEPQO73LeIBpRWMowW4EHxw9+N+GCXSstDzORg+NG6Kzavij/nl
7y/TknyS3PhZ7Q04sqDDY7GSJBbMTJTCGYh2pIr9gKiW2fc3o6t6npfStJqy71yb
pH+8XX8zGa8tMG1woVk+iZTQ2n6UhHOSF29waM84DSpeZOlWHaX2ZhZy+ZDEBrzs
Po7NeCj2IgaUuZsmJ0zEdRR8RITFZGn7+SRF3mg8InbOzN0GUo6b0VBlmXBu4AW8
oxL6z3t59G1orj55rDQgl0ytAW3iCNWOYrqA6HO9XcNOg1E/7gp5wnLS/Jnt+VvD
OWvzsbvsKhgSESR7e9Ip4axP2IJE3hAttCpZevjRW2twC1Ng4lY+TJLDH3lxSr/f
7mLtp+Qc/nJiW11ky/4C0kUq8dU7OcSuoEluuiTWqeex5tu5ZFrLBrObhJQVGp+7
Z6wXiK789ZrgS4XpXfyiYqd3OHFO8OZ4cwlhgaaZK36WwXKW9K7lvIf0IIyUIOKZ
khOBTFwUAVMjWORDF92jGLPBtk24usFeOD5+aE8C+u0TY0iXKwoSHAperjasbut3
BzUEi2pjpctJ3tabVN7Ki3S1T0UfPOBgVjJwH6vpzHmfPPJpaVZ+H6g+dGiSTgB3
JhEbU34QLa6D8zHpWJtWTRx816IMgwcl6rWr1urtA/g+r+sMAGJfUB+8j6IG+q0G
fFB43MKdJwuB7IXCJ1yoMQ8WhmPEBtlqBtXNP3WSE81g/JVPiTRNKJOTukghYrPc
177em0aybXnSeXw6AaypiYFwpZFJB/EDt/0poyLKXdElDmxlUvk5PAd2mH0i54P6
1v4v7dDjeoXRpactWguWHVJrE1vbUkyDiWAK821wNM+APdtUG9e6oZOQFmUeyne4
UErDAoW8v/ztdTsO3nTyD3PuWgyxd7XYQUEDamYCYpfNjSAm2K57eql6cmbRoeNm
TWcdyLy2co5MykWMf+CL5A3t3Fq0HN8QZaCi3PWHW+tYu4z5Li9JVp+tZH9YyAFp
mhvnbw2T2D/ukDfg+4ZslC7gw7W60JtFocFugmkUtgbvLqpn8Xr79SHfz0GJp922
qY2qw9XujLjeRmIlxPY4o8oUM4Y8epSnohE8Zt5W+dfCRl9zU9pUwGQRboPRcIN7
tyrHl/6fyGM/QTyo9j00Q8kGgNWJOZjG25+s+w1HUCEhaZQ8qexK5/P1PHrsyfTN
/ngAymY4IJjpRGCFtF+j7oV9qTV6i6v+RdaNBRu+CQJEAI7OvxK8Vrqp/wYn9eQd
n3ol1RSRHka1zoHJv17Jd2fGvHVBPkFxPb8TN5u/M18T3WeHP0wxy+LYYphA3lRc
G9Nvl6CEw3/JbJKAxP/Nv/OPrxw1sNEYruf2AYxg1dgEQF2/d+ETEMuBxFr51nmP
cpiu13KYUpu1ENEqi3YlHw+j8qBvm5jhDpTYJ5dQvYTYbKqCQLMd3K+bOug/ij6R
d07A5MPoCGysqVYj00FeLg3FiueGaRvLImIOblMipd0H2Ph5o+hLvMyugoAmwkaA
Q9f6Yplg1cuxXkVWzULhdAVgYgbrdaQgW9L1803GsP7vJm8/hdls1cgAztx1WFiQ
6OchAlUFopr0y7G7DM/nyEJUMn13gBCE/A42CrDvOteYuvLVmD5zDy/3ML7WovdS
VNq6cOmz3j7RnqpOYszAF9eVXeW5Hamp8Z1YBCC+619UHndHG8K8pfURWQu/FtxC
Sn58meN/Us33oR9TAeIqioYTpf25SCikeUqde6IfbN52bPjN7CuAiCxEBtUOc/he
Xkjj1vllTUwbBr37t1LE1LYzFcGG42DCPFhocJ0mQQQv/lsaRSKYmYmfFC3LCLPU
HKF5e29hcIMu4nwweBRftn8j4G1D2a9E7DZPAEt3+WEOmqGwPd/vNQsS5iW/mP0P
TExRIQxR8SFmcYyZW1B8MMNYMjuKpxXje8PW/UKFz47CWwMAzQ216FE3SPqdqDko
IB7492bT5XReWkMk8wrlikzuCZ1aNX9jLnbFkg4aafUbhMBJUbX4mRNvyYcbA46Z
0hFzVnHxKFjxH8JcaI9uadCLAvHty8PB/Ai+LDdjwl/+AaRCmL5Bm8jATHhSPnkI
eu/fq2RGNtNqFNH0/rNXS1oM4Cjb8JVrs9RJRRzozy41ehItKMK634YmhjDS5IOy
q3py1aTBha4IaiGWRCpm8I7RoqOv5jK+Eqs7lY4gxDndopyxlbt8bhuCgVHIYu6X
iO/7osuPhju1xz9M5Uz8kIPeRgFZ+6dDKPG2sFC32VIoXN3pxYayJHmSoQXfJJHh
UdNcZlxd33cx25vY4ZhzPwW9nDq/RjoI6QoZwlPcFjcejGrCfLYzqwRh1FLe77Rr
o0MvAHOIgcFKUXhNxuxgQCJUJ7RbUoF4qQxAJWgvKFXdMAhZDR4bPn1m4hhtJKB6
essFcBr8vgFf5xXbJ3aBxc1pnLkEs/m1Bt20LuNr3hpuXAOxZgYf27VZNQyiAyCF
DgWhpwEVEmPb/zdSR9SPZr9NNL7KkCExvjP153EWp8Bidb8a9df9JjfOcyiB4JU1
N8mJzpSJeGajicXDcvQiHRfya2HTdzFsWlakPWcd34jGgPmtC5o/132VpepeOQlN
+b3PvzN6ayQOwFA0pJdtH/f9r/Hd4nCvBSUB4W3EmcWzqClQ+HS8S2ljqKqYNSmy
CP7nY7RV4jO7xn290Lx0clqSzClOb/6RxHFnHrvVvTLi9kMfEJk38jw62conrwew
RKQVmwlsj2qxcxW/tAPLGC9hoqdPDA1zBvLQUx3oSYeh5U2xUvi5YhXacTdlpSUl
ZtCW9TeqT9RGt0Jse2GJcg+gZ2dmPHh6aaxLaPTSNxZ1ORCkXyEgn3xjIbfuqlsW
XF+jWglIxyjzDvnro3sBEQf1Rh1xuXAO9IrV8dEW1eqo6WJwTIqtwABFPbhT9Cv7
5EwKN8aGor2QRbPF2E0PsK/DkYhGMVf0uU4O6xA8c6RFjKFLpqB4P9vtyA9tgGQD
kn8CBfWiaZ+4eLSMw3xLwc8gJ5kYpUsMsYiy2S+8XD21BpfdQNbFeo/2JVu4UZ/V
mVQ6N1od0xuXFxDCcDUxyE6IpcOmKyOL/0rcngsqjXKtQVDsvPx0L4Ch2kvWj5GN
NJC6U7fbScEsXnolSAjP43zh9GCVvrY4pLL7IpjjcbiiqEowcSmCktm/3GZcN2fw
S5SHg+9aQ2B6RTcJ3FOB/U4ooh38LlcN/slLiAnwFyhci6qp2eTeL6m+5kh3DJ6b
tD20+pkKI/CDdAZ2wWdwiup1Vd+GIi8DlneJw9wPhPuF6L6EFbt24oDsucdFSeeF
en/lhX4pDA8UhKKRc/Lt02c861gBP70gOD/HjHpFwRyVqecicyJl6i5rSJGDsZOe
69GIfvWlZMv6gqQMuP+d+y85HslwQt3qmd5D+jXsZeOacL854u8VOot5OIzeB/Sh
gO+u48EbUwMw7jew1EsM7xLqvAEv6BPG+5ilznrxuuroPIh7IzZohhjl7sSkX9Td
WWLcWFOOBRhdGmjNCCPPhy+lGqGDMzIEVyAH5FQQCByFKZTRd1+KeHjTS+xmwsBQ
eAXREO/48iMEwLid8/m26+1wJdlGOuJGpAeXmnXOF/f/wP6roxTu+E1zjiuYKF2M
3ziMB8E/n3Aj5j8SGFkz8x/+nQfTAXXHoTF5v8bjscFkcOkoahLlb1Dglots8t3p
O0qnnEXGPUpe6gC/2FY0IXTWQHoXiaNjEP869wFyZznShzn7adkfAoNbxnqiEs0L
mzWzAXiIz7BRTdsZgrKpevgrqUWkFdkrchVpJdySlTojHaEVFLBkzFPAka4JCJia
xOxrgqmpcaDZFvU6p8Fbw0we4L+jQWGNoZp+uyMSuzuF0Q670T46BIDPAa9L8Su8
oaghgZ8A49+EBd3R4EbMOfrPdEgVMbQvGLIlgnxzX6sDi3nW/1gfO++QiwvQI117
qfS6iPjCSOn8nz1Nrjuzq6gcTP3yvI4JrJECWAqsSTX3hnMmR7ajyEtoVHeAWdfK
fMr+mzb6XL5cf5YZho6yFfC4AcX3+c5dkPePplSY1k63Zjha/f5tWC2TXLmy7UvX
sk7uOAT8R5yu0mDN5bK+XjwCkX583zUYsMb6k/pu9lb51lgkCQr9DlMG7+sGwdp9
MCge0Jr9CpMUHsO2Qz3i03oCEjI51kaQQmx8I77L9eRIfy8MNlDbx5JQRPkoP2S5
FwBc2eSakcr+IJAv8C/rLUrbF1PQgHvD9IynBeuH4ur/+fCGge/fZp32gUCeGNct
EGgmUyzYq+pUQ8fD/DPjUVtYCdbRN1rDpP0IKMNC8yilQiorwmGNHJXSxXnW/FbB
QrMK9GhlGbAO29kMp2i5XL3fVgfD4CvmYzZPwdIIDsdpjSCXvZWTZaRF06ipYi52
Y+iw5ih4uhButWnG5yhVlabr+oGdStvIG91T5AcJoell5zAfAmbK5aMG8b2vQWxn
7aIYLPrywNQBgMH4Ql6zkxdleAZUNYjgf/lzNsJHErM2RJXQy1BYVHTZIKzs0BmO
6POt9JBX3H0LzbZK1Zj9FptbvV0Zp+HuBeiSOuKvfBg8a9FJp1LxebaKYIgtjniC
qYwTPL5AJQo6DlmWDAdeLWOqXonQJPZvy/wiVvnOjB9x/KNwfCjD7QmXnvna780t
Ax4qvOeyexZ7OPOoGAqHFkR4QilyBb2SHEZUObcokWKxfenY6vRJtO1KGXtE+H8p
Wg/tAdn4SFUUi7nfF45VZIYc+xlOMW8/JR3nFJ3Yy7UU3DaTFTd1Aetu6cj1U7cw
xt9iFfmLA9CEej+70R2afMJ+1bo+mmNtNHM+mkIEa0MpHW4VQUIEI7NiO+EEIVMs
BIMqBVkBrw4XIR321lzFYWyRqhQX+oezGpP9Bjopzz5o+DysWPlRKSo4HgQyqKOz
8o8iCJ8l2bjEI46RFzhtnk4puqV/ZGfS8j3GRoCEzfE3Ds1k1yigtPIVFX3TJrES
s4Xjc7zNA83d3mFAS4hDg74zciBRM45mm0WxRZ7btq7B4ndyED3tZwVZIEA7AqAT
UtEGive9oxPP1TvdAFxrn5Gmk524VgIaTsrY2jhn9IzGV2CEE+2mZGEl9bFEEqt6
LpprFW+3b+4W2Hjp2vV923ictz1do3+TL3JeX0UNwE2IYGGlBTs7PONDH7svkdES
ztRSPEY8p1WbEMjZsas51TJ6jloYDE1etvpmIBUY32MMvrVpLUKtPhzGYPThYNmo
D9Qly1vs5GIvijFGsG6a6QzRT6GmaHZWUZs6j+MEhvz/NTGC6l10fWC2MOfrY3gp
GtSKQ/1g7La3HmyUBJbzmWthGolKH9ojXJgHZAt9bZ72GBhVyNvRRFsXgJ4QaUJC
vCvseawCuWCYOH2y59G7PIn7jpdYCU4jcgiSBOy7v7CbqNaum+0dPNkLxNW1wo/w
vdRu0nQzPGbat4ZfyBWRWfjOEPs2B127MaXI0fyr7xx40Ds1c21HqTw4NEzBsg+E
VvjLxBmFSGSli/3iy2m4JqJNTcyGpgrqeePPeO49ozzqcBHx6WOIf/ZFMIybAqm/
pQtwOIQe4R1kopy9tOR6eUGzv6NCejiVJELWM80I0e9HPVpgyubpu5Zbl7qnE0OB
0oJVnds/Unb8bg5lJL51gCxw+y/amzpNwPh5gBeH1IjmvRC2ykjUapBAS7GBZKrN
zlVUauFOGv0dBVBPwV4jRcg357qts7XAD2ML3qeYz0Je/nwEzsVz3tHOR3NypMts
Oe4tY0rhRDRKrZK3Y2zrL4y+70OAJcE7nE7pxTpbWnez9SuLLp5Hwg2Q6Q9Hrjn6
GpEXwAvZiKq7+c2npiXScGD80562oKVseyqA8X79XH08+czhxzERTZ3REne/mpzn
Y5jz3VDhk4FlZXfieFeUyr5QGCey72YsClQa/xbMPOMttchR9ypKIUEe3m5QJran
EWR+Ro/4SpNECqpfOWC3O5R42EVKwrslD5Zb6OxGcsAjKLbpAJy5CP4JHOlKN0dC
yV5UQLUhC/Tw/NVEXDwk/2nWQUIkpqJL050wKSLty8BzKZ1l+OCFig13goPy3hA6
C7h7H9InJhudC/Q7EkiG7KYZoWJTBtHCe/yK5MCo4w5qAG3tfV/OFlVbY4WnWiXM
/X7cdV83xaN9HSP5NUboYE+raRAwxKukTQ5Jhl0/iJz5jHN7KL9ixbzOQYh46MZ6
Ooglb4kkIjoc7A4EE/ck6eoHmU2DW7SnQmiSjlDzgKVG7BAp7Q7oDLGC0sWNoASd
j4GO/XbRDNFA5p+oWrKN9veFwO2o4cgL5RkEXzX+qviKN3XUD/ndKtZit8a7R3E4
X8k3tTwrdacGyn6kXOvNsNNxPN442xUrBpNUiJdw5wcBdvPeuymzm7US9GtJRQzO
XRDRirduQQ89RO7LFKnpcd6iXbw4EyFfR0HMcvdh5qRBQAatfNVi6XQufVRqArkL
RbP8+5f/hwYwyYEtzqo/ycHQRtIV2V0zHtoqvZE9M/ybsNg+IpuJ33MKnC2Rm3yu
ZpJsFHD8W2WSdqrI65DYfgCXrW59FV6AcPQx2npji2pNutAaWsl2RuOK3Z0X1/aQ
kE/Qh1sYgjWP3QZ3QmT4RSP/KcLfPUvOf0Qjyk38Dip1tYsUWx8MgzltDk0Ah30S
ZnlUNkowm2sUWYeNhgR5TGZB2AVe2mt6w5ov3EnY6MrhctpxHkLkf2G3h5TV1Sh4
OWwbS/gjhlW7KXtSSBxGtjTdx/UUpW5PiGL+H2JvX9hSWM+RVw7LtRAXWup6QdLI
5h5dW/k2jvRhA+GTUVkVPywST/LbBSLp4GLpqiOSY6TD5SwSqn0itzQeOCIT7eXL
M6NCStjBZ+0qH5Do2M6feWkoybNpkNBI3Ux3MihewImW35SHPCc570esLlaRc3Yi
hysE30Tevj8CRIQkd40vspHFa16p3ACnQVOCq3WG1PlIxLX0GOx6RgA8CDNX83/B
H4P9xKQbqaviVlY8EMw17UFp+OntmPWVsqrur3RWDQN9Ojjc8dEG9xyXWPqg/kJP
TjyipUPTj7QkHJ54pF1FQP+Ti6L61Nxz/cxA7nrWxL+UzyUWt96bEJ/JeF8v2F8Y
ipr2gTBh8Eu5OV8y689lEqMJQflHocJsmHxf0VHhUVDa7Xo6EDRdYJ6i6o8IY008
LBhYF0cW65mAEUOjKkLNUTk6leeC2KzYAhdW7sxu1szUDYOVEdQlM7JTsr1ieEkJ
EpZ+GT/bjZwC5zhAa205MH0k1Cbhjnghy2S/mLppovr8uFwtd/TxkCIGLTIdXWoB
PvUcwwe55nRp1KY0ZAiVHfej47XK54mpanOR/QK25LpVCVWpfbw0o2iU1XB8lEjE
QSYd/JqKv9Ou3402WzIhfe+BD2Ss+MOnBfALB7cgHj09ukpMyd3tesWxAIszAJjU
PiGG8mUu+cVwtKv3YR4Xqsqrj6NLd5YyvSUPsvQCeF6LjyZtInJaeoMSb/FIT7t7
ZJ557P9NH5OjVpXdN2JEHUA1o2oDrfmJmqfkVGGX9lWrw5Vc8fRdUvJv7l1w7Idr
FFsGEhaFOz55bfoUfdaZWyDQHvRA+/aJ9tDOW4bTVOe8ceqt7vn/LoS0/cO/Aqm2
X5nzbbDHQnoL0QO5YHqNjJevwOID742uHxXTjCkBq0Gh9E2U3GXH5xPHVr7DA6tn
umLno+FlreUCnIM4P3LhC9/80oMNpbv0NP24BFPTpAMil3Mn4OXZS9RypM+Sz8Es
A3r9LvNJxM5Pv7w5owG3EfQ/NoXu8D8nKgbmO2Uc8mMiXAVmi2FBNM8p6R2jls8x
Sd9jdXe6BF6iGn9fAjwdomPRi+TtbMO6VTY6R3c09lSvYnaQiIh4Q0+vte3SeTPA
IJKkWDNmVp+2X+yATLCdJqSwxeZMISqV85kFU7C/xE6Ki0BTcUR5bpVN3LsSmuaX
qDoWiPxBDY+TKGpfa3Af3ilI7JsODqLCC/JJDwVqr2FWnTC8Mn/0xtzTyrsiyiqY
Rx5ei8MagFLbW2VxTA3Hm7b6bM5lhZFLEoHD1gHoH86zNNCYemyRMAgeUGSiCci+
4OUkn1Sf4jw/mmaVY/iWCZrLJWLcNgS3wjBKpz937WLewvb1x96GV1SLwT9+wlTl
jAPU20G+x6VcZzmEX7JiAr0tVdhgjmmK7+yVlfIQiZ8FGU+4VIVK5NPz+ShxC/oU
mgdq4ACbOHzmFpmt0Uw19X2o1eYxZjTr23Wx1rm8vxF2QUWsftZyr6iJzDOVdT3M
F4B4PVVlwQJYD+dZxDMNUQgPRVxN9h3tF84revKf2d/Lq4FKHCgyAeWD1cr8Fv8/
cfsebyBoa253x4sf3qivksWU8jIjmHbO4X3HUkT7IfsfNCFdShVr/5RkdwUFYvFg
b08l514ZSdnEsbaDTeI0Q3YboYF5kLzYZnNBupSopAGfOEQsjbItjZBKt51g+naD
f5+zR34DY2AwcKPj7qSL7v7qX108QbiWaz8jGsjBZmSf3XUHKJTEyQwVeqfNwpvz
NhYhvmKiNwofbQVJP9m+FIeS5MD/wzaYt5dgsadGvoowYlYgIc1VCBREitLjJm+K
4Om1xIczD/NynJASh9tahosVHmqyBalujZ9wh8WzcB2Momh9pagi/zkoI7dp1vl7
La/nAuw3ZjxEWo217b5A8MNnH80h6m7jrezLz8s4KcYzn3WoiAHRkajIwcvR3Gu1
Ah10yEDhgR/swiDQWN+eq6rYbjS+1vwELgA+U5BAbFV7LYqQc1D0T0vxdtgczZeI
C+nbdmhoEkzWQBKWKpzQ2Xo7boSm34iwKamsShWjUoChu8CI/dQR9kvYZ+GniEQG
BHvkPx59jXe0K6b9muWFiaa2eS7f8CAKnWn1kba2WCm5sTHuGGjKd/3UxbQUYeBK
1HDvsooswC5ncZYzi6eprNEmKKJUkETMWPA9cl3mPAtjDygoAAwzKzqI8FcQw8ny
oCfn0pSNCsG3O75RW61GlWJ7cgrTaNeC3UokpBR4kS7z73H9oEVefeAcZ70Xng8i
09VgJaOF/Gc9Fw/n61cZd7iWDzu9hhxAIR8KgZWOgikrAK/ViJXMWAPgf185jnEW
89qm+ez2XjDR0wtWM58vmH0YcMvxC/GZwVSU3RoVQft2X0FTrt9KYwCM4g2Ili/j
24K48JoKsviqr2I/F1jJVX/lofd6sb0jt5VBUM0RvHFdFOAj42LNm6MANadoiXBE
J5TdV51jttcEYMasX6QjA3QpZ5mAF+MP+RA68uwG+2ymKWHSRvPiWfMh/68oyE8S
m92VH5JTNyBQVKPhxNjkPJzspbJn8y0LwKxkXJriapa0XHrNdI2OAY5+LRomskkj
Z2sCqzfu2qcDWVtC/ergLGKOlHRz3dUyL4KUW9cxg+u26ESqRYaLnpPkQ2MY1KDg
7MKKcN49NCGRxNyhSW0IGvHIjVciE4mxLVNBFgfjOyJLCfb/u6y2Bu9vRjdJbbQh
VXYqNOSuunppa9PYWYrAq3TdS1dSPusWowyGQO422ax+yBaYMicDZqLNufEuzeSY
I3aWP/ke+LDi503M2cWkW+pKPENdtoOujdcwQMp2CrgwPU5w0WxJnY/WPd1hkR7Z
dIpZpU9XlR7iqZlE5Xi8IzBnXk3HKQiaq68vodVLxR0DdAtON5ZovZ6a3HECBOnj
t5IU76wi+s/Ej+KjSJbeDpwK5cOK1uhKVzAovDg9W5Q1ANNFy7B4SUhQDZFTQxLg
VC4F+awgQKktgkbt2hGmUN176mi/Rc40wjUt5YSK4/quyHtthUsJHLoFUysNJQV+
dz7TaiUbUnG0kRQDP1gu8A2EWVM5mDoYglN7tx5yLsDcSdnLWZa9TBU7Gi9vGd2N
EisWslfcruvm8yLXk08XQ7suXF9iE+khB5gcKLF4PCDY7V56Nrc37tuTsrJu3V2a
NbMxC3RdtRufDnB8PlxxmOFAtCnvxwvIbasDhIYEjBW5V6ie3l0fOshRC44GQBcJ
0RDoi3isqCranpID00UtsvLEZUQuebfk/h39KiAdmO9heqdzXUItp7xz9bJsKw9W
K5+2i0l+H1t7Far5OEIFYvn6pFdl3IdKmxx5hqjFLV9K30Xe2Rh/OEuSLG7YTAR7
mUHyaY5DTNR4dFXlO8VO9t/Tlw+NfyIKPpjPVxU2b//pz3ZN8cXE9vjQ+YHbJv/1
WfXkyYVkbVm5/iQdPyOTD96SIxtYd2JVTG7gF7VV20WM16nKL4u6lDQXHvJRQRNW
MRsMw8ArrYvzfQ7B8vzZYFlg8Ik3gWVFlNDY/Iu1CLT9T1l/sp7zi58kqG4ZgkNR
XPpSg+qqLI2zdvZ8VZKt+pRPyuybEvLgaP2xEApJno/LdQatevJDw3SJ4CJZQ/vd
0h0iPd9UL/aPLQXZk/ArgfsaIArhvu9p2a8dPFJWuY+jwMWt2h59DBHtcDA0C1wP
zT2unFNWWBqc7okAaO9nGqHjIgCCqU5YUwKNsQI1E5wCq1Onf+1uEMS9oyWEmHWJ
QhREGCSFMuMty2/qNWB7+iqzRKOxy5b4AtL3Xrwxta3t7IMGImECFBj4eujnc07t
xbj6U1kcRUh0D0s1q4F6i19718nw4jLy69F5uAhgrEwpuha3rI5DPD6fb5OPDpvm
HIZDKlAXcLhUqxK/tJ9oDlH0TgPuXoWVZfh/v7NDEtcNlSymq+l/Ni43DE7BdDLx
1T7jmecNJ8Bvo3YuYDEqup8dVeO3Jjv3UWmFTaSIEeBpEeOKryHk1z/FIl40fNsC
91A7knVVHWuQB4AvG2VSQ5w36URjin1t/4v7j0Zdj/+c107M24zCjXpyJ7GTLGm1
huztyOw7M7UWfH8ocyedrwaFlOQS+6q2ps0doQLA1Vc5LqwpgIr9zNEWjEmde3xE
Obcr7s2P7n6aGXy1la4qS/JEiQui1xspMKF0EM9utmHuPJEGr4ua1mECPX+HucD3
4qumIrjr8ayutRr3/qfrsmXRQo8oATHJuqDXb0GkJI2NTUZw2PEVgHUVDlIiKy0C
XOa2sRXO5ot8aWD03aYrBRfzBp+uDb+FMtyoS9ni05w9/0lwG1M0YN/Y1OWIwwH0
KsDVTNBCucQmRma1ZEE1r6siyW02qqukwODGjtBEgCgOWSBAkSi22IeoYMHexN+0
tg6YD1mOWVekTEuPbejZuNUjADyzYxaav1w+Ls7AbGP+9tlVxT/P9N/pHhNOGWr8
IHd3TdtzjeEglYLYDEgsS9e22WKka9/O1wQ+VZC6dQo0S/+9S2qgh6iP5L9Z7opk
LZbFRUie/yGGYV7fzX92KS3lNZLnSAi/xJkXGhLFYn+Pp8BLpLWHuhTtD+WS+ZxB
9G9E1A1qBG2tyd+wTItMRxu/EB55dC0SZsP+3yRFasjzo9TlD8T7ndlNwjkdUeLD
IgcTArbPYmONjZVMKI1dskSenAqZLzqllGxMnxrlmsgVjvc/N9Opovad60PN821Q
6M84z3o248mmVTllj2m3zUCtCREnoH57STE+gFP8cBgpcyabifiPwzogqqmf5Q4k
VAlQfPdhDvTpCfD/gAlgNbDoCwCKnoqG0nCog80eckFkYkzRPiaeyl7TEsdsQZn8
za8vu2xWf/SPxZHtuljjLPSDjxJ7Jdwoda3RHrNUzCZFwlF0jocAJUcwB2Zt22f9
+o88ZCOprfGMjOFqCb82A4vviSH/YMJXn9g2tScW2+KJO9/Nc0YPxoqIoPmhzGMC
8K+tvNUzUOdRlRxL/Kjw7hXVsZ65F57D5pefuK6hl6SZ+kPkCKzNfQz50FM/6o5+
a7GVnfYkjRC7NzbsYAEAh3HWquBqc3xaXN8eq9cdGZDjgMl/ByMgmPfGcNK4P8kq
r78Ri+5BLDrpF45KNR+kjuk8zs4/MpThRufPdkOx9u4ys8VkB1z64GBD+v89pulE
zrJxo7d9AKfC043jG9AVmflDYPSjN61eUuWz7WbNW/0mphl1/r9nf8QrId5IUxAD
Lm05qR6ZAGrWxm5iNR1dsvKFwlVRotD/F8KlgKXJj8HQRgCemPOljyqicLQnTr9p
p9SE8C4k9SiZyJUVLI4zjtWwPFXkgGdrNtF7g4Xr0Ui2iS+VqC8/z/6yYcl+b3rm
FI/IhBeSEACyYXBxk/4yL6pOyi0XdQGg7v7BKescCPS1juN2KXQczwXBZSopH0wC
TUrprOFAJ74AeIPGyD+Y4e23EK/4+o/15INr8ycH+Ci+doiuQY4ibf1i5dMo+EBP
/1zSilNnrZcRwmVBZJ1VhrTmt7feJorsISjKwOLcA/DwQEy35BPyCu7k0Xd+Penr
Fj17mrox58pf2VYl8IWSymK8HI5Wob5RxA4XyBYdOfNlhfwc54UDiT3wcxpIx4Ps
wCEGcaMYShpYMsd3FYgd8zQsNRwuxJzAPs8bqGtyaxHp56YxS/sevWpzq5x3/9xI
mRBOCROGO9ooQO/f5gRdbhChMSz0GrmEzWhuitelGTT5T/I/8Gni9EqtaEg+14tm
D+z2s9FTmU3Prha1TjuZ8q4LufWmb2MxJZeg7fonkDu8lTAF7jhsbz4d+vZdPlDp
GHRi23QfE888+Yq8EEcix//TmvsNtXaE4a+zm9tGmNe+sFfET0fr8+kG0hD7BshA
Spsakjdl5KUNSxpAX8U2eGy5R14v5cDU5YFdPYaEvs1gX9g+L7xX+GML7g1U4W5a
3WO/1snsD4vKpjrdHwIytgaufbZHeRmZJ5RCyPK4oUC2XtpL3u6XPYJT6rBCdZkR
Xr7jrUO+xr165Hbd3cXA3QpZb5FsFUV5xIrGCrHI0QPLbsbaLA3GI51bJn/UhyR0
1ldnXNfU4sUe5EePrPkNY5bklKcx//oP/mmRz1i7bfEeh0B2sjJ2UZXmrQhtnNft
3+BiYa5f7OflaDLDae8iwdy2/8au5q35MFQyGJxp4yyIogJFc8v5uQ2402MjQV9o
+ozcLP5JcGCepdfohkbWgkFYJccvTBsVFg9Mnq8h88rjqMDM4f7PQSN8jeTvF3jn
7FMYXzm0KNJ+BUoF5/d0vLvyisWYM7+Is1bFon4ZV4878t+sB4uQDtiEcblzRkuj
sUPr8/qF3rKxf0yrVT+nxu3EbIIu/NhWMgh6QqGKY9yQOPhgUl56XVzc1fS1/vwC
Zk9FEkj5M436kQ4i+eH7aLYfmNx4QJotuOMN02OLrfVzjaM5YtmWiIn9qNvecg4V
4BVfzvxpnNNd9QI8katiWnoUy8P1HQwR6aeYQNVXmrf7sz7aVAqaVP00QVQ1zD9j
DfGcO+2CKmuURwyNSHGFifHKHGDied+N85ttc6sjMVKAJESClVM7UxhEkeBg1rHQ
Slp8HoIP450Q8nTD21/d9klZTVkBdsQHP89nLHTp/DdglbJHSVSVFf+JY9rEZ1fD
8xqqzkmL6QJVLkR4T4E+7CWcfkDgDq/YCgA+V9EYyUvxRhrCH7QLEkDGuGwxNels
JeszJ+Bjw8GeJ5YeAKyE31BfYdS5sFQnrH+AwknRZ+EGZ3OOyBcZgnbtNp6v7duP
AL2h14a5zyxjW9axjMIXpBkINXHYNO07LMYfmNpsFvqRXGVM+zNJS+xDUM2O9S+d
pBtMmI61ApqpP3KWXZpE3//XXUQotOd8Ti3lXcNQuK8rhzg+j9h16SonFtXA2WOS
SrNOcSD93KfnpXipU4GCDB3HIMefAkADBq/lvyOtVhP7n2v7gSjGkFKFqgeVPwm9
t0VpQonUq6uWlCWtRMypDqIirO8juh3Xe3Oh0+mcX72cu2BlDr0v7pbYlN3ya170
P2W7uwQ8kAOpUQ4reBntdO2DZ/Ueg37R4VZjyR3G0CJtR0J1Xqeq56xlZ0V3lx44
USd0d4AAcyurdfa5FBEWp1Zj3ehMq+pmJlzQK2TunJ1Xntn/5xrUQbp8MAOBTtCI
+nn282PzEZGnTHTz7TWgUdgTC7YyX+zpcbcKkbo++a9W9osgIfyC1ecrwgpnN293
+m+0iiZQu6KdScLLGflgxsnEtDdcdym4s9lFsmOPY3NyzHsIh6rX3/3MUu4mJTXI
LxSPGWzYtrEHfcbdVwTSa1H/Utu5YK+0ezPlTACpZIG9WPlfGll38QUqN6KKQwDc
scAlvlADv+SJCo7JVXJLis/3aEKTYt5vteMIXisCUCihMgtwkZAQA+88loECpVRZ
UwavpDH01i2mNzOfwWMvUkXGl0iIqI7EDDLQ0RgCxe7894M6xwkP3N950dEVSJ+s
i/YXFpIS2GNxPm5KULsJCD2c3B9rhkD4nxlMXB160ruyGxOHAZKzmbkGS+I66bsS
K40p8RkuvWVZz/iA2lgs0tt4xJZbMqUdpavcadrWXrFkq6UUz23RN32xG/NnFl1u
U+6QK9sSYaY+jjUibBqjrJ0GbzuQND+ZhM20hPjzZbwSk4LnRwknLSSQkrVeSzcI
kSWDWEfcVauBApUfWmayYb3YxfHBdyApr4ZDssCXVndW6MOoGurDs5XR0rntr6pE
yNalkSS/BXj8mUhR4o/nOXm0Yz08xeAf6FaCi74hceb81bsPE6ZDDt/TXY51Xyvt
2jnb1U9vXLDEHi8s54yuhMbAaIRIzXMFq3gQx5O6oU1llizSSmnW5fM/yYkDKomd
xY4CwTv/1In7ZMNNUGdze6LW1g3/0PH9fpFB6QfDwJNh+YNyqNRHPzN8t5sYNSl8
R5MfCcOYjGifpyhw50TCwigFJUJQ+OPoaf3wj2fjGfHH18wDCb0iyFuK1IHg5WZl
RFf5v7SOlvJi83TyK+hxOqS8mM5iaR6W6FQ1b/oFVHIXBdppJQtS2QOXrRj/z0WL
MU8GgsVq3ishBshUyZR1xruDHVb5QbWDrIF/rWL/gi/hA8ZX0eIqFZZJ7M1D3M/v
x0DpcSLq65oycXFRxw/a9B2Mx6Iy/LeeAX7c8Ubi0JzmeQoabS9jfQmI641AGNjt
Z6G/eYspO2k+Ai+Cgw5lo7vVpkE4Dmy0vtuJBdGmXZbDT2UQJt0CvLeP327hJ4W5
gAcMw70IutuyCOHsGbo8SPtS7M1z1OBpjVLNnnQ8fSeUbUWcsuq0XzfR8LNoUPZd
u7Mw3oV6KDGkcj4R59fAqQ7jyWLN1si5p/iEUUtPI33fAMaiMEiTO83o6atNC4Gc
icmaj3LNOq9mjUGlWo85GMKN4blY1KYW9X1H7zJWvb3frSQ5xaEajdAerINHOwpW
MEltX9bw/E5kWuX++651GUww9L8MUNAb5LNtOfcm3e/EO+9l8Z4F3d+fkv7rKOzz
K/mVQWydLw6iNseLiiXd/dUvvJsPEnpBqpS8tbQHtBb/Qo3ws0KjA6KH4yNn1OJE
kOjoZzy6EEqOCWPcLqjB16vZqpoKBrD3W1uqggwFFmckVgDGdECOQQEmgLpDsqIE
fbsgiZkeFLoD9YOdGVfGyCJZmws1gVE9uGxT0EvVwO0QjmmfBIMpPh4ZCIJTRL6l
BIzm7K14ItBCJx3IXxB7QVeQ0KViBalrKMCpCiF+MhE0sbsZYjPcK0A+/XjivHQ3
Ro0pAJVQ3I7frlhvp+bMlEYhiel46Dkn7pkAo/UqEky9qve5tNsixWOuULmC/DNN
ObSY//wcjGsdktVKPKpE8y2+csh8GBiDEfh5dnT+C3KaYw4mcdyvjA7qu+UVJKUa
gPerOR/RlPcPDnZDD3ThfSgxV8Yb+FUiC94y/TzvWBnlLYRoaYckq4sXX4ZMZeFO
st5F6hoE2Ya7L7Jo9iZNpeHwg5GZBvamUVqMKj/A9ms4Qc5HQrh9Um891ok0Crps
XJW48I2wSzk0ez40DWNhuiIrUm1q74EBRqg0cFmmV7qIJcWjJM6tBHwUKH+v8lv9
MH5UP2QWIYfWtsIKx/lcn67OoGOf29wxfYevAJeH46Wgl1nxQDDAxPmTqPxHyOsr
RvTD/izXHLqhigR4zSAyzLrUHI8+MJNvNC2e6FGGzzFh3MSSsg2aVrtR9JAnP1xp
L7aJ/2zvUyGwmgVV5OnlvYy01R4ue+mNaICCpCG9VKDTFFcDl8Hj48LkgWXD3e0x
rjExXqx0et6DxJq7nRjk4B2RQjdexPe4IxNo04he8Egl2wA5tcC6w4J24KQUN2+D
vd5YevCmhp6MpfS7Euu/sjMMbicAvrT08HMJVw7iSATUylw9mpq5PRsY4M1vCgnp
oxRT/DEH/eygumdLERhFJsV0vQifScbn5RkjtmptvTFMaOoGFUGVPLbb56T/PD3l
IMECSz/AnZ0W5c6clNv6NtJO2CXxt8LvAqvBnkftL6Vb7HtFCNuLMDrVDtMXgXje
rg2n2JTKsCCFZvoF1hhfHmLVjW5PX4vVot3tBYqr4rqhdw/9f/7MS1AggPokeXff
BWhkFbVdjUOcNdKKSoy7MZEQDdEv1EpxSZGxKAQotyTSzZz8xcFh8v0NI1HykWls
u4Wrkyy10I1crq6wlaMDNNSUFG6c4+smYSvXKDfXJaeNF0HZCkgWfzAsNivPkSgj
Od6/CI6rLTYKBPjwYxRQdQPtMb7X93CJVcbJZRlFZ89qbrmiTJyESj29ljzKs4/x
nYsVJkROKibrLpK0fC/YjjMGvGR3TQo3UJDA9rxoMdxvWLjQWGpjUCrg4dB5EkW8
XtfbfLtybs0iA1zaZDXtb8zcVseguuaykuyZKyYr1fSoLk3voVB5eK6IS9DWYomJ
y857i5/pu0EXfAEY2TpsED7vl6DcC9XjEP+qA3EjkJ+i0pF9nfRTUzF720iuhjfD
rsLK5cqVVyshDLbZ8VHmvS4FGV2mSlFscwuUTOf+1JFt8Q9BhHQIgk9dCyJYGgR3
8fYWSyinJL7s6xcaX4rNGixPS4q7Zd9qy7wzZXCjQpq7G0AWIxfHMLXPWzW6y5Dr
7ZMVT4J8EO5PCpdTFB6360Nomu6j8uzVIqUDK9m4lervK6OGV/jQhyKnfST7ZZ8I
RV6IqTWMhfs9+hiAQDA/63aXDm1E158j5eB4eRg4xtb93db7TgpC4fYJLfG/lSly
PO+8eGCiVT6Uq0t+3Dx21Rhrb9C4oswrp0drnkriDgDY2uOFQLl8z6o61ak9vohA
6sLnVOAiB8fCdggUimqlmgXM3tZpilR5QwQ9Mpfw3btH219B9/6rmROHrIIlKqU7
OJpLug7meDn+aVjWbSMru2tc6cAaXqHdg36O8SlvAADkMN9iynIV7BAxDMrY4Arh
gS1f4qtwAH8Mpd/RTJEDgwx6Fm9XyCY/NFFjVT8/fGaSewmqEWAUR9HefXXBrf/D
+Nw4huxx8sQ3c4KcCPdL25Es+NT4us1BBNINJOrHJTdNvF5pBKs3CDns0zh3Fu2g
kNqW5jqWvOMxXvfjcNr5xyD0dysEyJ9K0j7UZa3bvNnnXcdpZuv0vcdbVzCtQ942
d5JNgvtxydqEW/InhDERFbqH25gLeTn0Fv2zj6Y0Ws0+PG4VFKQbOTBUH+lKUmjK
8tQVH6xmLb4JDrAf6O3vH7reL6S7fPlks6Pk4PVwWmr/FuX7zuE3LvMvpYltv1kt
Gz0l7ej1bmzRXpineFTGZP27I8179DuxUp+BFuGAZmCE1O69NGWbj00ndmDfpRkP
SiRrYnhpXvw2pu40Bg51ZdATceeL1XXRRh16X6H0rtd4XrFtq0eE+PzSUA2E9Mo3
TDsPop5hn813EgKq1PG+Kwy0b73GO91amfdTOfsBxXRaHJOquQBMVAskSP/fqI3p
Ri1VM/L2tgsQFL73/ibJdWjuL0DSeLdTQ0i5X9YArUx0IhZGavi00rjS8hhCq38D
rVtcleRtXd1l3sQ03zhxSL2h52XY0FxnACm9DAPP+BFQsty/DWdTLoBEgI3GuHDy
J7wauNt6ttaM9TzWWPIdJW85yDOT+21E7liXkxXOoH0xxL6gD9k+MMQhiasRHQis
IzHi8pTH+U90Vrspq9LCquRxD5/bj1EBQApp7eOlmfX3NsbgudrtEAlIMBrP0nvf
uA3Hdq/JmK6qMmWXUW/hwEiYIa3f6ry5EaJwV8NMAQMhYzZItpfLixxmdsERvdvA
HyKDvQMdkFzLVy/50J89Shrgce1CIGvpYYTip7KzXTZC+9duCjTHfDn21VCxRiw2
E93B/oypn6VdEMWEMzXbl8hAudU4DxZXj1kpwj6Zi2D5HUTY3emLgOKKzqWaN9wy
dAcTmimsV+CWsS7NstYLETOql470clfFzYiJJTAtG2i5RF3GvYY0gM/yzRBj1L3L
ZbhnNBp5PPZ3KqRMyMyS1E1PnjZbsxgo0WyPSXfz9wZcLy3W/8eJQuc9/dUUDVWM
IkS8EYFGjM1YkLE9tvg70TCysdp6zYknxBcHBfz3Unw1xXC313UAHEwpcThyFZEx
ErAlGCT6klumaNdoEUt3aH7QEoiLoUD2X5DuqQ0gzWgDoKC3TIsVgHyKaWsDd+Qz
1rCWYGERmiDfYR82Bk/gfYbZm+/MtgrILtb5+hF8ekRHNpUQKlBmfAxVLSipQvE2
xL9GqAVIg5k0vkC5FqA/fQT0z01kW7dktD7+za6Om9tKCqxAauc1debrrD3zAp+j
tn2Oz3KzOUSOE8sgshKAF369E6exB7j59YfkpOQlWu4jeZxk1at43i6oOl3pk38/
w9XT2GifvWZeTLi5HDaYPIRpwXQxyipok81EdJxMWZNYzKVuLQYSZXaHKzEVuaot
u8w7LFwLQYytlN/g7SzAQHZKKMrKGQmLv0kJc7Hif8F0WCBUkqaerrS6oIXs6NFa
PjLIrGy4nHFpuH0glCe9vPZ91Jx5wY55qQNYQEKoSmjB1k6gGebPrHRWUJ5VStF0
F0tgF5qRyGM0w4+5WaFw2UGxCecZVo0xByvWxSFJZefAAuFE907pTl1Alrl15T9J
R3iKrO+AAN/22PW8zpOeJGIJDXQQDXOODsuVO0k7oKrBrrhJKneAtQL7JM5evf91
+jUMrKJH3ugNzpa7Y+IvUuYZmyB2OkGJ8I+t8CpAzgsnh9GjuwqMe5Qn7nk/z0Fg
AudJAki5m47f3trkd5QfoULL1SUk1Wyti+kxsx0iThv0fGyTh3MRK9D7DmTEgcGe
HaZv6sJVWj0Qf3ox4vPzhnkFzEs+IGmCLrpdyZfA547OZNA/yZmP3g1XMyMc/enE
DZrs7y587MHjK9E9CWdlbYT37Xz5xct2hE26EL9siSxmcjwjvfTEIW4dehT6fgsH
PwRRUtXUniSR0OSiZ/5sSoUO3f5nAkt8Rcd5tlHPLkKPJ9IETUMkqggZ+Bvk3loR
HRYB8yMFwbtR6qrKh6AvMWW+kGnVDVUNuFwA+WM76fTY+cic2yLuxL/VMncBVFoV
W+ZdDWbaDErHtcb6uRrBF41qd1OBUzXSP1OEvxcGVzB2mmYpKjRF7BCYWYsM/16U
rAmTwJ14KJvjLsfVJkVbBcC1bdhuo4zNBI5UxHAvDqp2iVHaeaeFnA2uFn9ASeIW
x0SO1/3Wzs2ZapLUTLDfoNLr8G9iXodNSOB8PqgUdM2ppGys5uE/1yfG+1b6o6qC
+QuZyigyTyQZbrD20EgwCkFTAbFaE5bJ5AKeplEJ23VfJiexpetiq79EFBr/fCu7
TjHTixJBnIzQ93tiz19VOZgjujKXsU9IkOGZcwqoL78IRTg4503ASKwlJhBWoW3X
cjVedNor6cs893UH7+eKZN28gtQ9Q6ZVgq+U1nfYs3NPw+Kt0tsnVkwf1ogQcLVy
xTKMffIDK/0sadLx8HQ6okWCmZPLKeQt5ZqptfkwMTn4h7xVjYGVRaqlu+3LFVCp
o5GnDT2x3TMIUMXcRRDolzHV59zjx6W6QD5NZ1etvQ1aWtExEf9PjdbxsglnfrHG
YUFTMdibeyW7uIh6/PoumK3nAxB1TcXGfqinODjKDmN+2KOTUp+15rW7W6HTrmnO
OLqgCp6UwAN63Wqa+Pm69WATImLVLmcsOyu7owHlteOoeOvSREXZZisVvcA9VGEW
4Ssq9Nn3WsRBGUyF3+vTAiHGqx3xtwN1QF9t9Mqb+GM3EM6+A0qk5yVnRcUCMwJ4
wcUsuxLdN9Fd7LTo/wAFzZMWiys6UT03y8seH/L2U4PZfOS2kmQ5pEoMFGn6CO2q
o/E3H5wdzrj4j+d6w6/kscvR1M04Thuu4GlQsT2Hkw/Y1db7Gs51bIe7lG0ECxTq
vOdiDGhsxuA7H+PCietVUh/3q/YHrAN2ld+T4QWvc2dAI4ps+xMJbUVW+JiRmrkG
GcsTDjwFHb9yQAIKkg6eSuFdvZu4Fzbt+5mE3t3DMtZM2CsIhBGPRQ/GtwsNPWRW
aJ0HM5ZCQZxwtGsh+OA17mlb/k5TeQfq7T1hKSubhTpXiZwx+uW5JEtbOwSoyrGI
nkeb6x7l1Bdjo6ty7s+PrMFw6KupDmjUhtpPbf4fuhYTN0IpdTRGsiD8g/KS6DrW
crMy8bOi1+viyPgjrwOGwqk6JX3NJ7OMVNoTu9mqHRzBqEE1K8o3YXoZ6GLL8WE4
IRVR84xvk6RNbS5jpsYz2cLiIm2sRfXmHW9ktLMDPoUjtlgMdiNULjzUZNEuMR9R
oqjxHoaLy4XOsX64TlnFfMfmnHGCI7Huf/hhadkcILmwTg+EymEwg9feSH1k2SMq
bSE+k+gE9rv4NIOeJLBdAr7ODLmhBlXONLXYB32xy5TXZNvJ1mxMMJzh9qFFOxxp
3/ytWw6mevkLl3faUIHOc9vE3UjXX3HLT12ppnxoSU9us183WSEC+JaolEP/XBLh
XrK5Yr8k2FcxgjLGL1LxZB8bcfQe5OZC7GsM87vT8ANgvTeyMGP76z3VJXY1hibJ
PDWv1yyhY5ZT+/DH7NSW0sq3ejq1YPpARsaQYTjTdh3A1p52V/uewiF3PTaqEDmx
LfgQ9JNTSfC2yGxD/kjhZh1cdBvkFG5rx1nQVWqf0zXWNMd2weu6Vf+PehRbV98i
vd/q1wqJa76bxBjPCjXRbdGjvoYgSrCGdShT1u2JkmKbFXxdN4ThOIff/mrWG+yG
gYSZCqpCGelfq2uRHjWZuSNVrjMbLk5uhawjRw5QvmXammrvahtNJ95dpM0ASrHn
zk89LhmzNdP+vFoJVzFZpntF4ORt+dncCfaXCIDZ7UHKZg62Zw2hfJyPVsnWAhIO
kA/Q/d5WSSZV5Xz7mWtD7FJSPZ0DSEXTXVoe6OvC6WJMVGmxj2D8PO66LJpA/prX
FcM30keTW6YNZikJarEWEJtYcGkpgzbkrZICfBPzr2xtsllAT5yrdbQy6/xdpuYT
N5PljkrpYWRADM8MOzwzWqencV5JIO/fu34CCUSm4aTftSAOJb7DVXQN61P5Au7o
6Ra25gSs1c83VfyWE+ESK5p7cZB7z3J3QWCMzVQLNLJUGqGxlI5YuaUn7iyNQJmk
lSCqvJfwBNB1tVxBAkMdfla1QMo45aMb79v4rgeL22ozJTf2xtp+5Hd35tEb1lM7
u4hl9uBCBTSp/U7DKj5dPRh469QSnDT5uIPYcsNPZbk2uhE71B9CPb0jrLgVKIqo
cSrP7M/bokzvIn5wT5nY2/a2S1Ht2w/Yoc2LYbIwzHySdPJAdmB0Fwht3qeYmZYw
w3FlIw+On44D6xOPOxTdcPJunYLGMf1akrDsVhCl16oEhd3iBzQsy1sQd4rA6rGb
/y4foqwVZ99rlgULUd+Fa+EEdMz0hISSAj5fWGAHj6B7D5FJFIqYvR6v54V03+1R
bh5isoRWPbpdoF4yVk59nwOc8Y04dkBwK+Z7LCJTsWdKv6BlAIS/vnuGrSIJx4LW
Sbo+1l3VqaZttKGv1otHkAsRSUO+hp5eRgJ9DogfAD55vOam/IzBnW2ixVen60EL
Flcf5AcdliZDoyb0YFtVIEykR9aLkrk9uKIFpvUaKpCPGbMzTnYxrPhzWMveq0Lz
/ZBrvRbLcEIPFygbLCR5nRmwJ2v90c3tcO7Osz6KdLai1zFNcga0onGOYpRcrV6x
Q2kOxWnd913uqA4Pj8KkKKcJHCS45MGGcgJHf6QJ6TkqwkJSgL1RbC3tvwrBUJL6
Aavsmk0avxwlxc8uPjG8FaFy39UCF/mi6eRYHS/YUBO85f2Wf/0rz3iAveQvCqeP
ZSZ+kxCSuKEOosJ+5y0FM60n1i0PlDP1/KGo88IS5U3jmMrsS1yL6HFIaOroJFr7
543C4ylfucz1/79yn5IiT9CrDS29s0dxFM1pq6f7GXs52qimiZB3LkpdvIsfLDeW
uMFqkRZ6Q8WCz1kMiIYl0e8L8eZEhHgWjBHZh9dPGo0tZIem3xqUh/DnP7LttX9y
3YCUx4eImDkG7kRe13K9rR/GZvFXJbmZZOHfEzHespyduPQ7D/ie1J0kwQw4wj56
AEFfaHhanmFlvRksNsh0PTM1u9NdfssNMlFVP+NWBf7UcwdHPmV2Ww1l/GGBlFpP
gIVaXKE8OfD1Ionhtu2QegXCL26miE7dsLJRU3IT+l1FMIkrsp04g8vm8pY5jgLX
8uzNf13rQjKkJFUFzgYWxjwfS4hbJUQ0/28dxZMf9dsQrnv5ErAXWQuRRkwfxxqw
PIUAzFaKJeSlvfAcv3CfMWhPRFDj62p5gyE2Nm04P+woASdB/lIWpb4l3BOU8xpv
SQIq+H5+k5VxMsMGNWOJl9Gq8U1hz2krzvMPlqGWKRtwUiSzKZ3nQW+A+rdv3/Kb
Hq6aQ+rC3vXNMOPyt5p5RfPPcxgORzNEAJxR9yLnlKXpJkYooq9shtDm3LF8ALJh
eynKImmcLGwNehlIoyE2RbCu3XVT2IDaYsfrzI09cYD5hqiBCtxKpSadxYbfyhD2
uGSjGUXf6g+S4+2ejny5tqx0GvcszT5ZHXWM7bHfqaJQ3bpDm0EJqETFAUoVHsga
NH5KoopPLFkOisqpNxnGba62igzk0n8WC4eBC+6TwsszsDbg+BzKRDD7WP3yK5vG
Pc9NmcMrZDPnYX7YbbYJpHHOEcuPFCTr+V48FGiezVDRX4GnJi5M+wFmF5Lp+sbA
NrTg8wjqG6M2z15ImHldz56xJ7J8Av58W1bD808X7Mqf9qLlcKN1gbT/eEv28ZSR
AlG2SfrCEgmztwjbgoDYeLzLkeCd3aW+lGcfHN7C1B8frX5hUyEcawC5RMzTijMm
d7fB86pRtVYoQT643fcY2p0ULKjbe+sm9kBUeyf2idU6Zms36tyo/cn/NO6A5jDA
OIqld4k1GdoGv972yqTsmCv0npWZDCt3mE2iv+OZsuef6dcY2jkFKUaI3RowBoTT
m6246qjI3+QueIM016rRRYn1UvNXT1r5UEiG2Y2vd9GMWo6Bs35ooySRua56k1S0
BBwKWcmqnSS4GxWQJEPjPyIbWgVwLWb6qDyVvi99b8DWIpUOn8Z4/ZxIopO7EkmS
Zd86MATU3sTi4TSJpZ9Bdes78NGlbdYde2mzOXe1G0ajqqrELTsBfZyAw5AxJ/FR
9K0q9Hy9VdLxs0sLVHUpNJWY3gRN60rnLmw4YNnmjhL4yi2j8k8Ymz53qAUxvtT+
j/8QIFYZMiaZKg3ItAKdE3F7JXL81mDojRX361bhYZKRD3dcoEpClWwooFfKzeJC
1qjmclUGudg0TPlJi65wt6t7gfeUjJDWmXyD66I52po74UdhD8//Bo+IuSdVwwHV
1z6B/pO/gwelS1uuChyTa9PQS3t1K4BOy63TKpBRQgUeD1r6ZirFYz9UCXxPrxFE
Q1vgVGNBixdYglrt6Av5QqkfLRz0+P8kzgfGDtCr0N3WFf6ZmGLPSgHteR9uKmnV
DZfaxsEoJolWooMB29nbK4SkRWQUylhh/gSW366kJy7hMX4opBn5rd9PxtJPL8Uz
C1D/Rq8t9B0cVjqdjQFLf/YYI1O3+Yu9o57mmWSWozyROYDXqIcDsa9/wgS94rig
zRXI31Qk+fXr32Hn7/wsFiu/7AEd4UBES0g51oNuu3AdUmul3tfF8tuRdqArZ26m
qTi85UgWPdzHyRwLqPibAtRPJwcg+au///mm2iK8QvEqdROH3YPbZseR2HTHJt5J
KQRUAR1FZKjcTBCF1RQ9trLd8QNVfZDu2p9FLlrh0zd3Qg+AXPA9atcux9+A0904
qdkXDxGqXSAAvLukObiB49S0rTFvoGOb+4H3abxYM5hBazanCyQr95kuYc5Ca9yg
wPYX2owRqTjPbFx1ddH9+XCnp9Y4s99QiLG5DZmcZbWJ9MOb0E7AVihLxErLuTYx
MqE+lz3gC+gYEPbINzHKQx1OC1kn8Y1/Qzq9GL/XS/J5taatcAxkJWroAq4sKHaY
HWl6ttkGdUKC65wlp/MnFPzyXG+PZfdrJK+4XGp4gLprPYQQ/3NkPq4GF6hvZrCB
BYH627q/eWgGYZgue/oQhlr8pe5Ckhh/fLWVFL3nhRL8XdwJ1xLmQbv+DK7PrR2d
bOVhJKTKHn0ZVYmPPR2rmu5YiMGygcOpdTJLlpBwLa3NcdmZ609usVL5tAHDQrdV
wcZvvphoWHpfKTW0Zdf+6rx7txNvD2pgljgcGit8MtThfWrTzmqMW460TJ4Sh0e1
1F+MXq3DgCoS+e8jbLYolFK0T7Ds2kiuFD+22o5lQUbk4g5tfsV3eilgI4juwAVg
DG5CskGORo77b2HBbNOr/wnJhiCVNsKmVB8K1yw4/BxupSNtuaQisK5fYZGaERZF
UdZpv/InAPVvo3RwyKhWqqG3c3ya90e4hIPWc7+Aigis9PjQIKiNbvkv1nbagm0D
xbfcOiAdKqqjb3gPFHyzEroBdGhjQmQrRP2Z6vm/Zc1T3SBuHDID74AaWwM3/zX0
q8HG8GTNOQPVYKQrfn7ltgRh2kCKeRbE1WN4siptpSb+GlvKLASeUB06FwvbAJCy
7iBK05JJXPoupdCIiJqKapGCXP1cDdvQ2l1568TYfBIHgCg03dZ0MzB7J5EcmM+s
+g6/1tWXVpouiKcfHHC+SFk0DRZtEi8dQuUdMswoilvyA8zGvPwDgZhd0913st4M
gRPav6chZTT8BmUzaHRldQcaWVAhEQerY/zXY5Z8beeadmoyWU1gbahxgGP0OK40
zzpBxXOTlwDydOMOEJlLlaNs1sz+AQUY5nnulkC+AtG81hys63rpdQ/MaZ1WaDnI
PLSAGAPiL7Y5053u6rDcl7It6Ouh4ua7aBFZ6QKt7U7bTkMXeegibqk7vb7wuNo0
n4DH70rXpTOGC3m9Xtv6VTsv33vG50CXzz7jjVMTl0dzgZoWCiUJNbO2ejR1kxYT
9zs4gA0fJsro2F98o3WEfECvLxQxl4lAFD9oeSd5+pstlRs9oNeUInFnVeIYIj5I
9GLR82AJgevXfJGvsPKMdlas4V++jTM6gY4r6C3qd6PXfOJQjLyj1UzFGDycIAHw
pb9n/RGvH/HxJAWEeuYGylZmn0Lje9r0Oz1Cofx6HO5ySrx2cT0TJj66bnJmfnHh
9ph1fpmomSDFeBlvwzkjkB7XHsJ1vYbcdosLpCosayQ4/3JZ3QtowxUF74likU+r
2LxFvlFi8OFMAU1DVh75kj1Fclw56Nf1vma1lrpHy8rTFE2ICBlvOszWY4U9wrY2
ubjkZSWFblBLarFm8py8Y4tjH7lhYFHstO4Z0ZLp4M/HHIoHvHAvYAASsfWhYsuM
wKsW/9aFQ6x0gv/w3T8HfxT4VsxZPHhg2QdnurNp32gs2TQ6x8MHKjsDLiCql218
sm1lNYqlt8Fe6Go9YnhU+RCS5chvcIYZ8l2AowgNpSD+ef3w/nqgG5C9F3oUaEL2
GJbMBoj0I0SH0Wo3qk6ky+EGdwfHYcm/2ekXrU+YRJjiKOuG4BhGNcDghvDJ96i0
YaMQA9EqEov5IlpDKYRIgOfdDIjMn4zk663osfpHJ6ovYJBT+F7GH6YhAy4YNmjo
FUY7tvl2Jt0P97E0UEeNQVqyv8xafw2iFXsMJ8sSaa+tp/0751sEVT15LWjNRUVa
IqcpCbtv6nXCJPJtmPtnC7SAvfYXwRsWGIf5JJpVz9JM+bXyL9RYiOCygEnbMyFu
MpGmifFkIUi61Rrg0fAdoU3XAOCYBumyo2h3x1FaZzTxb9rcYlBRDUqjU6+beGur
UaN6+uVH2++XqqVGnLH7O7hsfBh7fyWyA79Qs3hn4Wg7/uaQrSYhfjiTNMWZazF1
3w0vXgJzWX0I0wHKSvAUp5WE3dASXkww61Qhi0kU5BjD+Nuqz31QUbcwnfHoha16
7pbmlAxDrB06R4fTzSqHnDcFac1FY72IYgZ+NTIGggpnF14vu7v+0PvAgVP9Vh+7
x+HdHVV+9P1nhFpSHJSImFnJszg43eKRWzTqh/necV/Vd9m4XJLXvtGRmYi7BMJg
iw7ZIrJzqYb22gwc/DfvLXThisD1MVLmnR062JttRRXwTzUcuOSYgAD3WIqKrybS
ogqP72yVl5CVMuqXVL3MBI1wBnp1jK3M3kPlVYb6shhbQ1be54+6vY3ifb60zVUY
2qCKuAUQicfXKgtsJZXUbPBxfoi3E7X9TP94GY4PADDBVJ3PLyYn6UJ0EXlOtC3T
bNxUnRqMr6rjHiY1rHxQQ+nr6UHeCIxBhgEaLh6zy+rSq+NqOp1qWrHBsYy2m5rK
Nd3o37nKHhKfvqKP8Ydiyva86p1HLuJcWiG+qi3i5YWsPMWbi2H9gQYiBNqbUKZf
2k7S8VFahKnrfjuJU0NBslZO9C/ZMdSHkJFZ78rC5HlAl3HPHKeEuMAZt0+dvJA/
RXdKoddTxboeDeVnfs+ldSMcPK9CNLm5KGPHkbOPp/0cYu0xm3eHBwe7AnshUMmt
tgXbdcoaUtDdNTBzTdjJ7dkgyONlrWNORcWhbTsoh33MdZ8g3gYs1+TPPxWSy3iS
SBT0LjX5SdycNPJ6pNlTvOLjS2VnbNqVgQgoD4byy1kP37km9pfY2cEpbY7rnshz
2Sw6gAPrQyJChV/UBiAxz8p0NhaqrxB/XOvxa8l1nYlVEsbC1c9j5MxBybFmd9hl
rfd+BEFYFKBSbicVgzwH1nSQEg6ea7M1l4Au8HGDI37daMa8Gi/Z851EYuWPsg0u
uMzARwEnIvV0OpbSsmHuP8wNag1oz2JZyTM/gPjgQZcdeSFFI2BjDS1FXbYIYZ8C
S250jsvU1atWi0ZvNhcHI9VTEKS+bOdm7cwmeyTiFiMMR5axE2f/HX+A6+MBYYDo
UYJxn2t6Zk9uQ67lFuS0pYNFFBtMuK3TqnU8GW06LtsFTTBx/y1RxjvflkZOBsoT
peaUZ71szXqfHtn9O34lxdCqQN+36wR9qtq3WFurzar9MsWZcAtTCOYEoegJBPN4
srhUZTm+7r5LGOlEBd7pMEgWPaJn+adgeaz56zuz6Uxo3U8FHefg69pFh0Tv2nTL
1gJWx/R7g/H98ZvdsvGKg1cP8XxJHDpAmFBfTYTN8HzlTNjXUEpCQHG3kT9BrKfy
JKP31YMXn++DK5i4F+XKaIC2+MkInq2cTKZwEzdESUYZfJNu8yk0UfOdOKQ9cG9S
cx+bOJqFBS9Oq+2dcnnDdMvxlZItiYEhWgBDMtl5/DHIlmKL1DFx4Bn0IFN7AEaN
wexgPpJ98FErYRNa2valgkGkoudF06RXzqYBCd3gnwX1dJpuQ+OmsiUNSlvYkQXi
YKa2KiboJ3CWzwgcUdxLaumVaIDU3U9InznyugkDIivwE/etcjiVYWxgXtQGkb9h
lP+JuwUqUNDAFV5k2skYIL/v+Z9jPQbWNc006Gsl5bPszF4O/ntkxsUr0jCaZhKa
90W5F5CQjCnfV8ZAzhB/HdXxUSy36VOLPF7qcAOQB4DpqOzP6bsiUCmRGTmRh6/I
MzPKvAsd+ND8cwCrbvfTQHPLO5CW/4zP5v2G7u09UZk4gygcwHSL01ExrW9B95Zc
HQu/Hi9F0QftBTiCvxQ1P2G3FoM+dqpogphlqaNbuE3/7W4qZ7GEDtW4u6np2k+w
zRXHFJqKYatYehO8Z15KbEs3qKID7zBPJusg/Hn76KUmJ2zmqecU2USln+XHbBsM
4ckbacKSd3R9FvQGBu3I6FNhYkvt1UGc32dusP1PUfkdiDtQ7oMVCJ0X++Y1kgSH
1toIx1/r2nGvKJfK+REmvT1/VDYCdZTffu7WPE8NjgNKOOZTBQCB+YvisEEBwlW2
Q66x5IRVreDN6cSwYpmnfxhl1ej9PPUHiE4FGCkfSXkMNUEDLbknYp0myGl9cKd9
FVKgKECT/t+VCAFul2KkECcVGRo4PpYm9dd3ad2e+1CLUd8se60+IiHJuJt6FluZ
0oEtP+5wOiB4UnGvzkZc4gyOr+0pK/PkWKs7IEXgHZ9PAVJQqeS5nl55QUJG2HaO
5xe4kc2dAEPwuEhPbQifJ138o4TasrmopB3bAykhmamsm5jnCx6sfs2NwaEFnRAN
i9P2VNFrfro/Q+O3eYGkB2WP5sntYSbR0HIZmlHfSbUkNssdRcgEob8gqaZdza4c
g4Z94ykdYBkcR9RF3xMCnz3MMGYwV9UqgEqj9QpqPbM05Rr6X5DxjjUvKfEYkb3h
FtjrQskh5TZvXtIYiG3AnGs6NsbHSE5zOLN3Ekw1bivZ4Kat6Gxue4RMhdsccuxP
fBjZ8evkOiuFeAxgpxIj6Le9GDonrtp3FBqvS7PwNMCUEadm53PZt/9pX9V+TeWc
Udxdnuhoav8zc4gxuLFBrVENZ3/il3cSsoGPvSYbJ0NQDCXE4/v5Tw7BMdVEytyh
2l0BynQITthtl/3zJSbb0MDDeqxDXdFqX9bkMWtmLdRKj3qvdJIKcpyG0QtZoZIa
fvQ6CJEYX1nONx3vZHmQKC//RVYYQHHkvEuIs7tTgoebMK6f6Iitqnme9cD/zg/S
5ZBcK/pjTwsCC30WDEKExGh1yuGKt8U5RbxqviBshPeIRmPoJlk6uthw6GUb4tDO
hH+GYcoHairSPaisVCyFLkWKBFqo55lbneGrTQZA8KwOYiql5SYwaMJoSo8Jss9J
DTv3WRnL0sMstw3/WPsG++Lf1eRCVXBSqOIfKO1KFLEt04LeG2ScrdOMDKDu4TQ3
BDQaEf1aQjH+o18LcChhKlHbrASfidbtljm8TkI0lOaDg0W70vOJ0gAgIL3Wiyz9
RDOmKRsdE8ltBmLEVgS5NUgzoLJesuqNF5jcckmRunf9h+J3My83fZsJyqDuwAbV
P5NxzGsTf5Sr+31W99jj5KcqBFUBotw8OIJYBN3WqFZkx+UOafqJGdtF2ZHzNBIr
b4JuwFMpgUbkS2ASPkx+RpPHanNh6vcTCJRHISDScPe2oYuxi/azmRlBrfwyL7y4
LYw8hwnvN+d69e+p+ogCbochW7CMiTWE3tMy/qmyf9z6lgo7Qm0LdrsTGE0UYMcK
/WYQmD81xF9Yy4ShNwyIfVRAlJRvBTbF3ZRHbVKVyVd2Jc+087ICPWt/qQwSKEBC
2MxBV9v8SwbD+az8YTVbnV3WghUouMm43PL24rm0HlwJBBOYSdoB3i+aVNPIFMj9
ZZwnhWF5zT5m2sQQIlBC85rrW6KfV3jWU8e4JwAKKjIozAD8mD7/Jz1B8PQQV5FG
MWZ+bSrfYZ/JG5kPHlTVhht6qQrFSEqNPN76P4HUA71PGzb/aHOmH3al9iv/bMKD
q50DGqa/fz9s6fHKyVw3iNGsXp1F2+uCZJqQ94ZRLGE4lE7ZFVXED3yAKMgv4zX8
7rwVYs2mU2o6DT4wmgCwl/3PGpwx6Rs4G0QJRxI7vSPrNGPVZ/9F7HZLM5YkcT1c
N0hFgX9DW7eTC9c1z6uvEqgKI7v/udIw4x18bU1Xiq7qCz2VlWNAFMmq+LptDvnV
PxXWrzHWnDLqSFsB9k1x72mgP91bI/9KIq/WYZCYAtftelx42BISGtVWCsFzJjSq
qIGr531YN6oWIN2ainrQDeqIL6EaQhmqdK8soABeAsSg2+HsGWQoufQoBt6OcJm4
a38J9u3NHODDIZayuJrI42kTqTqF2v5hCtMMIhp66f3fGqgvCJzqx5V3mXcAkLAF
ET4NDzsRTYNVprrBNLCk1ov3EuButwImBNTURTEPhEqYwVmeO9Ofuo/7GYxN0VPe
lLFN/t4oPas3piUpe3ziowrbYVyVDfXjqKwNnrjfjqRm4OlMCUFEQzjJFLC7d4Ja
Lv+lFC7QMxpzNYWh6LDD5asvnGlFMOrmFh5Xvp9DtXrOK7eXMcLN2nGqDWNeQbkD
kzTnD9v3roZK+eDDlroUFT23F6jAqTRR1UymUh2oSnZIB1fFv4aP8sDLW7kozqTs
umqx4Vz8Lxjw81B0YM704GVa1zuplOF0DePVQ4PhUntBvPpO6DyAUvWiTj4g9zdD
AhWqBiSrzEKYtNDMqyQGs5+4WPSuNCxL9kMxrGbRZiIoGarT9d3igWMfHfA7Muyw
WrBswzXbMzZbPwgJpenH1+3QvR508D0pxkFEmkij+Y6MWbznRgiFVuS6oR9P+yoW
owhflYNS4YLQgnohoDnHZOAy1YSiCDLnzLbw1nsV+Mvq9jAusnAVEsuHld3eN430
xKcc1M3xJ6WOLIBP6/pL6Ls4xISZkv++gaGUxo93JEyaXC98kNos/JrPlgDgJYaG
8hZlWtlpj6K5ctEzh5M0sgpz/aIJJwnuqEePE1Pa0ZmV9MPtcSJhyE2o6CdXut9Y
9gtWGKCa6zYpWWyEGBb+r+EL+yrjB9+jX1FG8CTCvACvntVxIpjgAtN7o+gzB38r
ogQ/Ceaj0pvPPDSBigG9x1jCzEg3O835I4qP8kFjRR9B9VG+dSH3F3RuN/VcqRw5
ZsQJe26OqgNu/tCAgrJQ88/EnfzfgwnPIkTvaCXwa+B8UJXEF/Ouk92SryYC/FA8
g1HiOGZU2DOlpaFik6Ki7kGRJehHOfKHNTI2ZjAJUVvAHx7ejqSiDxNtnn72GQia
ksYI+mBuNNz5IJ4QrfRjkSJmtEgPj2xYJLWHX9aJnRRUiXgn+mLh2PgIVdonzsh4
aHj3WJnOCk6gC/3jcmBHQfaPtexkiba9+KT45GGK8evS5FOaT3bM8riT7SojpFSR
Kmg7naIFkd2AenIryo3+iB2fdhl1kvL30ZX2NpKEIYAO6Ov/7WwRPE3cXFQWx8oB
5uBpknAXsdsqLnekYMxT0ZkVEcFj+aNCuCIAn4ZlOjtmnCBMDLl87nrUp2cfF0eh
SQi7uIy0WmR3CRsd2+kYibJZYdnz1kaGrnLLwwBaiHQpEvhHFEBQ3ZXJAF3csXPn
wwnOYkkNk/fvxoY+bv+b5LLz8c0srHOr6PC/gHZyFT8kj+qG0QyQDktHyR/4aRIj
pIayEMOvIcxlMhToUKYdo4YNfWn3p3KQtkg2bBtbpp2suW2jU4qcBVbwRDjDCpHW
uuiYR5HLTg9oSkXc8ikLQUFUOYrhm0OJJY2meICXXhkD73+3qV1WOikqz+d24mPz
HTF69ynUE2c8lSAlBbjoQhNn6mu2sBPzVaaZcksYs1QxBurReuu3WcBgSLAiX6R6
onbtVrqImggOVTjyNiTP8RBkX13aQ7IQEtVL+h8rJC1BfBfdP4yaDLuqvr/HhWd4
dLT8fmpmG2srHGwnuMm8a+TeQRPzPLyAwV6xIxKBqXfpKjdS2Jh8Ja+zb/T9ZXjn
kxep6iLMMRazI+nX2/3UvVexkSWnERY+d+igl/07++ysEG7qwabAIRWvceV5FNKT
EAGg6MaodkmjyvoNW6u3wOdKNmp2hb3IjiBfgEP7ToIUqQg5BOw0IbIZTCAjkVCL
eJ3eP45g2kWR+EO7f6NHqxeqQrN2V6IAwNtr4B0JjwgJYIweJ6b7+ssFpQmoEVdi
mde/X0zl+C3dIYmLEpRggwKsAVq90OeH/ff6h5qTtPFFAS8+joiYDxLe2YGIb9kv
QodWvItPBD8EHPQ3wB1kz58KwltolsjVP85YdXeNL16B5IyRT6NnCvR7mHRV9pbM
m8EuvZ/OMivPGJsXL68K1z/ThclG/r3wsSgtDSwccrSFYHzaa7col7lZ0RWI3Hlv
jrLdG2c49Irk/OGKVe8Q7bpGZSoq2BIc1u0lP8HQuf0L0s4lyaIQSHDrn2ryKR5Y
/0+WbsMo3oaPZ/3fqEpMRent4//hrMdMjGTz6PTAiCRBiUrkk15z6ak/tSSj1pvp
HieX5MImsq8YCHFeaDb70wesQYLf506JlviBQOG6MZwPBV7G4GCSqFO0DxLHN3V/
i6RRh7Nx+QP7QEd5QKdI8pQT/hD4NF3/tUqr9LCP70n6ZgfigC69eLmGMdsdjve9
dPJ5hZErtTRt/4nTMRO+w4W8IePUnDPPLU2JtiKK5pDV2FM5HCN0OQJ2SYyEGMWF
RXm3yon4dTRVmvVhVSj0xoK711Rb9o4Bw6BwA6JusEt2e7tu7FRG/bWAG5F2U0on
Xf2lpSJWza20cr+3UF6dJxXn0Yy5KA19l1jDtqOQm/xiiFnAFeLVpQUSYK9vIv3q
685wiZ+iAgtgjS1Qk5IfpECuMW6wZvAy3zGUH6YVj2IeqRZib4sLwSiC1TKTk4uf
80sU9kTYKmqepDSyN3OfPVjLdV75Bc9B4BKpPMpGSQi/9mSl3RgrNwtlWbzRKlS9
FefBZCLqIYs+rfHQczubdYoekClklLrpme4C/TJjSIXAad1HYWQ2xj8ts+P4aRLD
9UTLeb04z7+SNo0PSzcRhXmuHmYZ37iYo+8zYF6iDu/hJepd8AEGMtmZQo7dSkwy
gTzqmGQwkeR/xu+bkuPopEOiYFGkDSi7xXaj98wK8kCWAZ20FpKA986cnLQyt6JY
aVJ0ZjCCaZuVkX0DU+OUr1knaWwvMgXzcgseX5Xnv+wmRKP03kfqwlytKwnhmSMs
Rw3B+9/27xBfwEqaFFG9imwSGcwuJ+JR4fdxttYXdaFtvqbK4BiXtD/cD0pgn8tw
4s+qpwgVW8qsLaEnSA7Zg99zo1Ala3c6RH6O4WTJvvQYolRjChTb8ul79J7Zc/vE
jHCgumHtwCXJMjVYm+mqNRTW0fZdFW9WTegkT/n3RZY6v7bHL40ZCZetPIqPGkJX
7ykWP/hnrCmxeusz/zXA8bKrsjMDa8uclGd4qH+CqNmYEzv4nAsApZ+ZbnD6JOvy
uvaCB565ocuuL+hz9YUNyfaWKQtqzlNcqxvcDUwvGRDQPMxGPr1OMetpUOONX7aJ
IgICtHupMN3UGrrTFfo36sviVdwr4rafSzZDzltWyf7wyRoOBrvMElrIieUoAV1K
jHvj+rbLmR8ga+/SUEwPpPUvpDLaPtMDTsBPhplNnY7Wo7FA3yhhvJyA34DE1jAY
qTFzeR+2UWhc8tMBduGhRvzR+HOx6yvo89/h+jMGGT3+6dihCbvhvRbHApVYCA4y
FebnaD+U2OkN3YCR8BI8RFUGvNo9pCcgNCbOhq71R+YMyd5BRtWriLkmeWE9A2O9
tkaKwg4xUoOj2RuPM0Li34FLrUYb96sxihHOhYpC/Iu3wPl4UeqsMCsIO7trn/Xi
bl2Ma9Kkxw8R1m32FCghZbL46V4QspcEfVC6KJUKO4Pu9t8Urg/GylquHesOGfkm
BdEBmNwxHgis8/RC5qa7Nt+A35xmg3hW85SmKLImW35r9DSmFBYtVSKgSo2gB1VV
0H8yceeF3eRSKepQVIfhDhERjdpK7ycn1wgmXS+rSQjHer3M6Pb6/THhkpZ/5V1B
WIVjaqZ5xBfLS49g9Kw+NS3VrTB5Ry8EFM4p55NLLYn2kxIkYZzh/bFgxH8jVyDO
orASoiQrfUHjAvUbupR5lg1LZ6cbkmKia1tqvVOgooO0C3VOu9RklFNwckuPy5Xl
4fqx0LL/G9EWmddYKJfYO2H+7kg4EIIhq0+TmadlYtWMaf83KRzlOohTMmFLXk2r
uA6e2x7JV8RkK360LD7B494RFPytf4BuTlr8q4Kf+zmY/Xae5NePVQr0uTb1jXcB
Nrbs9OmHwdEwkTxptIHlMKt4nbjwSxNVrdfYoN5YFmPBi9Q1sIzeAkn0JgPPubJ/
vTpuFuxQH0aNJmrVAb3FXZCoUvOrwC4dmFzMRrH0c1ORaz+jdtSAlslK1/ToxhZE
yLLRM2+KUiyVBw6/5TzMOJy80G0P77v1ELB21ycoNiDZFJ42XM3OrOWnJk9izLFu
c3jduJyb8a6snTCVtwsZZUdn4iNubTrF3NOaCm8w7gMXZMwKNlgMHlHDITtoJb+A
IznhVOPPD7heR8gVLqqn3O9ak7UL/UPQcdLH3W8sxx7/er2bnVLxo2UvfvKqR9tS
lqbCzbJzZtBCtt69wts03kJ8eE1cCuB8ZIDdYuxvcQJ44DpK7epyBV8/2x4hxaDp
C+683H2I8nbvNfXt64K3lawNbmZu6jBkwaHdn9S6fMiQkTlU+dxTAlmNYdVVAM7e
v1iOMaonk2ZtxKaOWq1K5oZSFFbrScZ5k2Du2zDf1yVhrV1vS5ADGbZayYupysiT
W/v+lBvFiOtM57TfaUA1YzKfa6lzLcMcd8118hqjJkswVkwmaMjCl1js3hu3YLXr
ZNew8zJvCtbQMTMcJI9BvdzgBid6ROJSVf6doLV2ZJQ9IiaYWdwjBDaw2+bi5hxm
f0RV/5VZzrpzn0XLLw6OoCzgoikEJvIYREgXS0RNHIcEEW/GCUEa4At3K/8qQ+Xs
ftchqTBV9SD9xgQHa//9Ib30I9aojk8VFp+D2B7XqrfPFCz3U8i7Ol5nmD1JZ5+n
jIVugNhioAEG06lfCkJcOwss4TCiAIyiqs0o8PZGjhBdPIBMOmY/hbpmSUhCGVl7
i81cm82s/1uQNvy60CygdaDZzE9Jf/ynhBQhfhi+sTuUjgqHEkpBln1rp6JXnFF8
xUdyZZJSjSaH4vICUURL5LAsPZvY/60jJn7THUdgEBh8zgDMBCa0X+At34kMkmqt
6b+slJ0R+DKtu0RT9fa3Z5C3NSzMx/lXZq+s7cfNDmnTGhi3jvMPLB1PtikKjVOA
tmsZMq8h5oon5pE0oN9ICVZrLanLPVgu/S6aczFkhmj3AX8jAbBQ110lnKfMNRWD
cqW4SrnDuUSIUVjkidpb3LBewEIVHPccUd+1VPVruX6YM5vi7hNfGmZb7T+aee32
wQA9Aae/2rHU81eFCCwn7HJOWuXwulxNnyk5Txm0kSZ2cNSVpJEWezC7oU1sHMj3
SnqAQfVFN4tuMO5TJZ47yxrsdLXUj86oiZf1GvpzFrPAurwdH5Bt8L+PAbpRc+4S
5b0K/3gliYpSKSoL5G5QdDq60Qi9YNysybEigGtnxQVumA+ByBwTGTF1jAQHgNbk
h1KREN/eT4euIi5dfxY1Ig7O4AoIB+JuoNWj2yigikiVQ00TmgwOuGgvbwYslLYK
o97elotBUFgL5GykdcqddvRV+/F1pUWYnjyxt15vU3dN1ef8pNsbYqi25fp8rajA
km4ZYdIctZsZp29KlCnqHLOzPdWltiCeRU0FZguEa39hP7mEmlm1qcuPXu4ZGNm2
DdcjenE3pSJ2ISsfaaKcyXe3zp576869gXtOC7vYrW1XldAwCaLDETd9ZRjOJfpn
3xFgH2kanBShgIoveHu+gdEh7utcU/GYwuwE3z0uEFW3MzmPW3H6niuv56TqYUOz
GgQoD1AGF5onSH/tZ3b2782D3xVAERHS5Ok8MoCcfPriciTk/yVdIbrhJIQCU8BP
MGjAzulm+qoZy3HRnpzjBJ36OQbEO9lCTbPN09vDScNAAmzfWge6q0zy6J3RyzbJ
Jl7Nb67KoF+Xh2RS1Fg05HYCB1B3oJphxieOyLhAIznoPzquBpiRJUV6D+a9t0I2
mt8It5fFtwg7h7aJhe46aySl4JgeWzlULSQ1RIKevV5GOdmYXj6c8qb7tD858i6a
+ITT9Tsi3DHCZsPOkV/mzFRBfZ4QYmwYS9PHdu6/+xUCs+3bEDIQECuPxMmH9JcJ
FsCyZSlbgL/2NlPrDL5REqefNvNaML7GIgpHWIZiFlmXXcHxGMLsPbtXDBuZYeW9
S9LaSzPDpNaZe9a9+7F8F04thGu8ViTSwnjiReVlLecownCko7I/bouamD/30D7u
m2UaUyrHYo/LV3s2Sm7SRM07Xc5TLMC5M+A41G86geqwJOMCK1GRQNoXWkJOSHe+
4cc348pcxfMmxTzTT/SpyqLuJEaG4IVNr5D/fd1OAL/Zceuyl+NMqAed0aw8ehrR
bwTJh3aossEtjmWakAJnooTHk/VnSJSqWvEzdfb+S7/6dAWj9dmor3PjznAJiC5t
uFt76X3u6MC7FYsquqZGp8Z6mUW2uMcH97IGSo6I53QcT47Nt9du9snQEANdWtlR
oIQoyQP/TwUNgtnQr+L9NM67QfZp0d7/jnJvAIxmYTktdQSsLJwKrl53lD//bgwO
gJdEnr446lZA/4OKDvKtfRPxOHIe8/UOxUCroLoHROf8pkggDTOQGgzMW32/0bpM
+8c55TghRgnK7N98H+FVjqpj0WLk1/GfMgRruX3D/7g8/cLFu1SZ8SDUGIVvkN4t
mi86dzd+sg7RjQ6rV5inSRpU/UkxdrS0CAfEEDz4jNoSGzvk9v1bHlXghVfPddPb
7ZP80/NGLtz5yUz4+bCeQbLgOtkWTzoVY0RgHAJQNl21zdwKzJxlaQY/5gwrrbUk
yECgOoHG+p3m4kcHX1/d1Yk1Ugi0gEd+BaUFNH7nEmq/rytPCwxIt7kgenEqSyCU
kAo+sAbFiAVCrYmpUt1jP3vW/Joy46DIOoxXJTV7KB+V+bdirZvhQqxqV7CdlZKO
0OLKjqacEMIOOuxzhWTKhM8wt2w9poEeIi1tXMX2KEu+5aUmRAYFaSqx1DiAbG9t
p//TqXFLeFsINznSMWlZYx2K9zDXWQf5wKL9sAqWrSJXcODe2RXPcel6Wb4gAVbL
+RBopQkywp4cB2BuY0nP9It19CSHUoX7eEmqEff7s8onUNDQAfDJU8sZuwb3k9QO
mAuZCDoXs6mnsOmYdCptQBHqSOYuKiGHnqI2nB1XGQGNZ2PcAoVdEWDR50IO5Qje
wN2fWNW+TmJbrlspDZqOelfcaC78Ez/Y5V0XDJcij+GgjSmZvDoOHFOR2oM/e8VJ
U0O+1oFh0DvGsX0qRBXZTAnc7TmhPE5XscD8Pa8NsRy66fGehVCQeugRs/3O9Fd1
lHVwyoZ4d0o13VvmFKEbPj6zcfsDamco+rBlivL398EHfMesufEfMzKDdcErbtNW
WIQJXyI7PdkR/fYPVDKlE26ztKgRKC/fBfq6UQ4/5v8eu6XvhcTyQA4Z4XSR6Zhb
2z5XuhpRl3RzWIXOx+U15vRH6/sp5fSp0ssBGbQ8NALBo+upJaEZvFHkyV8VFtZ4
ULquBxpJvgBSUSBmSN3jVzyQO3tHFJ9HLPRtjoSwcGbwWdtZmLlWf8UM8OtOSef6
rb1hGN+C/855usaoV2q+NwuAdPK8RksGzJeclEvKyxvevvvMGXvP4njJt73b8o69
jP6DupFS1BwTXoqAZebxZGa6BCz3wvu/XF6g4K/SUy04W8zPTYmc3fLV8NcsIdLo
y8vN3HGXuYHLwmDEbpezO+4fjHkyUhGfGG282BBPYZI7QNDvTFNHnAEId7MswQE2
d85HdRui36rHcEZm2czMJLVFBEaPHd4+5H9QA+Ti1UwSJBXwAItGTpHRUV8WGyyz
/q9DC1r7TF7qi4An+032dO+FKpLR/KwX8a0CBNELZhsWBIY0wnO40FJQ6LuVz8ni
2MTtHtLqmrWyXPMBOk7SKM4+Nz/oRPlNtmpzY4lskEJy3RCj2ugrFrEH4B8H0e3y
mbwJuyV2amy9DJDrtbZf2n8cLOFHWCXayUg4ND4gv+CIHT9Shgm8QBwHMajyVMd0
BbRUjSs4kKWer3vnop9bm2ztwUMvvy6pI/RGZpFXYJPUUyupn11uDnEv+a5ZS1+k
4zz2NwEputdDU4A10OILpNtaXBbSkNJZ78leo4fRX+3itMakPd12sN4M6K+nnxgl
cYVQ8yVPhzvx8y3EngMXQaz7Oqj7qHiWgVlP7hT8I8yy0/AfS4J2r8660OejInB0
36y8JAurRF3XSdncJqnV3Wo48YwMOFk0C/OuZs5bx2el0Uds232DT+ITtpsN+7vE
xgt3lyEcumnr2ehWTrISydeSxlkCACgZWILWjDkpLhWOFwEgMLuTwp4HmYEspfbG
MFpt9ePIOfAwLrLDh79p9eYWx56piM3l75p6MU2RSoNs8pTHetrxYohIoa16Sz2C
cE35pk1d6jwj5pLlz38wlmTdyJud4uKjFtsje53rzDH/ACwi+lH3T6NrCYWdqbx1
8I65azeT1J4WeQBdl+5YTp/6YO6yWKrTQjL/GyGjo7Or1f+vaaUpJco2X5RPnmal
O19iXigHjO42KuwpZcWV5UgX2rhzjVAG8GnzQZ/fCIVXWw+HiR02gr2Gr5HOnqmq
s790ynmebN4nbRxQpdZMh6rT7LdYpp3a0UaeqeX5ms+UI4HxVQZ6PTfdfq2LaPW2
lsbzBLcWp0feluqvzsuRJjxZ/K7eRfyZjoIkCZOttdpcU5elHQZvpS1+rpGE21d2
aKEJbVm5MDpBv3/OT51nzrAfZFTv1rUpRdilHm3zwlWse8kUijGWLUCJ3IgYRrC1
hYVps4/x6zO+cBzwpK6cqNxBirFOlPgSZ0gMUiDPkEOu1m/kOeC0ms4UmBb3TOUN
H8lN1Q+5zNsMbLjHF/DQzEMncvSdOtvlGxz35zss0rPrSTYRyDKbnu9mH/ZUjZ+f
8jBGQYx0ZTRkF2JiPRd0GTN9zQr1Vk3mP74+UOE4VSy7stuCKXyqXr8XcHU3eHRy
5bq06O4Hc8Q1IWG9iKtv3sgrqJb/dzocIFsJmE8r1V4hODXX6KxKlE5oBLPSAit0
OGX1Je0VpEd6W8K+zi7CQUTjwk9i0kSQGcZSZzF3nIbyjvSj6TGlA+LS+L+G3uW3
dnPrUoG4M1b7DXstEfHdmmXmg5CmGzsvTRypefhlaJfQaMmBHnmvA3xqadEHYm61
b4L68SaPSvwJZmBBodsAscUSE6oOD7kf8dK1fA3qrntI8It9hN+KVt7esR+JGtrv
5MLsRs6Xh+A1WV92GQwYg23LJdXu5Jq+TrdoeK0JuYShxacXnQ1g9TJ4PRV9l/wm
9n0u7SrgRmvyijOy+AKh6y8WCpEXzn3Ut2DmrTAOAXntAWq6aiHPPRZYDiR9a8B7
ZDWULzGto9BNKRof2j7d6U+LaxfasM/ajnsuQ3M7nqYiVKW4YpwKQbXbVC/IINnC
p90vUCRtB84hMHRlkEnm2WSQjPHSWSuaM3xZqksCK6h9EHCB+0MyEYERY4mCkRLn
OM/0mhmK5edwl9XoGREJXyjq94p71kQY9Nt7IIGYCS8XRUu9kt4jwC2OqDT39EHz
Kuh7l2qMkXWIuvQ2bOUuBZHmsRSA1wAnf7JphcsrFIUSEfpKRPm0E7Fxd89cakcI
fPquqS81/i0Hmek5Mfsu/bTqHaghaja17Kjfxp63iCdS6OGk5VrQ65H0lrhXRVzg
PYJOalZcJ7cscY0GH9b+7qz2JLQ/a9NTYX5dQQbOc7T0+jjtD7Iuw2lU+DmvPaXN
5nrgYz49gbfitm00ZNjD+h4um6Q+9PhB0GR6dyxYKhw1ePvzORSaLqKApL6UeXGG
93sNEWE2HlGBC7l3+d/RlY+5hAjfN6GBkmharXx1hmLNsw2BMTYm+fw5Ik36NySq
4ewfVXcIgapPg++XDbxQSqmF+CZK7T4bQSJeYAXMuOjdCE8c+wayQ7HZLs4kBUgk
uLdl++xrhCu0lYNHkplG2D0fzk6t+QEcBkcrSzjHK8IEZHfsn42jjCDVAaPbm1gT
iKkcF9EVCxZk0+nCUdgpDnwl7bzf3KOSk2yQzAeRJdA/eTnnHy6qdbEtGDcXFuaa
toKqAacOmJbPniW7QVmJsvgX9fTNNqBr//VewXSjy86t6VJPdLvXSNAfigIwklKB
DgoL3fhvkjtscnMNmyZ1J81vQD/4L+MMNGrEhcxjnHy9oxvvG6x6PGog89o8uZv9
YELRrf+kxIjeh/CWj1tS2p+wql0XeSZJ2nweruGbRnKNn4bLl+cJ8+renSOC2tdb
2asMjkEPEnXgeU6UhEzUVc//DcvenPDSHzMHSuAfnQZ7p/RSSqoGhgI2hjIJ6B5Y
/3YoKjYiJUYD/btxzkF6STKn1AVI3RFVqDBB7/0sRJIkBBzO3SU5Y6YmBgYWRl8K
ROtogXbLrwMn4l9LWFAYwCIOwCBEjOrzzNqpheF+/pLRpYpDTa8hj7b4VY4X5VZJ
VkgUu5CwWruy31zwulziS9TEUaKmAR1Uy+IUf58foelf3wlw98wcfuzbgLt/X7yt
mdCVD8OJJ9BdsFLHwHsmWy2IsT4zIG3Kx+ZONb0DdbGWGvq92PFJEIwc1nBaXW/j
NASzjM/6UcHFzNPze5W4ySBwg44Eib0fAwWaTl2hkyQvZ7J80BxnZARFtoDNn08Y
IAV9bdtzGBlsYqfGJ+OILqyhBkfN+xXxP7vwgwZpA1Ymj7CoMbjS5msfN+H1Rds3
SHUKqtZHSG9oBi7Y8/QRWQ0BQVzmOz6akb1LuhGVsnoccH9xDzQikSCZV6PwkhVE
EFaSAUtK19ZAve4XJ95KGzFUlGHn5tVvy/I31ySZbRmdoZkydeWnrdW5Ysxp1wL2
+7EdjrV60nQ4bBEFSIIiHe4mH3dHRxD5YVqSK5h0SqBxlO34GQEObeDA62CA50Ej
fv5R8+SqRuXMGbMWEtdzd90yiDJCwuR6+ajmWJKW+egeiHcwrTv8QrO8ZJX/lCAM
P/z9yXQLRg8SafDu1logXiy+2UFzNKH5g1VUNBRJ/ibUwTvwxLBETJQKMeOSzokS
APGQJl4Yslqckf1zsmWl7C60IswjrZ6zTJmpS6Frfm1N7XRSsrP1DslXg2/VLqmY
21bSYZiy0sTR0EJvy9xnc9tMgC0TBo2YxvhOjRdXqsC7s50Ukuns0u1PorNmIlY1
oTjN64b2ODlEiMMz7nFVulRkjQ5tMus+cY/XFOrvRWchnWLKiY7oIbdHOgLRpg8m
AeAshFb7LVsvBTKRtw7xbF7AnAXAg6JNqCWSQ7BxCHuUtNVMwvC4+Rgr8rq958It
OnutDhArBfFb7fUfzTnIvxqMClOvhC9mSA/Jyk19R4Le+dUVyxwV9a9fu1UwMVFW
L4FOxBQJyagaI+/b3WJEyjN52FSouzy4B8K9n+1D//z6V9OH6RxOycqrGF83MCfo
SRZxiDdW/3+HyMRl6sNuaE5AbYUhBD/sxc/iQHDfBuFA2xJdBgtPvQNuFlZLig1m
wKGY4KET46yU3TmA02EGCG0klGMphdYVT79OtVscwcju7D7eQJrIuZEPVpC8EG0r
N2ItIJVM1AK3W3lperWPc0FQJCxN0RihBd5dCYDQosiRUmrYXBT+Vf8OYGK4Xbxe
XhG9kHkX/tQYfq0QcRfbnzmjV5UAoMOtVpUDX2xIPSCqhZI3C2IzxTymlvTmLj5D
VVHmpBfyhCHHlDG7p3gTsHPSGraIDPldwKzkmsATJNfFPxJwwscDkL4OwpXVj9vT
A/KAXmJtZmadOMf5KsRBew5jjA2VSD68ylZQFjK04PxfCkAHcokmJr+xhNV/clDs
iUL1/HISjzsK+850MsHB29yif/5ebDkETEGtHtk/Hy/12eUwTo+qiRw1xy+eCkxw
WMH1tOmFn93Xp/gYoW/+ZjUj3Do7OkMxJrAUQwGbDev3Sz/T9dDP6moalThHs5s6
gvRVdDE9Lv1endI1WcjLfNIq5Wx7s/PblyRGvEn9Xvujq9m0kzvMkgDVWBCr7X2T
iOwT+P4G5MfYZwN1/psva8Q9JCTwiIgK+LT32+mka97ExT7WNWR/CJ4NvySugMDP
sKyVe3c2uNTdKcvwT0qGDfYRB+zATEBntzrjwCZPefKTJLjehC5lV7CAdClRPC2L
5H6DgkwWysW+QCxogkDdjUNlusL+5uVqIMeQrdrXI3LvaK89N6ve9mK9gcSqpEfK
b0lC+OV4yyAR7nJ+uNoYMrr5POLq2U7rTQ4i6Ne17mUoqxX+fuEhmcvc9Z8cpimv
EpyFwxCWh1SCbfupfP+c7YSDYbhtJkweguHjFk8dEBJBfP665t/PuCDzz0PtTKqM
j5J1EpkfzH+JVqKQk+tEYcVCIPDcgeTsn4X0lHXfA77NMCxe3gCtoDRrNNc9Wt11
uTPzjulhwvKOhdwR6YwxarKczdbSqHgLsbcTApCvzgedGQxI5A4lKoROwVnRdHhK
TCCmkjzGu+9Gt1AMcz0/mEncaD3CtoWRHgBMtOaAHhcq0HZueI3SUwe5V/t5n4Xq
U1Fw+UPZ8NqDbzRKeAPqKgYXPqchB+oA5kAejTZGO1zNvXA8RCdfKlYEm84lsSPS
yXCsMtRCceiU2hkXaL0f7yWUzD+NTYKqWO/yl5BvO43uuIEonYXxBxwFNO66s3B8
d/84YDiz85qBT9yHYbsZitik0bKsUKAmEfMsqv7o3PqCIxLZYZNoUhkfO9nFImg4
f7WkbyATpcTypaPpzxPO7hkV3C28lI1juavN+5Bhxe2DdnWnxDuz+WiBrVWp/QYJ
R9CxcCl1/wLmVcCEFJk//SzaSvONEdRuzFPdsYhLOltpvcJy9jlCVryk4xwqcKje
UnDPwidKVicZkLKEYWL5YVyO7oi//0efSr/hXYz6FrVpDIrGSIy2LQOgfuv0vx7D
rGhmgXb3sFrV7ZNRNtKc1C2v4idAc7RJH02TgpQG1gmD1QQyPZGBFyTNOFZtljXE
w+GxJdYQa5Qj8nU8MXxcdiyiEksk/j8oVMyFaIKcL5RzpbpIaOQ1ZASXzvBU0k+S
ZP+oXym6dEwGRP3rc/7FP7jK0WA4lHMpWHq8iLTbbPjXvsVjmaoId1KXOUrGdACI
Te7gzVR/r2NZSJR/5/VKB3AunwBGSeL+OiRFT9s/cQFqJSM8C075aiIP6GvN0zls
78wCImIHtRrFZxjnw0UV8btkUlyH/809pbmN/Y+FLAbl+QNVmlU+Ai40RLWRm+7H
Xaxrjl4qfaRhFpo/IN87Fmij50HuuL+upNwilZuVxe4qmFyYlNR9zJ2ZOsKeoKDy
ji6T7vjn/8KbsiOXusVgpmQCpgLochppNPJ7vKc6ASl1K3yni9F4xBnVOaT0qUjX
W/R2L8jnb+6WjG0idke04lEWjRb2glk2GNX2bbFCHGXehMNwqA71mx7YQiW5d+5A
T2YMFcmRjZo5jzbps0Sp4p9pmESKH/YHSO4DTM46fycgWtaqN9smr6mRS8AYiF3H
HZzZMEyoV1DklYIVPZnAgYElniTt/YBckRa8eBAsDzSAPRO8diNUX1t9isMYFnnw
3EfAfglFKsT1LWFTK7h2dI9GFyEW5n7Topx/X3wlt6mXvpXHLMGMvER5lVfVc2Qh
5gywhuIjQ2kIwxtmKPaLFweLvz2YAA7NFJhYkHjTT2Mf898bnf0wovRFdo44H1yT
osOTAvpvuUBgJWmfhdRfuURfW1pfPhcXlakkTlwZQBKx/TffksT8HnXAFmhxhD+R
kHDLcUZQWkisDWCC0M23QYUv+9L/30M7osnspuJjLoZI374QRwa1iUDnVMWSoogC
v6btHpyEWfFWe4dDg3ALfBejwFt5o+ToIldJCp7elIV6KtQ3P7Wo55dvUuhp9vOp
HjdXDFxm/rmHWKfWENrXogb4KhEqkESlb8GuP19G4URzpdJX7d5j4I9vcbWe54Nq
OBEHBJC9Difn3R8k+sFr5b6muyPddAymVn6HZPYq3aGgU/1VQGe8sKH05KtVxcTM
PcAN/1d5liByCu6yPZrDLeDdM2V9ngzw0gXgpsn1PAD4BOGMy5cwAG9DDjgELXlS
OyvnSLo72GywRIk8Y7ykO5SEBOAylO08lHjKfuluF3k9fGZrMfh2y+wGzylZR4ho
qTKVF1sDzeDOVI3QlpnXo+bHngJDruErQ9dURBDafSB09FYfULk5kPjW6rH2W/FU
4RaC2Hf9wQR0Qd1Rod3ZuiF3hSRtOwVCVttXG0OhiAZpgFfOJMizUqnVp4lV6Wiw
ReE54IdbFL5rl5o0aicNyJpmvhjOVtbLzPs0oNxMuJeDmSjIeziJfwnH2vYXt+no
5iN8gGxsbVJSxEuO0jP1iZXDgfUHJ/7r7sqUMlPTzn2I62fZcGSByA3Vmk0FDPBv
Df34m4QiXyh4n5u1l7mJQdGHdJcU0PyiOdVc7MiAncnWiXcunwMsLI//qEUfODMK
rnrjPV4lvUqbiUoEv84k4qqwWBk5fUz/ODGHxVk0AJ719KBVNRiXbGsajHhANj/S
0vn+sQDUx05nJ6bW7zJeDdLUrmwDeBYY1AZK4k3iQdAkQjkq6sR7JeV16DnBOjTS
iepsjLHnJ1GWsOof+uJ0woSS5iTk9x4SdZiZXAMCpr4/fx383u2BFJ/QXAPsARsg
wxANYXQbpqt9xCHHwRqL2rT4h6NH17r96F0w4i5tec43BFOreWgFO0Obi2FDxU1V
VMKKlPtFfiC0KGfSFUd+nBPI0FNyaE08GWxek70H91v8yQzH1lVD7F0Ya/e+eUKE
BYhMH7VHi3IzpxfNJ+PSx2fSFvkbXQpB6Fjs8pY4C4uU5M3nM81ubUc4Zc5nz2sH
BEhLaMho7nE2plV46H2VJGMX6YM/BKBszuVRxxqQH39gOwbEQ21RkXVDPu1ez/a/
4lwZReXdU/jsLhsa5zSA/vbxvNkhI+SyAlmH+Np9UMF8MvIte8uchBAPDA+SPocV
yULiJHPWkKnGxUpfV8X9oboJ6tKa8uQAftBDdYEhVbWsNsQi3OhY3z8uukcjWL4V
K49Sq5EDEntGVi2jUHtsYRyYgsvvVFevLnKiVHhtKsz2S85Fuf+TCo2tlg89sby0
mttBefO0Q9eRn7AYdXiW8oTIp8i4p+490VcRqmk4bfh3nn3e0XkjSsZUM7NLMfRW
r5d4SAAILzXVighoOSTPA/CntieFp+qfWtKQUKIH1mB/0+lSlt7hOp1fsTWeZfWf
oKB5Ayq2n/RiaDlM1oqQdZhQ/pkSKPsH5pe40nwMKZ3vH/lQSHlJoiP0dPGlJquM
7h6nBZ9WCuMjH67AlPej4zXkWDNrUzUgqAi0D1X9xBjrGb1PzFcyDgLS4pYxr5+A
a66eoGkbuFJy4nPU7JUIzJmHuyBQAJmvdMbk9/fhprVTDxxcTTi/I9dBJMZMJ8xQ
CERJibdeOkvvs8jMsf5ygrEHcQ/e/EgrIZ6pPkd8dkiHcT06NVJ9pUBH+a9t9ous
Nk4D3eCg9pArwQsJK7rJlewwTcUzSCfnxHFB9VQMStj0LbWq+pMjJkf8P0jpmLyx
maQFF68KnrHn8N4aj2xMNUD7DQ04VJf4K1InlB+kryGupA+UA8cKxIvqjrXZvvBX
G9wQoeQl2x+Ayn+Yl6ickLZOp7tBGMiYSloAXfPEsmSIMWKLnMPX7DbEMkjluYlc
8zL+ae5gl+/9RdUmgi5S2oDElRwaDbCU6g8GdVMMEKZ42IEy7s72RMsFFllXB8Z2
k20GW3PYMP/jxMd1bbVPXlolh76JqCVb3vbLsqKUT3a6b7hWN+gGZ+CTtSgZpT1B
/yQDmTI0Lp4fDyfnrijSRa3xm5NRfIJgFpYC9ZkgoYVNMQCir9oaPlC3hVw50/OO
ah8OTf5DW/56XCuiDNEOrEf0V1MSg4ixwjcNkiiWx/RNIEM0Tw1UBVSK0S4RDdSF
kOotfoc83eDaTljfm4HiNAx7gQfgzK5Jkg0itla4z8uDsKgAY28M5TdwzjdXmwtr
+f7iZnbC+echlozxULhAhI2fkqXe3NVQhgbUpq5x4Zv/jXCu7WVNwwMHc7HzB87y
hwjdmUMjhUOtwuXun8DP1HJzmi1TRjU1SVhvNkckY/8XuZiC745STODrBJa6kCXD
OkgtvV+WazEAuKs9ZFyjglijC7eI6Xpt71YDOA6kS4LcNOnCwieLZ7Ya9H56zwOe
3rkzva4q7CBvWbG5bEIzmwodmZjQ9YQPN1avtZ3QmbEZcIXc8I4lJ0kQHLEtlkeh
iTIlV3fLbAAgIHzxCTR+PZy/SE29e+8Hh1uuH3Cy5EJW4TpESbZZ9NI/rbNPe136
u8fheqH9C7echHAmqJiPC6nmlDE/I1xorNNzHQL2QYmVR8uQfLcSSLdinixL/xHm
JvgpbVnIDOcyj4pUn22h/a7pZQ/X+CV67LXSGBzS1qZNkCUtJHv/CSNCFv34R2rA
hTMc8ByLNv8nsOpr/MBqvntQQQpnbr2MdrlUFMfKR1C9aMBcJj3RPRzjG3oee6q3
Zuu6tuaw7X0s+GdLyf5PkPp9DIPWR4sWs+TgzypIIUFjG6FrfnBprwMwbXJc5b57
3AXu2g5MEPEe2uXpAtb1UK8yz0UjIb13eZ+7K0MYyeM/CQkc+cTuSaNsIoDJcjtM
MK2lmDMNE4CgiQwxapqJxhnlPZzQ+6cWYwl7dkCd/CFNU86bIBC0wzqjq8HO9a1T
bYxIUFQ7kUpitBph+B1arWpLS8rVb4Dijcpx3A1ADsn65r54XkznFEUWspKUIHh8
Z3EcgeVXoEsatuLI/m7cRDu39bOFoche0xPIuK7ah+ZzGM4Nf1diyVI+scnfOkML
vf+4yQ1zB3NBhasnouoqdr7pwGbOtFk5pvla8YHao38OyYaPxLYSUNskIIjyYA7R
aQ+QpMOSx55Qp83cnV5JLe+24jIFnxdGeOxELivlQNryyosQVjeAG0HpH/mDBdpq
wvLbLrdHzcmqjPF6wHQ8emtREg/rRsUo2Fcq9OnAR5WeRw8bK08Iy8v4fwtrDZC9
ZuV31n0geihNz1NkinrJutQ+YBg+LZGFSCueCrR4CuYwdvxoumClznOIrQzR1Fbf
a+2j0fiT1jCrtKh1fd0iSnDvcFKIt8D3XUdEwBjgRoVK4ArUb1/8ROdhAUv/KIUV
3zlprBvFJycVxRxw4VgTsxsVnBYuBnhVbwtWA0xY3o6bE/R0BLfSObtseZZa0x02
gg5CC9dMsI+TA/B3mfVSnRHuw90bKkWYpuicZdR5Za49SqSSv2HN2+IuKSarsRfw
3Zu1/aui1hGVEk4lgb6ubYXh11GYlyX2YN7Jcy/NMHmncZC8q6fh/yTonEV63r0v
uEKC1UPkYt54IMoznQ1Q0KkAnLCDgCMSbAT0rNladriEsPA2s4Wy8siOS0RAJ070
N6HawmcvpZah4xEEYMBLoNPEAlR7KKYUXiTnDKJDc/N4QcthewggckkBZhKNCHaz
OpUjhgLXCe1gg4+sychsavaKwQcxY+5YCASG4wMnppM9Dhl4TwXbkutvWGMmTJir
6dvDEW57/hTzD1+TKzwkPSrpxXMs2QXgSNBtpX9uL3cAbaTuSMBUxv6fMn+cU9Z4
2Z94sGMpznluUFZcXrp+nmQTsezSicC5SdOOdWfyVF1vm1x2+iAimqr5yVqMIGGG
8qdIzB27kljO/xeDT/XPQbOlba7CjELFUs/Y2OjnT9gq75BjRH1NlgeOInRuSVyw
WiQSWhiMDcPhMebd7/ROJDU/MSyL1sK2/M5NqWduLDgOyN2xQj/DppK++xsmLbEG
GEr1fWgwBzj48kKXLW5AOJN7gpJNKFUANS/9LlBKWVI0WBZ1EGOxNEpqI1I8jU/1
6K3SKahQ6TL6ZzgerDrQciRanuePAWOKddaTior6aWR07IvD2wUzSUKac4LaHy9S
lbtfcNJFly4msbMfE5Yng4O8Vwo6OzoZvybaG8aGVRp1udoOpkSeUqXSq02Aao3C
Bl/O/StjU8srPTxl97mRrYOyEd06s6pK0lLVruzouryJbawf+FsJd+r1rpm2Jhu1
0RJok4S4aSw++lPcaxTvm3oEqhiU4u7c61yGWumqX8UZRRb5MmzG2An3VqUbJ2FU
kIr2q7bCZ+khTy8ldJD3wUhPhpITzZtHUL0y83OfkcpZzR6nLe+4SQazoAB9XY3z
UKeZeHzzKGKNT14f+hhBfZIUbNuX5XRt49SGysI3CzQer2+0NJXFMycnOYhfLCwC
amji0ub24WS2+2hOCK8KwVlvYZDfSYG2PUCiEbq0JsxMyVDM3MgFF3rRHfAIZibv
cdxytOOFgYRBlYkI3NGkjtl5LAqFyiyaBTb/cABW4GfjdrU6vYD3Vv8RS3yA/5oc
NaQmrHk/TkYtEjhD1uoKmPjDhH81hC45vhBmp7+Ij0uFo+rZ6D7DIeBYw4l3sdV3
DCYwB4YPjxbDV2dSbEWlliIph70NVbWxAr4B8xKIQlvEv4Bh82+Q55iDFKjEuwN0
iUi4yHLIv2IpKxZj/ozmNI09W3hS1MGcxJX44STkdCk6vxNQXVAWUhzYqWxxGvTW
38AgnmKLsbpa5HPQDE8EiNdDAJ10kDDKpt/1mmucz5hnYL8JO1CjbGA2IXfsH5yY
bDkeHeGLLzFHhlh0BVOBxaCsmtGaXecvmxl8jOZErogbzsz8AoJep0rPpRk1qXj1
75UPN8I+mD78xx9ww0h4jRaBGI/qFYL7vTbSRz6Z23HoofUCj4B8RBXcniOWTe/c
cO7gyNiey3uk3TnghGTTyb+hPxpP4m1oZOt4j0Z6mqwo48hF6sfJm2E5VU6dTaIG
wu6pFDnROYYXQQYyg/Q7hDLpjS7Ia8aGKcysm+xuOErmx+mFo3OUqsaDNlSs3eln
5/uZYqBbU16UIxJfKT0e0E5UdB3jpPvWJagRaK6CACyfgkmbc4ESXnRL9wlkEmv/
Tb7k1dJa44plzemnrV1t6GicUdw0KutRgs1zNsq79pjnpLAlMAQOkyCNnJ+lWEWR
979fAn7TvQ+pSxLuiEegkF7W44XnZpDEmNPJc4v4aKjw/8qmgSjE4rMvZq/Vyv8r
zmgI3PB/rt/MUrNI5yqMlq6+iF+EXOFFlMjdeJJPYnlXNFBoJ1POqFKniG392nXy
4Lqzz3V/fsKcCFlVMUZo8RFKoIbkR6jWfu22WqMpsPqOkbqVwEdkmxuPWC1M+x/h
fQlcgjON6oMkIdUpnZJBGENjhEVy498ABV8oKoA+W3Mi3KEexV2GJkdtFfqkXJke
Qn3qSrHz66O0t9FTLSs3ZI5a0aKKXz6kCM4klLxSHPGpaf4iig7NY8ZXRIPEGfHW
btM5pfIcqNq7NlAGHUyerT8Ax1fkrN6yYhSsBM+WQOmTMU3dlIBqmKdp0Ck4GpiW
qbojVBo5bGiJkkeXVdk3XyOTP1/dNaAd50f8iZrirGO6lDgNipUMf/FUe7fKrp5P
SigquVKlOR0mJTQxAWQijnpRJQvqx4h/VzD1D0A53NcIGiuUQLtUajP+tdpRnOx4
Cgqx67nWSPF37+ntngdGPqogrM7M4hgcBNDUD4PvOjkNhSYywnrFE3Bck4oJ/DoM
QLASRRFjVSMaXifoE/0toiBV7gMWqLwfTAqWc2FWrtJOafdfufDCEof3Na++hf1G
+RPVwdYCm0aD2Vqw2s+gZAK0gf35eom4L8FBIMAdZ0lhnMkTpeshHnY0agr5aqaz
2HO1+pM77Zs89uhLfMMVqr2iBVGEDhokFJFdCBNtt96yIgn1u3qozY9dzZlDQ+sx
DwxpDQQb3fDJ8/nn86no44+zjMd4EYyW9MGd3feCKbX21gabiN0q+4S6HyCNB2j+
sWK0cwAi3ni7jp/z8aYNcvnNhMtQG5yrWnnwcNryKE+3sWLQsklCD1GHhGrElp7f
4WXLNM4AevlEWd6DxETvo81EF2N9KbUZIsT1dpcFiHkM+kz0f9KG0gGMslN3eGJp
cOvlA8G2WTqdih4hbgYax9uVJ+e5ClamrxNNvGtxIvnzSqM/+m5R+KMpHMaDiawi
/ODe8RyIDFFIJFm7KSR5dgEInFIWbuqzy7HyxmsTAHdto8/ME+uwdNNpoWm0/GR2
FAA3noAD5VuwaYu7n2lan/vigi0+vqblmSfapwG372gZO6q335kBr1CQXxAnO1xW
aG9OfP2MuYoWvMj0+2A5sfhD6mUDDWvaN4mWggd/S4svnhvlOuP7DtNQHsPJsv/d
w2TsyVrORZ5KJBjjF66L57zATPRPSYljOLSUPz3Ub5gfdMAq57bpqeZ7V2KbPjZm
jQ1wQ7HsNjB8ZCn8VxdaALQwVxkLefE1gq/609MS29l4r2LD2tDUeSDVHJ8bKtc7
8j/BCkhYN751OfPNFZ/QPV0JSXNGihuRAS+iw/yJrGHZedU88rHBkfMYwBwnIqCQ
QzPH2gCs19cuUKqeec2ZZmrTZOhP2weHHLFiVCps4lqd79IrLFliO+sVX6B8xfwS
x2t6n150kj6q88LWSHlgPacPoo9RTLDk4TMZGGEi3zNxn4fJ+RROSm0hhhRkr8pt
6mmA18yfQLPLiZsGVqMSa+qeyMYZ0Iypjk4rXaLqa61OxFIdHq5Ok2SNplwzX1+f
2agUU7N1R0NTwoZ1ZwxDqxJT1Qb8xcbXeJTRqoq9dx6jbi4jhXh9fAo7cxj9L8RO
6rOJyDlARPat1V2CUqqBHDZ7henMSAGRVR9JtiVWg7juEYaoPbViD41zYl4pDoPB
STURVjEdIw6juZa7x8vuhi0Wy7aDRTZkh+AnX+lSnrzPR/fuDyLE3t8wC2RzsJB8
MXl6hA5ozosUoRIWmaRGyRUzmzczNqJGBa6ypt3C78WNpTZ9CXJ1KaflAKcLIDrH
6hmBKwyHXn/S7w7foBsslNm3qoCABw9U0bNzs+EoIHbJmwb7Rj3JUphC7AqqDgGd
Og4Mt82BKzKa/8Fq/YYPN7tNZ4ToCHuwNhqZnY3H7k/kuSyRd0bEIw+uedGVvFwm
PfekjozA42bdZ6XTfWt+Nz5+pxB8E+8g+BvltYxnkT6uLuNQnqsb+fIOFDll/CBf
DgvzwFUEw9cF/Yus+rbQWoLarOzAuL+itnqQ6Y05qnecSJeCT9srN4qOziLCIdo3
H9ChQEnV8dfjC/iC2l4UsMBrA7cZyiYGjK77CngTVCnnq0IqJGZyxC6OJIS2PNYE
vmDxu0pjExG/MvDi7gngs5c2qCw5gvxTVE27Y+VlQhkBMWpNM+MX84e/h/q0zXeO
MoNZl9i7vG5jwrm/VX7HY2x428xVVzE9ddZrv5dzxVip5a412K0YzPGChi95ZqSH
vNx12dVafGimQyK0+AamINv5s1aOmGPlByv548w2/0Gjg79BxA4KiZqobQsealMa
gnD/iEPpoJyT8JejhU+RhFznsmLTR3orjVGtGVbFWJ+oJ+M1plbjlWIA1xI2oc1k
aCkklvR4iyzpjKOeSV4i/yTrHiN/nOy0NKfrzGzytrdtCKpDoi45kv71nUXer5FU
8mjyZwh8PTNNDb68C2BfOzTz8V75u9wqObqWEewEUFwWhfvi9pn++/J6Q3pUXx9K
p6xai1xBwh6fOHVZbjflBsWnsMo/H6sfRW3t5QTMnOA6rfeHVYZ5/E6W827PKDCK
B52++ZB3jOcxNTeJqmBnb7GxqFhhwFpQFwJKRLcA0o1YJveh0Jk1KIkepZSvsxVy
/nyUZwzJIiCEOG7hoNEDswndw0O/idSmC/SJpDpzuIaXuK8mqeDszAiKUdLGmtj5
M/YWM8X/NojpqmxJ4hp3WaaJhPBqwPiaobDnpxkoOElbXYKz1E+/2YlIssFT24Tu
nxfouET/+nRzzHLEaSmH4nQBWCHLhc2Mchvr8iFO0CPa0iKIXA31u83YMwfuRxgf
tZ7rNQaUo0e9FJdkkTVAuqtkTNBS9TpGLu3FtaCX1ifcsgoIhSXx0p8RQyGhCYQX
V/ot1b+YmblEg8hvD2fhpt6w2N0p66PMXvXT6OrOlcdqOrzpggL+7o0/Fqw8WwMV
jfs9xmWaa3zAN5TkDLLGEL+WUz5yTooNUKvKRY4bN8MNNHidRyU9LP1SIDxEbSmV
vxe6KDQ9RHoUfoULTS0qLf8LbEjdz4EmTZ3lSAzolUsfbXrhz3uHB+UZfGv2t4iX
jQLz84zK6twM642U9/7yEzhHTb/0Ci8/9AAuOwW2cluEfyrh73WBShPVp/tc9Q2N
fifSfQimTWehn7HAYIp5KTpEg2EyUnh9immX6S92zfa7rd81ZoKxl2cuE6u7eJ+F
oMmDKfDmpdm3Y/M08szQ3MpRGjlpXcbufJN92NEQ78qHPVVOrn/awAZlLDlmEa4B
5Mf9UdrZPzxPLFinsNU3BmLfwDUXBZkjVkgya+11ePAgnmi4oEAzdhhG9HXXMSRb
Go7K8CBv7FVyeZyollDGCvOPYAw5cQVl6dMYcVWc67VQ0KFO7HhqEn5UtWT9/HJG
8kOlPuU26F4x9YrznV159Gs9hRkNezM1YueJpXpU4umYmDQSqpxnhZdguolx3+D1
59gHGMqW04vy5uNLAowUdvLzfjIFLMAaZvZBwHdkSp5MgEfwplBJbZbvtGmgAqu+
cVnonNBDh3pPcdSS4wemg3//fChg4Cu5jDN1UxZm78KyCmvvdPVYjOXMvxpIo5fa
5FMo2GCkcVjF51HCXwFWgHbGkbX2SGtGtP7sX8hoBzh0VhV3jy/IQGxi1eTWgudY
Nx0+7tsSrxfsdiMfcS+0bWeaduIOSrAgNru1vg+VxNh+uLVw6yb7a5t6eXWrElgu
4dZDVAvCQ9uYyXD2QSoKNstfAI5QfuZHGNpRUSoyjPkwX3k0fgIU4Edkl1+Tqxdc
m4UFbWrpNsOlteHeeskpukUhwPvq5shpBwoNSy8+O5U0S8PP4/J5DxRMIoI8B/kg
ytXikq1r4BSx2C67F85+EJpE9rhj2Bd75vOotq1n0xhNbvWT1xfMP21P+bwO4NvN
R0ZcSc8lJpIXJ1Qq0EQrSvvE0NSZigFe1rNsrvx+tpwRtVFHCWn/mnz+BonuIptL
RXXDxbHKfGlhp2GjjV3AhhbO2QOGxVe4RWFzwy7FCsnP6JOvkZt+PCLlTxCDs/VD
1KtMIda9ni6NH6451xhSgQMrIBGGciUn7/LK75f9rU1cwqX5RpakIt+JLC5ZndX9
qYLbcz4z1Ig/KvLIznwUTRI/CILJpi76CtcuCqcPAou95P1GYInz0hdJ1vMopzKw
jpfyeDeGDsNXGhSXF4xrNOckix8Cc/368/Jx26f0PLqgEnK+Ow9GhuQxC6HDzYbT
3gWKTMTB4+n4n1dBG8V+tgv8Txyz4RrOF8NTgeYkQ1+MkCrQ8ecZkurn++t7gR2L
Qd+DcNeZId1+x2NMcQyez+ECRIKhKe06wPTJs+rUvfDQZn5KuKm8q4nrnGlK2Xd6
2yucrqpEnCydwVmKS/jD7EJqQkXDBYbmAbsOQF5BsOHIP+lk9Ak2ZWzonIuEdXSk
5hReA61mAtob1CKVAofnIMOdglBV/Z1jlPoOcLhe2PruG66X4yru4DltLuqwg5Nv
smngwFW8cSckLzO2ZkVh84VoAGAQqB4/6u/FnHEg4l9eqUTjQAV2r9jMM5B1Ff1m
pl+wl2OxcJLYZv1nCcSvSHjJ2dbKqO0Vj1MnC1h7s5MjD5GJEbdWzffzrtrKDH0z
6IzvGPYz21gXNMzB6TFSjfJHr5+TKx2+zGCvcYPBfKz3lYvFOCGg1JvGZTia3h4y
yarjleWT+AI0Efr6PFSPaZPlMPQFgJV9IrFtBRynKINaGYoQ8dREU2/C2DKPpt1h
9XplkESwbRPDAKkNMpOni8aOnyR4qzBYfhx+DOe15hLdtOgMLd8wT5T67gDMZbWJ
tnS58ilQWSNLetUotda9d4yx2fia5Xeetuq7Uay8TAgNXzRSrllxEObNK9AVWDqy
2q5e1oGjY2howwJ7Add9hrqm0msBxT+dT10BisFCQyr4ujrc6baRYiUY6IgdWjil
q/YdtCXRDIu9qfnOAaRqUVpmyw1S0tOxG7XCN9kbaqEl/Tv7T1M/0iLWWflaQ8HA
+6PGgmODzWd4cTGpH/tmSuklXV9/3vZZdElxC07Snk08wF/jmwQ8TK4iYacUInmO
0+tXI34gzZAySIFRtrrJskJ8MdGG7s7dBkEoWXvPl+WKFVDitFuSbKg63FwF09XZ
pibRql7pFf98TzK2bzZlDKimhfWffAvSEVcfTWA505jTPW1oFkMEYOWjfDJbydMs
BbUwCfu4uvZx7ptl1p39gaHVsc+6vEEwQB1XQwTZ/n0W3IxrLuq3AlZBtjVYgp6m
ze1r/+hzdATuquf6XYF8ulqqxmSGyYQYOiDiI5CWGRooGn3rxRaaUsUWj1IIZSsP
pZNWkSWjdEyjtQD3laZBTJ8mATuhWgc4282S40O0UGuf9e/Yw39r7MvkCc2CaCL3
3/6GCyxwoPZE0mjjMnzziBdFlgTHDjeQMU2UiMqDjcd7CcRjmUWbfPQ2ZoZmOaya
fbclYvTLOwkyGBiOXMeu510oVgLLZFjWDyqDWUMepzTsrWYkP+eFpOypIn3z07SV
sjDlE2c1R+H6mt38wMd1LOCNU8Cx1yY4via5Vju+yn14EmGjjfw+y/Q7eISeyU9/
I4Z9QvSf8IRJAxA2XT23BSwdSLulYrO+BFhn9GlPmqdCyM343mE0EpYAgINyIdme
AfeDh0NtIiPOlofy3kRcC64HHocfZCtuk3UNC5996wqrNWqAJaTmXBgsO8xSpWgU
psJRzefU8WHsIJ59goEPDwxYZGB+Xz7TvnwWL9RTiS6VkaZt9IGGBmVpKMFZfy6t
+8xrMa6hfejTcx+7WRj0RzHr7SxcbJSQ0EzGV5EvFjoQJ63SukB1ECQEy3KwID5E
1oR158ABwInxR4zBXr25C0q7fo7lwsUuKDSqe9Qa+2z/YQ8iW/AYSby4k3gahJ75
gmVbBUYZfyvHP+zdjK+L2NDt4a1iKU5t/l9eUtvVRDU5ewXo/f78ZcJxtqR+BajR
PBbSIPYlbFb5Y7To4gyBMqih9GqTSF3nNwPnr3LEcScBCWRL0IYGNZtMc/+3fFKI
qWYNLvP8V6tQwhQK3ED3TcFAKIhGlT9GVcWpRnPSiEOYmj7GCsso258qNiMMwolz
6+LeBnwMwqHQ6UZsfg1RjQ3cwGV/CM93xtWydBVmMFlhr8aCK/qMGOgV0o9fk852
P9QP9GVTVd8jTzQCb875ACLMbkS2j0Hw6LkHQs7Wogbia7TSylPBuFtzWjA6cndn
RL4y31/56Od0EzDaG6xN1LW4lSmNY86sQvYCe5OogqCDvTmq+pF2hKTrP4+KCwCr
CEaX5CbTwwf6U+FP3M1pj/nJq5vcj6998l5lZ5P7rTMhT/+nKTQYmB7H+ZfuT0F0
hX3snGwBYkEtQ3VZsfT0vumK8hQHZ7iwHUbfSqOtodq5VmNyXZHEoYoMiCnH9OQy
+U0sHqZoDctMw72SR6DmKzjGLzlyEjDv0hz5JpCIdE3APT1UMTfviRDG67+kwSsK
jC4Po/3tZ5mUtgo4i5YojcWJDwVIZerfFYktQBb70xcsZ1pNYYJaByyDJo6eFPt3
djHB5D8PloCmQk8tUmmpj2f83dPeXCfkkVgMs/8AVHftaZstrHYotecmSjuNOocO
vscHuy0/aANjHPvb/fzU14kg4MiCGlWVq4bx1xPN2Me84GCi+bdDw2/CD3OBBdeM
ajF4EfE4LqjSRo4z+7IKxWRvKvKzTZrz2bIL4JbE0oBWVcdl+Wzxrtt61RXHj410
Cmdmrd8I59f7AKJNTktaw/DGinzi6KsEFTqNd+eAQMLPJmdI2jo0PNNJLEOOtMIL
lxH9900yAikyb4qij9yzXGQylMhP/USDH4RItoRxmg/FEuUvzaxMDP0PEmYYAcOB
OZp/w4d+gamOe7X6ZUlbmrBeR+1KKz/7iQnvTI5RjaJ/clqqA+tdiJfyu9PG5i35
Uxgnk3K45bjgx/Wu1Tus8xWbJRKVcA1WaicEZhuLW9ahRzUB4sZ9A+iOzijzzDTq
AIML1ayFJdDzQ3p49jLUaCSJ6nkF4mIaT1xumrcoNKcusFErLCdj8S6rhifMfPYk
NhQdpfyW40BM6Dfo76hEKqSOGsd1Qd0iTxMPkMTJ3Pm5MkbHaFkkfENO8KTxVN16
+QuC77K5EZoH9MuoivMapSqdvRARlyvEuizG5X/AFf+/c8B7FEpfLUj7BOGcTpWI
4mGbH+OZJhTs5NBSWZDNQI9cwi6hW63P1nlZZMjxlevXV9afZmm9a7qmwTqv82i8
U/esEx92WwmdSnNoMPENCpfpp0b4DhHNe++y7hCE4f0sCyhHJkbdtgpKDMzUkhDD
P3gzO6phN8DqZi6hbWFiqrFy3IpWN4SaeztBeEaayp/EZB+a5UvHA7PPf9rzpkFd
ASs3Oga5VJfZvLxtX/kkFlPBYUNRXWdVg+2vczYjvx4f6JoNMSqPcqzOtr5Xnz9n
Ola8bv+sEgGGsfIw8B0a91YVtaNlepQa70CtZHA2FX2pGDdxZuSZYSf/cLzMpFwF
PWehnXnz44/nONsXK7TaXTtsMAaoYdfPL99g0uCoXaxKB+PINKTjdDI4lCqIFTEI
iVcDFsWAmc55F9KyhSgrWCaRepVaX+Q5X8YyvyuLuaM9PaCT8lDrPa8Rt7cOKOG5
mj/jD3TrGTcKxHnrw2JQTLDAwvM0h5tpoGqAmQXtelNaoV80K62/miJ0GuOVqcbY
Sz4RSaRsOFouzJvkGSlkGXliwGl8qt5KXJQ1WoinyRQ/GCDcU4t7rSvTptBCwpT0
f14XwhM5l0H2v6tzJ4EXIE9bn6Bk37ad82D+LCpNzeAZkT1VRocgqixT+KaA/m4N
hShS/LCcFO2iLaxjIbsPPzZbc24SLXjBLctySOv6Lrc2oJVAeOR9919ywnF/PiU9
XqgV/xNW0bk/lUrKPNbHJStiHSRa9XLYH1N8FKmjzQ8z3E1ENBzwAkhK9hWBvNS4
IOk1s38h82i0aheE+03VW91363GGjrBZeySUH+hzGJEhCtr+0mi2rQzmuOVKrQZk
kHw0+tNumVftAmNnXjtFuxgZmCYTzknQV2ftqsZ7r19O053k+VUFBdykTxbLZ40y
mIFtgjxqb03g2xrrcE5vPTqyNxchELXu92Pk2aGKmQgI9G7Py8yOflK1hcSbUQNw
XpYz9STxE/+qkUGcC3SSoDHlv08mVXbId2/iL1YvgZEKDPu9DTGt6AB4AcPwWi92
Mj1ergEyGflr4LncDbLcLASdhHs1peKOy8NqmmgIT8R/Pfk+HfN56XgTQob54ZCN
5p4jnU31y77wxXd73Lm9FAxKwAepk+oNs25BmM7cdh8JktNkLJe6bG1G2522rARR
QilwujjsmpuIrHW7w5cZXu5fgiAL2VWsObOSMVE0t4nscwNhQDJza2b1sf60XKCr
Z/vUgIB3zPGBOPSIVm0APDqJ7HzMysxLSTMCCJB4CE++qYrYdoMXCO1WsBZ1AzSO
O5Rpt2ZLRRN2LAsR+clrefVHam1B6frWTROkRgU8xCeDGSUndhLEh3YprAW7nryQ
xC/cFC7H7kPaFeNYxCpPSkpHhXIXikatNV/NPItoxterhrNvQl84H1Md866F2Rmo
SReY0QX2ma50eUvq57WN2qmJTzdHczkPD7U+kKFJOinDlnZ5mmaXIj02mgfw5hXB
Fbj40p1vszgvGzr4ww+N4zsSGq/GmOIFpSFMV1H83HKdl15qCvgeU8yzwZztOTYH
fA+h5PNFB/F4EWiZPUAirBVyVUqN9awd6Ik8k8UdPa6aQl9xrLKo/X+zeg+V9CUH
hCHK30nPCsU3OQsIsKTWnZlUIkpTZ69OFG/BvhCv6UNy0/eFGhx18gR91DD4O/EQ
x0+/8Eh4WoGi2NOwjJCvvgUOfEYz3RSShTv+UvP8doGwQnVrve8II3XtRE6QfZV2
xa3t5+zEesEBz+UfXwvJuEU9pJIKo8UFz8+nAI/vCbashoAYLl0bln2Ezy5awE4q
mCfisX8s+YITRMsgG24ekrFilJtZsIk0KQ+dvr0VXiUObXkBRZz60ki8mt36jpr5
2X6tedebAOU2gcUm2tmuAJFkXuacoADQSCdpz2uS94xppRw9swnseKl2cgvSrMCl
nBwGr3jUw/qlh8PyDF9Poej6L08s3MQY26cYxwVFVAWsNi2Eg6L5bvNwtZL2sjYz
6X/Q+7pw7Gk4uxZHoSGZU+81fnDvkxoS9yoSsmloH579nSr/yfB4XgPYHMeEuKHr
108hxkdavQ1LcxCuU9b8VcHcByiD6xWyc3auRKrtJRKaM77Pa7TF/+AYr+lNpPr4
SuVmTPqVGvEfD/Bo08sQMeCw2+r4LIP8f3sq1/x5I4eHlAEFsYK5pAfKQHeCA1An
Es78Y43/kp3VRkVxNGIhmb9mJHXJWGky+curIVFBcJzUVZzNQh1Hx2WVyxrum6rV
dp1FQi8k/c80kebeQUFYqsv4drAyuitg2oO3GtvEiWnGjnUioWxV9J3srXP9DRbw
eMS/8VWOA1oWsM8f5r4swoSXkd+etEz9Np+UVKCUPr1rhA5bwgfjzFWTJO/graGa
YpLLiZpDRtJxrKAsvi7n3LJFnC2tN57TC8MoweyZ3l6mviL9tNuaf03qR9PgLWMm
zW91uO6iuawEUeQgiBipTgB8ybnDzwqu/v5YIPV8RgwWlor59XcdVoOAVer/BbGd
Jp1b+mWh04z4Zyum1IBVNpSnPS3/Q2NxJtFZrTJQmXqxj7B1jfeSD6uugPVQHAlw
dIq0eH5vRO98qGIer7uPTh4lOUVovlBk4gypq17hpQ2zpc/APo6ik6KmOkYpiDq2
2WxMxM9akBZjAaoTrBA1Vx4PcPK3XSCJEVwq1dNB2tdaHxE+3foOW8QpOLReHypA
3yULyHm0lIfQP89KvSpQx3loGnBszZHXthhcIn5V8VRHL8eoL3xaqvH+ATh4HT9t
XrcvAQMLXIvumYL2i5QJg+P5xHVAAuUnrtbJseflbd+pIGXALgJykE6M42XFqDrE
oNOzFGrzlsBJLKpL31VIMqHohMguhUCumiNsLQ7siiFIUznHwCLsPm3wJCuFFskC
5M4HKMZ9I+hK0SGdoeR8FEtfXfoBHO27zg4O6GXQgrrbfeUMdbs1fHrbgkLzycA0
iXyfMCGVaJgvvzbRYBTmarz5nA+UtJGY13Ef/4wh2P9/PHf68N0wruDh0FNJMbeW
pomtqRr9L16vyxyD4j/Ehr/qHeahQRDhfvdeem7R6/1ukBR5A+Li43RP20CTx/+Z
Nosu3cUH20Tdd7Yu3zUtWOZVfkPQwndZ2Gf1XR6f80D0yk+Oqu0o0tLgjysvhGlQ
6L0Y2ubTtgwfyKdRkZ+kwc71zcmx1kjUi1n1yV5dTHZ/lU0YKFsdOSDneUQfcqcN
ycAOg+9l7EdSZPVHGFML7JRLtWx1/KtH26GhLqupw0HmcboFbnH3hgft+e2Zqsmd
balpGyzjwYxXJxGMXRY62VIbMCja23tRa04YtQzSbmqWGZ6W1rSvdePOgGKfo0T4
GAN/GL8twc5T8LwWegONc3R2ST9Aj+z8C25louhR5fpDv/Ri7zQuPg8bLR7CzCSL
q+QLWI3XLHUAals6/6trE2zeEF3cMXFSpUViVJuNKaLxa/5/7cZHAZiH75/On0Fj
rRWX1bqUPb41RA0NERnTbVqbGKwczGHx0vEcKvkZF6kMyJ1dRaCAe+kT8nUWIBKw
SoOHk83zcO5fMJscQYGfurzj7P6XP7rGdXEDrFudLIqOn6H7CebNCS4K0Si973nf
pCTFR+6toU70Y5vjVJGfc/a6qIbKWCOTxBbH1QqZBzPD8kvVK2xtwZ87pPcZ4v0w
DyPn1aCN0pHj4WoIOhkfQwHi8n++BQ7PW6KhagiagEikkc8+42+BwIv85tebSCCl
J1oEFm9TFobtlM3RMfTcun63G3Ycn72VUZtyjbfVPrCAfrOvio2dPFFItPXZzAgf
vxK+cdcAXZzFDae38gZIkvE2QvjOrYapbbEaGvwNU2quUVUWeU22L8b6ShnISSqK
OPHT5vNRcZDKBsscUPrzBv531S/DybWdeFgIr8Sa59kocU4nj5ncZc+MPRu9J/2D
WFoj86zxGEhavZz3uV5P6YrQ9Xs0K4qH9DDc8rO/peei+wFAjGxDd6LKlGArJLOU
WCpp8TnYA+NIK3v4bLb5fDH0drx24Zxwvjk3SU2kPFVj6jpFhZYaqds/9O8lbh8Q
LkVnjVCXyvVEdhSeePtcCc1PY4ONAmMpy91NAPjYJ3QpxFXiQh5dc23bZUKYd10G
j3Nztji8t5BsmVUlYs2py+RSTtRVtJbZ09NsJTeKlZTFaNFqVGGcUyRLnRkTwUiH
uA10LwIa5sWFFf4E0MMkOax+pfKAN2OTeBQl3uL8lZxAfXktZpiBTNILR/8ecBcv
NbzGrymbyzFuonZS4CmrttN5ZbIWn89x81GjwzQ5Gs/IIg/n4r4jI6dsMLFLokZN
xpP7j2d7RD9CoaXp/llnt8H2xM7bmuFjWWRX7bTZKEjJ9Hyy3YtQ8Ylj+wfaqdFM
IO1ojf4nvYeBq1FUcehhwffVlHUM17UC7ESDMcIucBeMzTSDHvcU7h0GpashJ0Cm
KT4+D+cahSVg+ZYJhjevZnlO0R4I6tUjaWFDnmtXzLwyubCJyygUi/2Sd83g0O+I
dhsJLiMS32xQlqK55K1e0nfMslM2lzUwsmz3kVyDTVECGqEPyxPKzBIfDEe2lN1z
R6xgO50NVmIOQhDvv9i3yAsTViolLwJIFu6sRa7zshaa//+6+OaGTYabt49+vLtX
N3MXuFOlrHefCVTzi1d1ZYWdl9klAjbsdYweWFxzek/nr88HG7T8Gu6cSFiI1Dk/
u6sr9dYevUbhiRv4+WXoZhrw/7w31FTFMUmbnKM5EyemOONW74cJKTcncViNXtAl
7D+rQICXmET2czTIK4P5BegPXq6M3t98iqIoXRtwr++sApzXZNaK39R4O5OrHjfQ
S9JY7H10OfepvGzFGLIyJKzoc3LJ/RCxqA/I4syhJ38GBMbvmEVFI7h7c6XSKxQN
J9hIUmN+6xXGI+eAA+0XQ+emYI2ybZQhrIgPWfLxNyBPCy1oMDOJhk9DGH09/iV4
wkSHL0+4YLM1kdnppZYyNfGwGthZFHuP+4Ksx2FNvl7wsfT/UEHjmjwVPX4nwUlD
3MPme7rWkehjUEwy1lYj6vZigccAN+DoE/Ai83awCL1wYyM1WedEs98qZ8WChgm4
AOcCmzHUiFEvPFjuhtbqCU2zqDp2vJXG3nZZVE37iIFCAgPApFnn//5XGpAa5LFS
02xS2xaAykzK4frIU3CZcu+aNn+QzdlW0XJykJlyyZBHnIqJAM+zfbYT1evUPh8r
Vs3N92rR4Vkj2V4ijXgm4sG7tW6Cp4ryD11FSUfkCm+mMxMje5wGkVaDMersBQ55
TIxXrpjC+V3wZJoVwqzIhpvfiLMCNDneCDWLcNRvIEOHCK4ftO/RLCwsM8irVUlO
UuvyxK9S/NsPvmvmrHfMxgY2s7pOup0RH2nbbp9Qyu/O9OhQRJgEr6vIeAOUgm7V
liMpMVC/5hsru0W+5yw39g0rrvcbRXWIeks7xx7nCk5I7XpqnQF39F1I9qFx6Jym
Qf5SgIFYpIwTL4PgvDbKKuXWBBf1sKCHmqmlsaObqkZGCywYpTm/cncKvfxL9vuZ
9dYWnVCRR+T9BuVpDPm8VEeMgyOwODVL9oULFg4iAcp7kG88mq+Dnr8YpE+hqML0
8unldIQEsqPAPU6dNVJU75KxfhfF3p6WNHu+nUA2gcaSHnCWE4jJOGTI6w2OBjSM
m/ydbqprcqcQVmxUAJWkwlU5YvlRGXhj/Qr6Gzhn+uB6Al53B7dVGa9w6fqZ7PED
3PvKHhCQTPMW0VPhcQ9RMGtavU7Bar3zh4J/WHNUbeqKqFH0xeEXffnUuBsb9Cu+
7YYEz1X0HSgYsJ5HpbK+D52NzlJU+1C6WaKlUzXwU4A7UpQbmTMql/LOSVm+znF5
QZNflpowj1UiB2LFz2TPhVMy+zJXtzyL+DazD4ABJ3jsGRV/DYI7+px7rPJ4VxYn
1BoAqBvsg8EdM78uJ3wd900Vo7/sdhVJhGoziDX4tinpuqXvSS0aV1mfUbV5Epck
EnSQTkBB//GOQ8B4mFGXG2bMNcguZd22uMXYdpgdkS2ESKTlFWjk1h87h7BFFObE
PCmx/QJB/A03xjcXV7TMPKZ2d3utu2X77aElRPvTr3oo/RyfdysvhKgh3g6oFLoX
ccV/qyhATwoUBnwJ+2JvyqIE3mQYzqqBhJeshGjAoIxGhiS2DNpkBsY2PwhspDBj
zpscDK9M92I02JTYDu0cwiwfj1Hs6oyw0qgCNuknCfxgEeRterl2tWgmRERYo8Sv
O1sDG/zuSwTQUc/E6/06SI3ghKSX0f/C+h3HH/JGRjueJJx8LKuWbLbJD9ZBeEkC
1jj3Nk3940Fr0YGUaEms5t6RAtmyP72hX4SkXmAlh8rC2I3Zgxxbmk9ffJNuPMIs
Fya33JWebJCjCZ7XqsFxOfuzyUzbsGnyYtZpoYmsNjtzRqBKjE7m/ijmLo3WIPDY
aKQ2QAyJSDjip6VXw+vqEw5goPG7GaYia/GcHnETx/KDPWXQnGKIEXLYvthrGutf
RjtZNPxKIi/6GV6y9r1+vmwm0RuOPIkDAOCpFv87nFzjgQM9nXnZfcYG5nIa/J+H
P09s/fIxUAG0ZAzdiAxoNMQz+edhV3ynbLbUyNTOHUqlFID41k8LHqvMeyJlZi4z
R2mhPBRltzDRr3xRpzCLINzut4I60oVBLjaaMJKO2v+Whc9u1fOS4ZkNWL8TkxsB
RB90FrCzXtScCI9fp/T6ovwmJ5TnEjk3ERDHu+rB/eVySnbYBBObO8oHjAwBSD/Q
Vay28SPDKCZVE7E97ygKhD9BJ0OjSGXHReECJKi8/0s/m51Yt0rAp58co6fKQPbP
Q0OIdXq7nDa0UElyIqV1lJnRNqn8azjT1Af5kBtvAWisG4HnfmqILGF4myeHhPin
l20onbrKUgZBIGjLNqorLUTwdV77PMt8xnZbJwMvoJTcRaI8rhyHX7phuHdlEMt/
CdpogaGLvBqklrtcEA83VkRrdBqQwqtiUVEIeCpBOkOlVy5uK1L/Uo4kZj5it7ec
rWCe8Dc98LXuJU5QBbtcRfUEyL3n8uRQm4quqSqvSvQrAJ5skpP7MWNX3ELTo5aw
yWq0wcnvTeB9tRx6xC7SA0nYfBVH+KJsbuIJOXgR9L9SC3Io46o5z0Mivc4t6hkW
W/lAQO4Mt0ogojuUzCYwGle4ZnwfOweAs3AGgtbjEvYGlhtTSNQ3FoXEjHQtpmld
CxFcBAPd6JltiO+6655io4x7FBGw7GSAUrnPpiFFAUH6s2n9ISGecJkiWA+kHr2y
2DZjmnjXl8+cVNHxqEnGs41fBG0PKqeTczu/aG/Pr9X2B9xCwRalIraFotg4LWV9
IHNAnGnUoH+hMBGCrdk8+d2JNzcSEnpjIGwRjwVHgbGrqDQMJuOq//4ZwUGeRm6S
L83wIWdiTYJVzgx4gHAIehGUaHTPmTOqbPtZjTaZyeCLVbOLz7/ygdz9oFVhgnwQ
MOCBo+QlKh/zlNrONG8E/TPkmahxSRHN+rk6DodxPa3yM1xU1B4M50glxaunGzkM
+GQnSZyKPC20T9sys0YMVHyZjTO+gDjOtqBAleD/Ur9a4cNRzfLZyFD7r5BLv1mm
BFPPskPAgG7Hq0vOJz0mbRf7mr1Rc5bBjCngjuph5g0ARK5/huqnI1KnmxAcbvJ4
Vnt31S29zuF8YJFYn8IKWZReQLrWDJmZJuU9ttTwmKZzjnBCVwsyeOvX+b3RRLak
+HnUSN7H88lWtUl7TO7cx5Cz3/aL5WjFgVxRHarEisMDxTzBKv/gks094N1uhf5v
qPJhJT/z4iY9bAJHOfbdcQMCxksS1XgKvAgxds6y3FYWtD8FY8Gdkc5N+QM3ulFl
uMhisgAg71Sw5x1Wx3fmeiDwfgpi9tsZkT1vhiNUW74DNbB5ylGzqCLi6mSBRYIU
RYRjXAguBSAxctOateyjzD3si9Y8Ayt2nyeEsTI9vsYIEHxEJETNcP440B55eCgb
MS7E2dQpSqbR0CI+OzcpuNUeJ+jOtG02aFyGzmLI+84tmssAAcxBGWdN9Y+nGrON
aqiV3yWpMMLpTLoqdvnaElM0L65lajF2Ba+yd0FaJLKj0WSuRr0OA9t8zk9rWBf+
uuQHdbwep/+hmcSZQiKL38I9pWesUNwffPgZ05c5pEGUoDRTysEtKdc5vj7L2xni
V0A69S/jGH/uoY1et87Qs2HQJF/wOFF2mML0bXthiWYB9fLNfh7uejvTUqkQKmxs
95dvhnQHmiZibDE75k/W+p25dxA6FcfsmZid2CtbV+BOoTbzMa0YhsDJTc2E+cd5
sRJgrgHI7hcDJKfvbrpDtjhLfn3w2/EuleIxY4EajcSlT/PaBGstbA5je16dtcRa
pBnG0SqsY7bJrgvwc/3fxyncM3jTqWC+GL0MLREI9L7DeIlAI493k6UBLsSeAn9w
7GXzKHlK/rBAVGbOUU988HkdBJrxjapr4Ctc7olnwSqgf+q5wfrAjFHIt6VO2Eg2
ZXMqEyD2mjgT6wTZ5Y5FKaPaRIMwKjMqU8OVefpOUbwzeGpg0rGnE7mmwanF9f46
bPJukFyJJBwj7BybXkiQDp3MvuiUwkmTssEP1wBZFDL81yQhDPgDfE4Oya+3nfFB
942k0NysAXxgUt3WwNPDllqGriJvBfSJUVV2+tW2pWzgOYsUvAZPyM9jOCrNWXkl
zO0IC231zmzDmFFFTc9o4WqjCA7r0UGKQYzhDleOZ/H1JTwbEPy+rgxvDFKO8/Mf
p44RZncPN5Et5ds3m/A2niHPup1FcwzR6SqL+QS++m5ghJKRTZhZHEBxg9AkV2ds
BqRauu3Ss7QOfFCPOhATkmNishKgKAcyhaxKjpPEIDeZd4KtbxbhS9YdvLQjCFSE
VhCqDcqmhsu85JqWNLceXO/1EKgPeGjron9OKxI0n2c0HJ+U09neQF62uXZXTM1r
3huppdF7YmxRZ5FDo+x8NfkxPrIKxcggUGZs1ER/4st8J4MYZB7deTAaw+Ox9pAY
7541S6CPN4voQ18zyPT3V61y+bQ9a8np42yIRiLgoQ85kP6PO2uNjjTCQjdN2G2M
DRyz763KuQChbhbU18prTPSjKZXMOQkay8n6YbfsBhwtBf7k0z9+TRk4CQkU1DCo
mvzTZXp0rzYFqyspIkC51WPUBir3vHoiXelckwh0KzwZXDVICQbixoib5SszsGVP
I+gvec0k3WqKA3IWHx+X6Ci5IvUckDlrrggZ3g4S4Dp8elUf90H46W5uay+cuyfA
gPyAXZpcqF10LdyGTSA2T0oiLB1cCOSyJ8Brj2sM/gsxBh8PBm0lTzIRbQ77IAHu
4MfTZQwIDgOqKYUIFJkQX1CPzDH2VDHwBUtqg2kx8SmcGSHKTdiyCrN10AHq51Sa
34lz/MkOhjhprs5TlEeBkrjnqAYWxGkJO+iPwCGexnyltqAsmHwrm5gOEJkzyR0o
TS11lJWOb4z8LYhIpbCbfNMh2HqYuf/OYSzGHyTmmL2K1EnBt0Pt1xyLWZSLRDO1
jbMU5JGgOlt9Wiv4qw0KdJoHWglaw/Km9pbju6XambT9PUzHJewEGPFuwRv8Z43u
gF20tAq9DGW3uhg8DHLv/5FG503pqK6DvV1OO/uJNz9uVY+cUutf9Eb35t8mvhfA
wWe+CbLwCBSqPcLL+nprAEnNG9BgGxMXdxyNgx6dPvurE4CcN3KxFcxuvv6CPsqV
VCk9et8gx4UOqyMrhk7y31ZNBfoQsn/8oWsIdr01jCjnr3wRhvD8hvm2bq7FoJoi
+zaap1QaL3zTqPYAcZHnna/abFQtUhRmgDZDkA7pGaBhzkQW2W1rsPuQ1hs+GbDx
Ue4rWkklq4ovCyClu8ElU3CypaoLoA90j0ANn+sSPxp202SEDEkD93SXefWuYMCt
34CkFtujLE7FZ/uFfUZaPyqSde7EHfXlLGNMniz9il/AnITnMUAJE4/vvcHHzwz1
xX4ked2Fw19qoDIiCvuzOFqA1s9mm1gl+b2SK/f29nHlG/zTblE87u71PrCNKVGk
m2MFi0tNLhn3238pfPzuCSiRNFpJGnRJG4DOOQTXVVeQoyPUCBTp8Fr0qMcpHLDR
fhJOcArzAJ5M1IdEjIiVAZVQ1p13j0IQIanpyxp81lxJtWISIEk7ZzJ5STssYQCz
BiYgemuT4ZCvXzKnfI+FU6OCahNXLk0xQQnPhU69/TsOq8G0kjqBvLsW9Fsj7IUV
MJ1PY+AuRRC5x4Euf5XFyQ4sLXmP6okhocQBPsJg30UbYFfoE/LerZoG1EX1N5sp
s7VRSx/eGOtVAOEN5okeUMJmfHJYucyzKsfiQRTBrDAV4MdpFt5+SOQynGzfspdL
tTuyuNjF5TYWKoIkaEvD51kS7KsXPpdFBL6Ifjuj3f0vaFhLcXXeMqoTR7S0cP0M
4FOkDakYCBcqFCHdSj8bhY5y4ITI0xePddu2W9RxDt7Mz/r1S1jo5y4PU5VjaDLV
QB1DxCsPUlcwXHy5rhUmB4cuKV2RBpEKVjhc83WbFuQSCv9Ne5badfwdPfeBgW7G
0RCOR1LztsfjmctZqUJ+kb39ec/Y5uHTkKOntIyjztq/ZbRlHC1ul9X/9w/c0yfg
3ILQS7gDiEOJ4eiiyK7kwzYrPTX8+bir4oyehkQV/YHLtT1e28Abnxt38OuNWL5N
aE6DbQIxkMPO2g+B6N2uDaL8l922VID1pyIpPLt1DlGGzONDaFreJ72PT2CxKGpn
LcD5PFa46XCF8eU1SPEP/xK2+x1VftYO7ExbX4jRTc8zGIRZlFOxswG9VjrdYP4A
ZgeG5SPbhnkN4+HjX6MxL0trDE/uCmio2yrt2f7frJBH8mf7HcqNeZOG0P9qjcLL
pkAPqmnf7G35O6p7GokEesNRYjn5GZP4E6BfCyNOmfpgHdvDDFTSvHqfPNJJAh6C
Q6b6xBxOud3TmGDxUIOJot+xC/sbTA3mM77OguszxAF/3W5qoRdigTdrRBy7bRjg
HdTdqBnYqAke/oEzHxGplSy6sXj8jM2DBkPEZQDCdi27/uUhi/30ql9xQY3+oobb
N9RuevxZ9fPjHY00tOcYRewFhIHghQ0dptQ0iXxE//mhYB/8TiBTasVAkU9vVxzm
0zkSxlPKGVX1r9YfMTYbbZjUUk6r07l1lIa3nG6DZFCrHXD6fO0FoUCMXagtGaVs
d2nDhaDoNsKKCBxHkjaQj6P8NeI2M8atJPMt+oYK7AYUM4sBTpul69ZG8FrsuOpF
vLqt/e4CFVT9/Ao6lryI7wa2JZumh8gmNiIsWAu/zidQuFJZPSQytC+BGVS0NsT/
yLLbtG2kBM2yeKinaw/op8cIsAa4iSI/yLxLmiXeACIOaIJ4TBx8MD2ql2R/2aX0
pag6NhyxXlgEjqOKct+7Ry9Jq07R4vLFDME5MRV8Q6Zt0kJhdv4qblrQoN44EYeV
hDgss4ZqmpklafJ/BL4Tc8HX9GRW09UqoOHw3zHJKu4ghii5fxuan6uSsmm+EK/X
m/8Cl1/tMIuI+45BFhvYQrMMtETw8jvxvZvXdNfpUp0Xvp9COVfyZnIcEIUG+ae/
rsw/1DLfQGVSCZcu770Q6TiKdqUrEENNrAYk/3jmH3UDOJ1ccAqqGigbiklOkct7
oeR9Mp+W51mFach1G8JC/m2gzIL4MOKToNN5216YWqUGFseSsd5uTBBe9UxIol0M
vzAGMJ7mbHINFlZTl/6VVIxG0+4l99RVyyXItBpKfaWE1Rp36Qs+gh66faXkpTwK
GPylVa2ACGdqfnn55v526rcgzQr1ygSomN7Zp97JfKn/J8y8nk5YJLn7exMJjYiY
09EM9siYR61r956lFhPRYmFiOOpT4v6odjyzw8jWB+kMmcgkOsaMj/M89RGqILwt
Hk0CsVveRkrTQPu4Lnn9wlIbzg1sLXMPWUR29Ik6d7y1oW847xG2kC8aBpzU7zay
gmBDOzO2jqpT+afHy8gr5nUnKMcbroT3GhqcN5QS+ZMN6mEvWQsyDEzAXbQe5JjL
A6+2254/XRP5qf/KHbJtezxLg5PZi0VkGSCT+2fwg9XdJSxvy0Ek7cAwns9cNR9i
GUzChmQFjZKM0enNoVEA5peoiVzy+k4FxRZcz60OI3fr7Iyfp9hq4Wp+vh3m3uwX
i+3x37F0XzxamhBGS6u8PPwUd32lgLyz6IOpUDQNaUq8y8dDD4n5mpIFaSteRK82
ZYA1jvl2Ai9GXwe0UPq9zY/xSl8c3vKs4AAngF0XUxRQhQhC16SAtEFbYl977uQI
IacHhr/ElGSKb59ICpJOzUl8IA/XhBcRV3wI2DX8XMvX6p4NlUEPNjJGndkgSqgp
78xDjJQ0k/0hoVvnljbiNLywEIxkHZrXfcccV2YCk5vp3DiP6M+jLs3JOxTL5yzR
xlZbukgseq944ujNi6l4BMhsj2rfvJcQT5WqNHYvoq5UaIPd0xl6EIZAUC6WiD88
s2HOLAgcyTDRvEzLjYynG2My/mK8jCIlGBFimng4MqdhquaFefbBHokmaEiXfMN0
ENE9MIqlauYLbke9gDCuo8eWYcWPaWwsu4bfckNNPZ8s5OC3x7RpqkWVW/Bliv4c
2YSDIsgIEPFY1bawT1jVIxwQRt4xSh2PTykX7UvV5OHWJQlTyaI2M9oDwUZstGkE
EQF6r2KyReQETCcf0RwVFgxbnqMffTA+BMSJ6jhmaCI3bkSO/avIZYoT1AD4cAFY
IMuY6UN7Z1tUszAEzv2OIszvc1S4ePsmwGtSJnjJyibTPW2fXRM+g0IKEIovzTAN
6E+Josu3A3LETNvEwUfK0upQwRpq0D3g3n4P6ENqfsl2u8NP5Avwi0grVJFqMXk3
iATQB5GRfxpniDMYTbzpOF/vjBb9fQdN43NBUYZdsRMzg6o+JWkWENN61e9mBLXh
Gz4SUkxw/HyKvp2PP49cFBbF1H6k5xwSvQLrrmewuj+4s0CGhwCxSsIb46wcMYL7
UILqNlzOyKNExZQisDgt+XqFiKeQbx36R4WEWSTyqsfzmlK+BCnJuiFGg8YwutUU
1fK/oz1PO0GVIClWPdrnXFhFtY62JA3Y3UX4/DDRSdjw/7XD0BKinuORtaQCdhOf
OfWsytFPmxz/abTF4LR6Y6g5ecBfW1GFxBUVlLiSfNLkhlcr/Yf0lRX22pyEV3a5
6D2rku6RHCC3EFFaUGCAlgg8r7uLDI5BKlhW3X5JVxCDW3/51VPOcgENAhhxhup1
e2zcYdUSno01i67ZiJEam43D/TFN92QUdgvrAmcrHW2lGzZq0/0AyqW7SSJVhipw
MWjOUW/dhv1dxbSjA6zJ3XC8d3Q1GfWr+orK0QMePnUawsByQbBHAAEnh8HdN+3R
9aZ7qG2qHb7tFFgO7TABEr7rGIZmihIUL6xrYG8u9dqBLUkZqR4ysJ8CKBvHzUiZ
w4TKx1VmetGP29vbubYjQxunfazxegBuZ0n9oKjPSQBdhMWSdc1LfhIM71tqoPhc
bhMsDLfKQTL6RJU/j2oM91Hh2Bo+U06WDTkhigcTqnxOVryis5+Kkdh9tANe+aS0
tETQGmjfd8arjBmElYwa7VcYasyq2nxVBQc4XQQbQbayBgJWzHKnjvomMx5DE/qT
L6VF2kEu6ui5yXbS+p9OpT0mjI0tCqnascnHF/kd0hTXnzbjVwyBqow9AjkCH5wz
vNce1FYL7ESoYqvcXN9wVhO1nahqpkUwUL5VV0vAYx25X3zbeW1Clj6GxxTpla25
jF5o3Pfb1J3+92GMFSrL9KOft1Sty27RnK0OthbChss6OYZhTLZzjWD3ET4mT9AC
uIj1P/k2Ztx2w0afvC8SDh0JHP1qz9V6VQLrPSOaEXlp8kda+2DfPNtzC5oOvKa6
KT/RQqGsAfGgMCBXiZfkQ7epVJBjaikALv+drBjRQP06R0waVZ3g6777Mg/1Yq1p
iaxnnyD5yB3HG6uUkO/Tik9PPYFO2mkEzh7gEwDCPLhMb66AM461nyyIUQ9dx/ka
VSX3qsRORYD2QIZQulICHE2RCSSXjDqlhRjhW693vTR+DURkBR+255xXYf5qK0VL
4oNhux/FscCR0gnnK89eLdseVSjb9HXugC1VAC7ilZjIcU5jrqjS+/iYgJqnK6Lk
UueC7BI2fWU5tO8B8LfTaZjg41qQOeym6WmmSZ/DoqLqooeJosyny9qC5neI+sAs
rJUs4vZgSFyyK5H0qhBcMWHfbWVwGRzzSQ0Ou4qYj3fWF4N1FPRa6DddzlSJHm60
519bIVSQU8o/fooVlIJehik/PqktvshF9+YporuItF9GU4uCzDp9JDcV2QRxiurP
AtBl7TiR6uQjqQBAqncRMutaWpn7HLW6dxXlsX3YMoQkQjY/1lfl9U3GCkfUI1TE
P7ihul6bcs04Hlsa1d6YYSPCqfFBEp+LveENnEtknwXybwZIAiAeP+AgcpiHXnZx
AHpFraolX6KuP3h9ZvxhB1ISbdlYRiz7XqOBgb5dEWrk8TwCsKAr+G5Zc9ZIU/Lj
72+Ar12GdCrE5yMpmO9k9wsmqWFVhbzRXvRUTViACaE7sEHVd/U9I2QMWerIa89e
bEA5ZmXyIvZ00Oan124/1IM9Fm4PVc9sW3ilVbyhx92vq6cuWgCh2jQDFRF6z0Dw
NzMDL2NWDJ3Env69zteTGYZASUm983hL70+Ya1ZhQCxoY2mKAWw8atyBFxS2gGIx
UU/tBwRh3AIxLxzpD3kUq1RFCthWUtKAFuqP/CXoSqVvcnw9TCyio/awvCWkmtSf
QctQhZilKC54oKli3oDfC8q3ndBYhLZZI7JfGXim6/jGWL3RUqkYDgjff1XsnKaW
jAR39jYobHIO0Uo5gh9FfT3Td/DGAs3BI8ifQwoXKUB3jvcuc0wBYjbaGXDF4qu+
Z4Pv46ZNMwJDz3yYEEdokHdrFT1VdYqO/CnYL96gUO2rO14GkTKnXfBKg6yTdE9D
Jdfq43xO83A4tRx6t9eOiG4o82mxaYv3LbjJhGBly81jdVWnxEkB3ndkAv/h+lFF
WK8QH4wAXGMy/A3Cw27Ckj8ncXCvanPAzurA0OcG9PRXnkiXx442vf7uz4bd6iZ4
qM5UZJ+jpPoYACXoxUqGUL6L/3HF5hJCtYPAvXwPX7iIqIBmqfnN70f0S5Iel2Ii
M/4SpC6fOyc9COMrahhy1Y1MXBMdWWkA1lRUouhYm/D9t7rZk4IxtudhoigqCmnn
Tw5OjRZNWqdQUnuXvB51KeCKG1p4PBuGsWw48tF8d96qiligyTELieIb3cnEjquP
kBDi7T5Vctpp4UCx8vQEoK3IfGssUlgiUJWLyUQA07w0GJheZ3dSMXDBGSk9nULp
rvEFuPLsfhiJtB3u/+UGilz0aIOzHDwmV3+38t/xcMicrFEzsjwAle7wP+abfB6w
GqPTdZhZn1PPtuRl4+2Bh5m1yT+k3gPD69xkZDI5FWOmHINRS01Mub5TQi2/G9rn
L7kJ9llZavgAfd/FFTRt0Lba4oEHS/x7NJMrTttChO9/nVsRvmA2e36PZZJEQTjo
5D42f++xErIHmgKPr3NfAThmocFhuT+kH67FcJXDl6TxbTbZTwNUjRn99brdnbG0
DC4xBs0FjOEicq1a1O0oqJUYSkluNL6GY/my0wFL0CI3RpN4Wv7F7qt5lG5ceDFH
ga98KilY0VnulvFq01KisTvUX3UQrfM0utrbZn6iXRYy7817/Lw96weFwWNL3ux4
YNxj9UGB+Qp1Do4aWwRoj0QoRE4WienxqYpIP7Acfc0yA+fpKkCHPF4tiWO0C195
XARNZ0pcFyA4N9cqTe1A1oHndxhsLsRlET8zN0BnyDOurZSxfcfLvffxeIPD/Gj5
JJEPyVaQUAKEDMAHAHB1zL1KdMsvQWIX8K+R+YRhbFMVc+yPtg4YUKjqRaMhJJNF
WOradIVHrqTu/ACqFY1pUEu8+mZlLW/ku2x6yM9TTahV89ox/QcMP1tijMWVLC6K
NZD4Z3n6AmyxJP6uYV+PEzU4+HrPj8/z06ePJpVMZFtquIXu9HFGYbuFInekktnZ
BCUWmoQcmbJPA1tExOG3fGqLBaL9/EHQ6my4xLwRiALdTsGQX37j12pYz+txSILb
boWYfh9GWoZMuTVRrkVvFcNHkOZ5Lw7wK3VuQ9jP3589Tru3AXsXSWgRxVxK4Zlr
X8hh1wqiyQaPwtCTvVAv41BefsJw4aMpMtLM1hIg3HTZpClHtXDjiJJ3QIzYs4F/
qqMSpjgPp/kQl6K7W3SHp32Is2LA3BKWQ5Zkwu08oikKHehiV69Zy7gT6/OtyFiM
grvCAf+i/4iKVDYdHk4OhCAFVR1EF7W+g09vue+xgnKBQUuDutftSxSSaY2rvx/p
mjnvXKVfdyuZIHOOQLnyKN2nfaCeYusCVZUvmQKQ10ISLaRWy4WCedIiIml2Ycda
tK6oe4IPHDcRyup+wLHH0BvKErgHQbMRo7sEPxHq8IYshCS6AVuR8uZXXzAfeCaf
0Gn6qseyeZHJR92zSdTiiyuUHf9M4huVqYCzr8WmOgtwJkLYM6f58TYnnvCQhHJY
rELbS/d3n6OflRgq1ybsiMmGfUMHFZMzw9pwtsLiH4Tgf+NvKtcBQc+0xiy8Pj+b
pphjYONP7WUDNWNi5+gdVITfYRqVgGf4uyU3QhmObiZ22HIEcKZRYEAjeGOzzIYr
c57i7P15QWUe1G303eUrITAhnwYIDcOpJez5n5pLDT2hRr3aRYko/RZX/bptfdov
JplIqgTi01MmcP7tLNC4rGzbjLQFMFufBRW+tqGX9q9KUl+wQwxpDe8e+EJF3QdN
zGtNDtt3g61cJ5WqqNi/MPZ9BDP7YZGctSx1YGMwF6zUwCuf550UIRa0VB1JbT4o
mnD59KJgQdaK8VulMeOREbpXTUCT2lLB9Fj8isDacFeno7qJTpLBcx3tXwr9ZqcQ
ZEpYSn2Xf6IgmUxtUdDazaVcPzWcS5Pv3YXQY2vtEPUVsyRz0WXcx5IMCrLoZKR/
hgGjqyyTpXfubRU1vgdxE9PBBBEyhg/9nw3sF0mzsgA/Kjcd0C6Y+i1MFXSElhRb
57ZDIT7ZHQQ6039ew6aEPC0Q4UVy6l2pLICuU65cFBz5G6vdcb/v61HrOMkikD5M
F9nxoFEbqb77DbBvGt6s0XT2b6K3MVf7VKJvLzM5kf/HgBq7XBgYCwaDnykhgvZL
sqUvmWkCwYcYpYZu5rk2kw9jVPkUOyoyuJFsbphD1I2U+CB4c4O0Qr1g7o4BCzWi
28CTPEr8zNZC3mxErN+CVaZ+bBhpEeLORz0SIlMwRUrdYc+5qs+KsPX8dxGeeTpv
QmGzi/6iieNfp+GhSAqgxpyDb1Kc9afSFz4zJKQngO2vxzvHCkyNRNHBwuF1Iucy
8gYELtSrTgkmAagTm53zBYKCTYNrAjLiOKx2atq8NjKtkvFOxCBHrqn2Qu+incj1
MCqkrQF1WktitplSTAQB5qkMozPrMpUXUZD6/QPeED4T4qwsPzDMLakW0uZB5zfP
xH5/6PNAH+KwcAbSFgo4HAcQwka4TV4aW8xk0v/44VmMjxBKcySN7oRSwkPWDsW7
0lT3KYS+oHEPW/7+QebQ4KLieruSf8JQ2WqHrKR99HbOKZFcTu7+b3e06WFt6Lyn
c2akO0zhy3UgOezioNemtxB9FAJBYwwwdgJi4Uht3QWNrK/9jyoGL6hk7h1O8JAI
Wb0WmvXZ3UY+1ENhQVhhi6oOuc1+HYN7RiMEN7BDYuWNuc2xfYOFEJvPhHMvWO5m
evlB3Pp0ET6OSu2lERpxgopn4u4nnt2nYujShtMY9wAwKXLHFCE7FVG8pCu4DwFR
BQQxgLtmnPM8pqKz7wvTwpThucHCzUy1JcK6KmLiP6pacVA+VmGGJhz/lPKIzK64
+5J991HGqEQDxQmuopQFbP/TMqdXXtib93hktBjRsmDSbAsKM/06G9NECgKMCY7a
DdcjCB9lzNgVHnXsgyB632aAB0DmJ+JJlaCW7yMMLsEd5+rlZ9vozUx9HgTdvWVJ
ycdd5afW31Z/j6lpZ9QTzTngShfyRRW9Sv7a3BoTZKWGSeF9iWU0e3+KYGJZbhCE
CLTf0h/idyB+P6pQMgHGor8FfivhstqDpykbM/a1iM6UM6B4GFpw6UeabS3TXl9Y
ArbbMPsWdQhCc4se+85UixTSkwxuE+dTExVx7D1T5QmFOizp2RG1xz64n3fZcD3G
JMTEdQEumm2sxTJw5PmNB5FnIraRvMYfPsSUF7ckxerRADfpUAR2jyVia2aOTRW2
Yk9RERSO4Y1KZLsml1He/0JrnnXmKforx6FSbSsElYYnD0+6V2XjX3X3Xdo6m5NN
E5U9qr+NbopZZWfdtbV0lV7qNKZ/Wxk+CtYkAt6eCV+JI5HERSHjMJzh4/dC7snG
LjKmVBd+r2KwgYAJak7G1ofjrrZ3MJTG7uATRbzABLtRSCRl2Dz2ZHPZNsCiR7dN
Svp94LhMSx1tF+OQk1a/Wv54eRDXAmq50zDzLFZQLlhoKI74R9Q3B/WJ2VTugKmi
pbs8yC6m5GbhblJVyXiNrxmIz7zHVKvJH3djGoNu94g4ysuPhc4vU5mnL6TVGkMt
EnP+Qq3c9KRUj+qPnMPL9ev1M7vLH84FZnZ0/p83i8MB2P4YjaGJg210osb9SCdB
0RATq4FUCy+c5e3IjlO/xI8GG9BCHCOxEbFJicum27L2FajB0EXzD0zSkLfpJOyT
r/3J+ukBBMWlc/1feq6P/k+Y9eP0e7BPWwe5z7oTskISd43wq/AjOuw+0DWtQA7O
z99iQbzGXsdvFoV8SQpHczRzGnY+YC73b9aAQk0GmvUL9Ilc71awf6iOk47bbFWk
t3fV1yQZ4sHqbJJFy3hQ614gKhN4a739jtaWi5Ya5WOmk0dCGFY08rhTI94qBRyl
2qDwS5fjIEG20qt1YJYmO8O51jcWj/IUhSOJ2CK0UZsktrC1uv3cP4W2plLFuOpY
wGRjmpddlanbwHveYJ2JJvyCfckUUL11VvdXkmEFhVWjUkOzgLF1YERMhTg4hDko
m7kvQqJw59HKKXYXi0njFLY+RhbCdgJeeSTJWAqYcw0/3m3Xzj0Dlc3sckDS5/oL
OuYf4Dw2GI/WnuQhBQy0FUSaovzZnh4MS1PsNovMdwJi9NT3PkLiLJ4IhYuHVjkc
GlVQLzR/9L6FYL1ODQI/FiL1ml2hqCQxlzoVhZyIPyqQByc4L5DxZ/mzUpaUQN2g
LWNttInvMFMJY6qjIMe0d12uRiuiV/zr6pGbBtmMnDERkKJWzONGsbmfGsTOKp7O
bxZLG7im62PGS4EIl/DBy0IO6zHG6TWp0eV/NlIqUv4A5Z498BtXI6nS06hP/DoM
bZjTm4pMiZTWBpqYPRS6EJA0gAhRn+AOcfYaWnIWG7dIkNxeQkAPsllaSM+jJGAe
knFopFVKD/EQLsOrqteWX+ZIlDLzx9nUmSGakbflK53rsYHSsV8Nb0vcnmDpz6xU
r41drvlxOReLsaTHBFNyj+Z0Z3nUM4YWzMWums4TQ/hPsxWay6Gn0HIc5sW6vAXo
oBdE/kMr9VKLi1UgG0qgmfartJXHn+e+c39Z145/tihNhnp42akIGdn1IUZZplO1
M/K1LwQnrqNbdctwKsdT4+tjUNtdo8BdnEfimP2hdKy41q5XZFleSW+/uerjH292
YfTHkzRpMuOIXrHDYnDVnVXzgnYgcsME96VwJZOAtb8u6zG9gRV5nb8DMtClhvzM
NGpLmgloa53TJgWnawElEu5aMf8+NxGMHleHW88wmXAVa03gdOVFbsEGHwtpXsZn
KBFuGKs0GSpyO3oUk+YxStAprE/Ur+41ttiRswniDn0KWiooItEL6aHHgXELDN2G
hzL8HBZNMb7WaSjPJxD2z70GRm12eDTTY9web/GQY7S2W7msItKqLFlvPOcnik89
vd06bitZGcADt9mIoiZaKO/SGBQZxeGYUpTe/qebggenjWHQD781mF1OxF533jLf
T2ZxxgsqKqze/gqrX2OdQwA+JcZLxrs8oJy2mGKOjbOxwxLitvCkEBZavfN4xlEv
1AKr5dL0dDGdq6krGoRVu5pklTUGdsixyg6VZyLnSHdd/LJQIXScGteLFhimAGz+
W+X1kIgaooHR1oVSGdPwNwdfNcWFcRLZEHPCe3rAgFt5pAEKiolkTQQhm/AH23fq
OyG7+vjZL6IW+NZygg6a7BglQqhNYv67KfYVmQt181XFYyLIBK06M6hgL+vJ8aQ0
rXexPRTVmiXVX/tiu4ksW8aInpZKWHp8LbhInclEPaRKLMk4N+2vP6so+ScTBIYv
ZMqRopv4Z4H+amPLn8WYK+kPOEOaoEEwWunmslVpXqRxJYKTEL0Kznc8ye4yEOi8
SdhzRS0Q9UeY74OxpeEoi7ekqycM6fseL2hWpp/4kHhbZzNE7Seet+eKjbe61MSv
EL+bEdFixTiwP8JMFJoLEWL0VkfnqyCmGH1vjZLEPyX1Gt2AieZ11Fe1msQARj4L
573oFqiGnCMFdx/KwEu6wku99ozJo8QUlQ0xX1Unzd+LAkOSEzbaY67JM9u+oKdU
zTTQmuVfmc+KQyrxE5RXS9ewrNWcb1hQ3nnOg4F6bI4cLv/lj5EiaXaOUSwIk2YW
2STQAMa1C5l76/NVmgweHsffb565znH7z7L++EiMhnpPaO8xp3VBhPmKRRUZv655
H87sSUmvOONOxWR6C+NtGc75Xq474Px8P6BwRMq6AjhOzSs/qBs62F3LSaGv/7CK
G8tmW1f64SplQob+vLk+v2dyL7f3u6FrMT79a7f1qQsM17JRCzEyEcWnAbzIj0j1
Qab3xEUSPSKYjCw5EtEjDwAzGEwg98Qd8D+B2UiLTP20UrFqSnPogOLEKFZpMYxj
vXj7T7GP2Y62Z4+MDsN4JCgjm7M5vF6F9jn3j7tu+vZH7UKtGxh9iws9SXr799uW
C5ICxc1yLZ9kM/48bFpZfUXFqv0zisLiQbAyK3nXij6IoF6OcW3jNx599KZc7cHq
uDR1eZGOr6asJJyT4pui3bFoxDTM99wS1gr+RkUmAUIZ5+c3z77+D9rg7roKVlpo
ts6df4OqK8PzjlmvK0ZspRiMf/jgW8n2MwAo7YZcCWMdJ9HpU/jhSry3AsUCeGRH
yLgUrlFLNwtvrHaGCiNeC9yEWmh9MM5tsGgBio1s0AwbQHz4EwqjYeC4C1qdZnwG
BEn9WuJZVz7tbYTBcbLa4vdCcOtP3rtUfTWPXcd+hO32bARFXMj6W8wUArVv/xsq
Qm/OUy3EopbHmScBcc1PWadLlxEFC46It1RENJQjSQjaMs9DCduuh6xFB0Qy1Rox
fI7pOg6uOcf3rJFcKSbgOj5FxwGMmm1Mx0hsbF1m5b2Z28gWu5TwVXKmWowCNYQd
oUTHR/xoiaxiIApOChpNY5CiBJUb+iZT+KAMpW7uFnkMhuptWlnQRVDQusbXymn6
VIy//0jdT6tAZOwQ8NuYX6qqRXUu/6rY7yLouiOgAycuUn7+oRJsuEhIFjDnbIil
XhHJ/js1syIg5SfRy9jneeS5RvTcoLrU8HIln0yhu+Ihy3y/OeMcRQykjjbg5WjE
6lgkCT46Dv+sJDweIVEuUBNsnEGfl/KS01Ahh1YYJ+59TntvGMSqdiXCGW8R+UtL
aH6NQuy+kXgpVjEReaNPsvdWgRzz9FI21LjLf5ShBa0t8Q5NfVBIwLVzuLLH/AVo
IVxGpP+I8bzhTDMNwmy0SOnYxWLbmBAbhzyWw54O2gnaoP/6IsOplccwu1HR3Iyf
wuu3bnpegMGU+tqxSBYeOJ2XGsYbh7GrBK4lSKXY5L3S2+zPyZnOeWmSohSbcyjO
I04mkzgoeamWex6CWVZhBhw5C5Ma614UFyFUtHp2l8edikz1hvJ3TyrnwFiEvpJK
BP6ryPJGhx/y9XuUJu5SxHmgiiXbI+KeqS39KmMbugTDfV++HZxJEgaUhJ0jzUfo
5ROWxP4xsBh30F7dTTAeedJceeRMwtKICOPOdOvXsHauJjo1It7Z1+nhWmqGDD/w
O9oAU59Q/IFHCs4q9S2sN3LYkz7qWm+YaWA7pAxc7XEi4fwALZXQ8CLM3nysPtO1
3iULb4IjAQ1/1VQ0t7qlXhMcnOVOLvs5DxI2PztrOJ6o/JGzYsMid2dGdapDZFGI
Gx9a17OiKXNGmlBCqvFpcNILp3GMGZYdBZEk0Y5D9zdlK2EYkNACgg9q3M0s48y+
zgYOB2qXESHmnsrAnU7JBp+IxU2Dv1VetNYFkq5M2P+DTmjRb11SqARWazCn6WUH
Rc21cosJgCxVsNTRBVdt6Gv6kpmzK+pZ8Tlz4VGJ5PbrrQyLfGxOkgpNemvnE+4V
JAZCsoAPdUZ2cT7RoZCCyYB8yg6hJfWYP0+2RqTZ2puCrc2As3ntm8IkMu88Bu3Y
7z6i+vZ4Rfvea4D1k8XpIglfdTY/Hg0fcYF+P5cmZVwTj3eHfF92E5HKDB7rpMYs
wt95WJCNbfXmZAUEbVdqskoTUd/8gg/UvhPqPATmyEdaA6Su6UKU2Z5hRJQMb6D/
oOgdjXBJbXqTsyG2TJ1/hueuYOiwRVWsLsf9pG7Bdtxqmqi8UY7DAkolbEbbEZvT
AiBNpGsjB+tXEjcDX99Q8QTLnsBW+JIqSsJi9zZoxHPB8vTYG84cBESIdYxaQwl4
sUD/8+v7L0UtYg89spUw72uELSGSyushsYkcTAvu6CTxvaq2QWD94HgbYE+UtHHk
arnRlc2+U7HfqaDMyb85rLO51amcuTWwliDgMfN9/T7zki1WA+zSqS+06XyTuAY2
39tcWzppepGg2lbZ6MqLJ+LU4jMfDle3HBxNP0Sv8ry3skkh/Q9YxZ3ia9+LF98a
+O8RQL469zOhIYW6NwMmyatJHw7HBMOinHB8VxRu1NjSEXQ6ieXpoXjoOslAJM6E
orcfGtPI1b1kqdf34IK5W4cWwpThF1XsTvwejnSq1iLpjFJ1TnWIDJTAC/QMcUxP
QsIMc6dhtZWaQ9N5YrXemdqBldPJLZRenupIw/kXog55h0e5W/t+IPVwmaVbNlOG
T3/ctShQQ/yMpXcKsEPJEpUpIl4rbPsCBouUwH7sXpFyCJMVKy8oTCh0UCowU83K
A87p7rulqZNAAnVFKR6rgIh9tpgTmfrOiXgtk+5a04YGxJvV21wnixWL5QgN/Tn3
PNe34XIS7dK8nZe2SlLptJgxioZyGXW7IMf125LmaHoC4uMQ0g1vuH6im/0oqHGc
tAOpEzvdVVgI9sP7KQNP8hPfHh8bblQO8/UYNz1lU6gJrmdbyBNJe3M7PH5T4Mz6
CY1gbTLLtXxrpZ2atbRp9ct8mUZIjsveeCF2xGyevoQGFwi8Ph4c6DgrlQq+zml8
zpOjwEKg1q6eP6Tz3b/G/OHhABnxdRTQuSJDjlLHfrqTnA2tHh41mnn1RTbovK6M
6T7J8f//NNDX18xLqz4whxDT5bwV0FVmKVxJNZCPwcFFFxkDcQ8imKYb3luxdtr6
r5WfyAA2waPKfOM7Hv4ywMPrJar3pP01mH9OrvOjQwuEvofyIUtBdMMB2GBArQTK
IviMNJSQ1AMU5Rw4Tt2phz3tRCw2Z+/4/6EuqPA3AE0tSQEjaHBdo0oE2u0t/t8E
PGb36TD0x40HZqXOAaOjD8PtQLRcnXVSQPWZFFwDfMHlVm87aAKgOc8E4FcbDkez
hC9v1NjrQEgZIAjDp3aE1YdyNd3ECJA7qwvju1gqJzpCultLUgfBONg2MPmfnsrs
2QR5iH67gdwhMFjEzQARAwpoSRc57cCkVG8pqHBt5ox4T0rM8fGpeBPLWpjdwWOa
Dy185m1G4aWEo3b0b75J8bzSfO4ZM7S58hn9sNBEbWS8GYMyZXWNcn8PfC5O4YGc
rDYvC0Q4izeUGzC7ewRHtF8XCSnp6M9oehWwYzgUa8cpkd5NkWHdmohlDKopM6Jy
ymNvqPOw9LwceXFIMLoZjz53ts3JpGiTFcaqG4b+oxsGnzRKGlJa97Pfp81KR1ix
GSY2gWI/xDEoeYJCYalbM0pWJzHshgdOp6EedLPWUhersiCZ1ZkxBvyRvwxfiTtT
kfFn+TPW906yv8kNHxezzm8qbsBfeE6WSVGCjW/WfAOjxBlKPXRi8OoTYEdXn6pQ
jYcxw1DxTE5z8G+NNsEk5G8yX4JvpwJ0yy567cU6/2YTiTdePIp+1Mmff5Dt6wcu
g9cAyOdp0ubInRTcsUuw8heYgawzLr/ClTFiUDVxmseLj7MJ7qSbtNiYqhWzkquC
W7qVeSywdSZM2GQEHldiz5r9sDSLRW86tsUmQlX+C/3lDKazOy4DpaUOmoxm4uxJ
hJyOaJYQutB7DsWNH//uIRP7nakthzxHRYTOik/GzIy34NpZm6ekt+2j7xkM7KjT
CbY0sl9WNxyJA/4W8T/Zg+M4NkcjITtTpOZ69J6CFspxw3Pz8iI/KUycN32U1ajE
BDNI68h3uWwI4CccNmnxLEvrmlFYg27OLpZ9ZEVivJPiX8tCvhbo6mt8+AQrMxqm
ANS/K8KcSOd0cEZuvkKpcbigd85f7mp6LYuiIlNrsh+JAahCXkyZibCHi7dq01qM
9WPf+Qx/+Tz/OIP3wZmiPI8assAy6yGktH+zl9slWj9sQfB2iT7E7gZfOd/admJ/
cM6stTLsXvaZ+iRgPIh9enuHw8yJlQFhs42JtdnCrE5obz/qqmtgYHsP+RP/jm2R
bvaqEhtEvxk0niSSDtDEqOlpimnJPNHwLw+xyHCXuKblwikemhz6Xm855uwfgRBZ
4AOXpcgRgU3eyzW9L7ZEju+13Wy/bOMjuwvrkc/Yi2tWTY/N7RTblcnUp8NQEF7S
D9VvBr3goy/8vFftUIr2LdeYPWXsYJZRTKxToZ/xrEfbtWF4rB8CCwum2gCRHn8Z
6morihN60SAkrEmkhfXtGLt7mG2Hb+iBkYHvmMLYOn029JrRJoogupX9Zr+1wBwr
bbXYrfQ1VIhD+GrFxcxFFjCp3uQlyDcNANq4/RL0x5C44FGa6zR4/HTpdLcPbaYV
krRfM9HfNvVPmXk3Cdkais5oIJh+6CiRHreKL21Fk1tmvzq6yu5AYzMpF5mXFGz/
O6ALaFNfvZ6K8uLdTEZqOW4SnEja6isYUuXuwPEu1CKTdxH5TxFOuWSM3h/12nUx
pUqp34w9kY2eOv/a737u7OosTAIrBfd3uh9XTwF3j80sGMCF7awJkpiV3yCUXCD0
yLLOY8PmYhn2ifLQFdaHohkJyi5Cgfr0voSNJ18Vjyn3wuYZeyjqZ0sG9V2FECgV
P5Xb0yKxOzaynYTl8xIy0ZJXDxg7sDsy1dS14qPi6uVyZDcHcQtuypQJmYIiYkoL
rkSwr2EKl4pQuilauB2ZZM1sA69sceyh3gxzVfB4uU4tX6ewJmM8QQk1bYsualsI
016Qqnv+s/CI/CuEspjBhe8IBJM+j1habbwYVrg7gG5OcbCcrfZWKyuJGxQvdztx
7ND7Ndl4DCb96WmWs7NRMqxfsbP6cPYwIAyZf92TG/j/4DzaYU2zZeM8BXC5KSIv
J1hOADlEdoulTJZ2Jqf/Mc/DJK5+N10weHpk5LSWllYjstYIKszgewv1pX4sRg67
hmsS9s54pf5BspIUznY4S72tulook3S5PhWxLwhdpJ1sT/TVVQAYERlLgpLoLxiw
GaKvTN7UlRMDVK4Z4vrX4OOXVBdWOXPgQ3uJZQMkXDfH4CEGhrXhOLqVd2D79+/q
4L5teUQJmgH+9ByikuGrKW/eHAFnmNBPi7770IJ+k92Yi7skAuCn1e/i6h+U+WLv
G3QJzUN7IC9QYt+/zyshCuUYDSyjEMmVKvNB91fmI/cIFC4rpeXHP4/9ijegfPq5
5pOpF9lTqVwPNSiURIyYlqxLe3KJ0Cq3+pxfSfgCNJ+UvEuvLTbpmd8pSdp4+xdO
app/ZaJAtporxkElt0ujsSF5yScjkDHVNw69daNhBrOW2VfGw6JPe07xjZfb2nfR
fUodsNPASPBHqoixmAPTOMnwmzJzcOL8VCwcwJtcyjYSPFZn3QL4LZNcsgMIwLq+
X7TTSycoj6vjDXXmS1nMCAcYPV8032j8fHwePk/bmHJmeOGv37Of3ipRjEYTT3/f
RIYOVSQ6qURGNE28CLVU528cY3T65J79uD9dPpve0VZ18g9zghOB52Az7AMM5dgT
2LrSHg01yYx4YcE1HfIZmG1LioeF5umbZzlKomEkxNpH8U9GKn8povRA9XnAp1Es
ZJ2PnSI2Ff9UrxeQz0sR3zSjDUf6L+23z+Dp1N5Ja6uUBCs+YQUAr7sADmsNh7jQ
t3YrYSoetgBdZO46tT/MqKIahwn8p2OHJasME/1RpxE7izYXZw8LeW0iBzXAiweV
QR6rUoDIDtENPGM7U6aKH+TDETHdBKhaiZbNAsT+8PzzioxCsOL+W7u8AF4mcHlg
BbsIPEygibTW+IO6kTjdRv1SIxId2xN8pqGozOp2LsNbkfodahvmCreOzP3Py7jv
MiADX2gMgp7opOMbSCihNSTNN4q22veqCPJiumIySI+fuj2Cnh7vitJlmsDd7EDt
RRgPlSutE/7ma/0PNYjBy0YLWLlXY9V8HITR0ud1PUrraiPp7i4wGcp9SzCl4hAv
3sHh/AuDeHv5euoIFTiLeA16MMayzPTQP2NHz1ltppc5945Q+b3ZCAJrMpER8reG
PIqGo4RBuiz+fVEIXHe2Jwz+6eCW3xT4V2ToCJ+YkYSy0xhS1r6Ozg2ZabvtJGA/
CrniLN0hlmHR0k1vcK8okFtSi1jWU/QJQSxn+e+GfYCE5njQ4/xzrAoo52KMP5kT
rMz1JvhaIN9ijrzi7P9oUCBKgZgrPyohsQc6h6pLz7SzG/vLpdAqRSM7niQ+6OPh
0hy9MfXBfWbNSgNeGUh+7uFFdApB9zRXaZdNSikulNwtlhxm7T78xFLaWSJ7pBrs
QC9I7V0kWu+LM6cUC9cVPt115KT5scwzPw5vESAhXRsbrN3+mDsLSJ8u9e/dAH8e
1mFv2sHPa9kMp99YHlMcC5/IMkufe86EkVLTZMb89+MmVfNYpQxisnoKIlB3xBSs
fCbwo/7+/jjMZd8ugdfnv52H6mP+xOQS6M4pbmfZn565FPixIwiXp3ro4IbzUR8P
IdXpYLZotAx5xDhwoZ2J/W/IJ+BARy3aY3kn6Fs8NicNjOuvXWtXe3oNCfm2sGT8
VtNISw7Rx5dQrsGBhiJwm4u6v3zDtNSB4fWEmpENkHRwsxVryedDnjLNC6E03CxE
lHaqnUA2r2KJi0gIgLTkmB5SQ+iwOGf5l28hxgczandqKoJJpPKTizAqA9HRNZKs
x4ovsfKtE5dKwM83bp9XuTpeq9TZOiu092yKesxZZfrgvCetq+LrfKoa7crgd18W
SwYQyuB/IZCurFoCN7utNuWVKbsh5r8AdObi3hQl91DEZB3rNwDQOZFvtv6SX8u2
89ekDZ82tKb5Ppy/XdRBBvENtw9P6iQiuJq7fjlP/EyIb3aRKYmXTEFN9S7Gl76q
Nwp5qYlZvTOdtX5GMaTs5PwhA40xcL37LAKklYWKSwNVedriGb7eLgqfQX5TNlDe
fbsNscpOf0cVBVQYK+7EbRTOjJvGSCvxuW1UJyzR0adSEr+GB6oKwWjs4OvvnzOM
tdem6dRlxBFTCsCwZwr0RD8kusLt46HMHYUjppzsRmxpDZHeCxbDRH7abWPmGn5B
GplyhPm6tunuxOpKUNM8dwn/sYFnzSyIc6YhdkRqx183lG6xPx7gDU8KBBy8EhJv
YQoDV0GRr5aP/kv/WHCk6H5CV7rEXzND0+R0ldpkie2p1g2sZD8lkb1X+3AQdzxt
bk2BQchUzwvHBGIEBC/qjo8GbI7E5iTzbzj6ocHDvehK3Wa/o72awM/g/UwD2myX
M0odWMNb6UQ1+/UHCkfUqC6J2ESA0HqM7rkzCFcahByWC8L/lbvgCPMZrb0glVjg
LzLWdd8LO1ITyshUABS3gP+izsv8hd5TrP41HH52hVtAGXXOseoMHuBSvZj622G3
tw5AumYtlZ3wKcEsCboCaN/tgwtvw5urUIj2oq6BFgGfnn3t86qEMybPjdP873uu
R3VtYgEvHu1jhFikBr3DVYiEz9ELZ5ZwsmgQKhUGrFeWCavBpcKeGyDwWsPBzq6C
l3PnNfWn/Nh6JXy089Y8LCWpy1/upVRbHPMR0UQ6C0oojeqB0ZvqGsG6cuA87i4k
7YnM4yxHNBu4+ZkTM+INjpnGPUHM0CFPNpbGx28mp7/3h7pf8LcwJyccrFtjEXwW
KPo2TRVreHV1AhjK/qMdzjqEXTjeIiap5elaZAoSy4GCVANYwEw4xdQ3lLP6LCSl
OeY4LdXncsx4oQsPMjMCPrCF91eikI2T5m6Sw7w2s28aLDj7Ugm1vbpQ8J+jXbkC
+4K8+eVCTxUBDnIaUohBcGboBkW/cGsnt1Ikyf5MNS/YRKzb06ke5hs6aLTC2Lzl
KSEX1YZHgD/gwpJpKOIF3UI49MRV89kJuBb6HpMwR2QechuxQtfPOPOOylhwwApM
aslMeOKSjx/BIuQu6iqY95THLb7bLNx7YM/ulcFNc9XyfdQ9rxzWM98uNyH9Bt1s
wYw8K3zRTNZeVqHpPOs1p5bH7Uo4VO3Y0rznZsR7bk0Hby8gadk/4EIroUD+vVvi
tKKcQu+tcH8Q6EgGRt+1vW3UqXni3c+J/2drj66DKvGb2dcvDFS+iXj0XJG5ettz
7DLTKCEbqlri6fJDo491RkFWSIkCVK2NPdozhQy3d/3gTqAwKH5/nbxUNqa3/i2m
TFwvrjxoVrnVUpbokWmFL4z7Zr7DSs4UbmD2XsD2UvnOkrXWFbFCP1fkG554quz3
i0t9RYIWwvkni6UL9nKLQf19VRm6bUMzsvKF1omydjpXd7ZbQLox/BKDPxbXA1ZZ
VIaUM7ym9CV4mRYxiFOSC7zB4ZAaG1L6pKts70YP/wH6SZQXPKruo51ecm64VZhb
PFKmT/XfDUF7NgMA2+QEK6zP7Gb/bO0eedtQAKC9mFWePeCDFRvWJmASX4to8xcO
bRIgz6aAE1yntJjfX2LCB1DOgatWWVJHPH+BMrh71oxbAdNqKsKmLFoe2HIfwxZn
BA1pEFRuZm19zkcLT7lQ1Vi474z7zOCuMu7jlnWtgnIBevwAo5XyV35KPFAuXXQ+
4Nnl0clzaQU3hUCtQRDp6mhHslYwairjoyTD786r6M8QeKolb32S2iNtNb/2dUZT
0Wa9gfmzeO8N6TXgykFs2qIBsxtrvWlpQAlTAa1ErXqGyl/9XeC+Md750yYSRRGQ
5rqJCpak1/ilw9H10rGGTjUem7yQ9MHE2w6ZLVUA5oOuRujahFNKonLyVqTT7tRx
paWaxq1Ekab5Ij7lD5Ys2rZi0kAGftjtWM2zrpicfx4sUvaffoLPSSZ+BfAWbMho
6RCgaSrzkq0NUkaaeyFGMsQ1VF/cVjtNquuH2kC7iJ1/ZazCmd4iyk4IFFZEIx34
dVa0otn8RrXS5xdqdeeL51mydqKdOd/anJjFjt2lzUjEMCgkbHThRYIZtZBRnfrQ
SusJTdKa+ysG+qrJALPBpuxgXQZC5I4a2Ruv2afjmOqMS3uKAfVq1ChP2rzMGkCd
FTIzqXIRX7vYmET6GdINSWhcYQGvNiqzJoIMPm260WBp5MlQO1uBbMvRc9lCNZND
dRaVhHxsKc+LAN3P8f7/pjHlByxhue5g/f2j5UWHYPWr0v12M/r7Zz72KbKHflld
Y5kHpuDPU8amAVtxXZWNH3qdEeRP27fT+Npc5Pw0HRSs8T/HOGTiIaBe8LQ7TviP
0/jSatMP7JpfJ8gKmYUnJhRFqPUrpWqp/y+NzTkvA6eVH1sVGIO953ZN0la3dzsY
gZg7ulQc6o4GjSXcLInGk/i2V1mqAAfKae/fOxPgCUNbACgTR9tFtoEaqbDRuc7G
K7hpGKzHOarJy3JheqmU4b3UYeRXNwq4ZfXsfGQJcwa4n0OmhY35DK5gzycb6Ay4
qwhvdRJ10SCPmaTN2Q32X2dqMin6+Y6+N0ULlaxXZVnIRONMaDllrRuAxM/2F85S
J03Pn74LiV0uAvN8A/Nl87rTP66H6Eq1ckMK1O03GiiiqC5kVVEW0/Pk2DuVIC4q
b2+pvHGFknRFyq7g9Mm4YA7mgRpldr72aRUw5tZjddfUBtvhf7jwxX4kj8FvOE2C
BDJzyWZJAtNH69YzznTL4PpG2joAftJi5RhoSwez8ZBrxY3FuX1I0nXnk8Ql0tte
E8IPjrBwd/7U2Pf/O6ETMnFNWT0WjxIwAO0dKKehrvLDGKLfcfxlxLVx4b5W0c70
IWzLdqSJxO0FTnshZ7r2VrUeYR8/8O4qlj7TjWzy0B221rVVPdBabc+C2XPdAqGJ
m0VtyY+MT0jHrSMtXKxA4sAwZeI7SJJp6xDRA3xL++bEGhEvnT8tKrVHgUZ9XArF
rUO+KQJ3V2qpwdmWB2w5ufo8GBr11r0HkvN7tG9dCJ6hXRt570mtz8UgBEI4cQ3T
1wKbriImNbSnF8YHqu9YVYaoN2KTQE+e27a5MF2ITvaNog1JEsbTOcxvfQ4gL+fj
3N6O7TZEFYKoBDCTZAXTGFr/IWa51TA7UFEJXI4izsSkgdJr50Znq9kywexJ9j4O
CPqNWcVFwxdoYhUCmW35K86Ytn72qDcumUEXdW507Pi8eg0hW+XoFviWwDHkwk40
bRzitvhQHzn8WvoZMSUmIFY5DAyri+LBo26hAyZrGBtsbulhUEvIRuNjQCY0RD5x
K2I2O6SLCUH/aVJl7xj/sUOfjqmyfuxa1Uk1amE+CPsaIHjgGe1tWgt1ziu1iUqd
vXUWdqBw9rHDUv2NWKPRMhrKgD15PHwpBlnwYJAwxIBkcETUVPDYYqXgWOwNrIRg
WGgqJaLDe1ZT+C82AyXt4uM9MYiFKiFeo9JecXbFbo0qXfzYO/xF/Bh2p5JHSz/l
HWOXXQTaQn+Mhj8dHtbmz+sGEX8ybN5+WWztht90H0QFsdrJOvQmA51ALcCsjZ/p
cI6hD4dNOQvD7aBaqsoLNMBDZuCc+svjMSzI6txOBamgnD5GqE9tPCAvloXmUDrS
yuGGcWnc10miirtkLn2QIeMxa5EMU/k5n7NpwJy1DYBd8ofLz4UOWEu6ul59O07c
qsEucjoX87CxNmUJbSEi7a+WLoPbYYbCeiNReEHO7t7njz067fxtA4EtNn7J8AJG
ZkXODZfJL7apaNKL0AdM48/SSegsvrFef1rR1C0ZbO/gEIu34tNQWl0eSjI3Tquu
VI94PpV8BK84/eGU6/UkRhsnJGTHDjMHv5WXI7Y4t1RTT3zb0mso9r7UdYO8+Fo0
9cReTAlrPZ/sj7pr890/CzuG3H5FURWcMzagnWrfsTvOrPyWKXN1AxWVta2O9/pc
bELefDx/afk3l3Xk20A+rNClcvDCZTUA6HUMrEi7PIAhp1Ek7U7kNtXbH0tUZcGN
R50G9KNuz1usdHIcW/m1fIefstLlOz3jKt4LY+0kT3MwdbV4BeZkpgjstBWDDddd
5ZqwHutuZaXMDPDzZCOGhNgkuNhPdvtTwhg99ajqbb4QJHzW41uaQD9KN2nc183N
T/xFJhkbON6XNpXifSyBYo7a4gUX8mfYZTARanZSEsVVAY7Uq3bAOp5Opt4TJDOr
dtkM3TtNCWCt0/iuLNzBEDlWuNlfLbZv1kN16bRlt4dJL5BmENijGyNTZyx80JTH
JaTy9EXPMRAVYNGZss4W8Xegfk+l7Qo0NeUQGNOdrl75k4Hc2W5VIt8yjbd4mUsU
97T0qEO6YG4Un6crYKC8jNCE/Kmz3V4VMIF9ct42KZ4cMZWFlS9YJUUD+bFJp2Sb
p1lRxItJ3rLHaLpxyH0ffAd8quCCDGEGN9qZ71Ep5ClSWSQ7LcfJ7wVtOpXC+mKx
NfI2EKCF6nIT5msOmGZK7VV6oxuKnBA1mH0ojVAVLQG5Dvl0vjy5uL9UMsQH9B5F
4mu5DMAOpUHX1JrJY43bmhWW1UxfJ+4/tZ+yam5qkSdTFI0QIP1xUKS8TckLTY24
htOBAJNF+Iw+781peh0UKUmZQ1wfp1NGt4ls6t/jZFhDF9h6U9+qwW6Ld53u0SEW
uqtDwAbWww2QwOwoUkGT6L5o6dDADgmoAG4f2Bwz9ql30D3BiLtWaWxxsAqNeXZa
MrfGggR5MovaBubWfSCa0QoLrHMkoFg61YahybmPgpYiW7EwySyMMrcwW136lzhm
xOQGnuaMY6LF27/prmerhRqVrCqwtp2kdEKyH6PTimMcFrMsm1XoQfM2bbl2N/t9
N00PEoKAUONQeLrjI7dIHMxW9lJ2bv0YaEQwvadF8Y8MTR7VGT3xrgq71Ekiw6vg
T6GKxdGyiDBiLQRPemq8jaIITHXvd1AUlhCdVOWXBF0Rwj0WpyqiQ9Eo/WXF6fA3
DLV2xUgYFRGZmCXAZausZsyYyW0vBFvl4jpshHVyU8i4J/SI9z4va0kC+j6ugaMy
/hrQYBfPfIi7JY/GU1Q0c37YDE3EzmVVr6pCz4aNHF1J8s/GZL0+0OobjcCdKVw0
RrTyO2DvJeZsrPlnVnK8CmAYbVi3qsiq06Rac6DQNSpgt7N1TgVRJ+VS0eek0fmu
kJw2hBe/m0QayOidSN+M8p1sJs48p/GQ9AkWg/Rmtu1iQno7uQo6TsgN6ufp7rLx
9V9aNUybUuILI5D8DX82g0IRkoXg862eES1fk0BQzGk8438inIYnzunX2EQeWl6d
fEVD07u1zccZi0+jbKjomaJ1CdVRAXKiOfR7zlqi8vMn3v/Sjq71et5m8SE27F+Y
WEOQVLu8O+ves/DYseocEmV2Q12i5sSl/mA0mcH1rX/E68fAPTVaDICqhXlyoOe1
KkUGpzQYu2oegOgAc+opohlZBbbqgAdbfNpZQfGfpzoyUUf6DKX/3CgqIXSqugck
oFARCj3rHe+fjXmFIjsXqq4WILkK4RUVkosXR8XX6Ixmz8gxOItvUiGJsTbasfpp
P9TtznjQveSy80d/7Xxg9GIzfVG/GE/DxIfZvcMQxt+ErN/3dAYmiS6++sTDzfSI
9x3vTz+KAKXD9Hpabadx5KeQ5LjX6sw4oVir83J583wkR0TUBiZrifhYO1fz/fJP
/p4dqF0xp4ZjPApJrSrLVWcLoPoJak2iwMivxUTv2w1VzBhbuMu8jqupFIBZjKE7
bnKyDKk54bvtVg0XFjTmfJ0a0MPbCZjUixHNycRdQ+jelDGQplRXEBYB5eoRu7Qb
XPzC1xdRq8qXNvZwNNiUqMpQuXvRXY+mCI12ZqKlzZ0aRwB7TXJJaZKSMU8LnjD5
FeGtztAu588OvxJFch+S93FCNTD6pI+K6rQRiEKeFip5Ni0bqPdzyi/bwhP5hrtq
EyuXWMnnL6SRkSu4tqTYTDEqWYEO5g+mF7Wh1UF0ag7sI0h4PyWWHKq0Un23bfYw
SWiV25kSGFKhKUDi/BHTjzEljC4HxilJhm9Tz6RoNb5x/4cT6WyXLF6p8GLQYG1f
w5OP1SxeOfp45YEw97aBZm5n9YYLh9g5LFIWkg1OuSL0+ZQpkYgy+v8GIfmIzBhR
2WX8mAKSg69KhZm7kU76uH1avIYh6iGcRIBOsIR4JEF6KSKDImuT4B2t0RiqQAsD
k09u1d0dC1SLlFsrgaPg891aiHVFjJGuMWUhseR2Yu2d+bRfVPOUzz/6eSSb7vBi
5mOcp6lE5j+PaZbowPdSeyX0AzPSulHWaPMmG4hHKsYH5bfiawzqwt4zsolIdrqJ
A5JkRaE6ESman4VSwJJdirA3FDlUyY2qRy9d02pTdfUarr79bWvxrQiS6LaYBzlf
QLhlXCMdPwht5BLgIwpKbftiBwprWhYrUoRNQDIZRdkkN2SDM/BF6CdnSIAt77mu
5ADQj11MZAFnqyrrKHrc/6Y9ppUNRJzATWBG0Mx0btFTYvI9h2HGBKJwaPKMGu96
x6M/018IkwRa3wDKFnNYwXO2vdO9UiIwKk0AbbURd2lMWp90mdt7z7Xesj9ItohA
cF/JZy+h/o5p7V/moJwwgkfT71ZMglCz+ldhg0Gs++r6CJUyw5+Smk/xo+Eyf76P
6GmEJD857A8Pd3/Wa8YdCcKxhgv7CBYmZiVeKL5jBktVClytM4vARDil1tKygorz
Ztbnh6fTWZoZf0hvt8vcQbRgrt6AE7EvRK9tVyPjJ2NEyWLEuXifOQYYcK4Lme7v
m+WRZlxkobTqS0zCVtbnTNLo1SYYh20QqzSwfj5xa97MOoR4XeE/nWwiVcCk4Eoq
53WeCIV3S7Lnn1xkPsojF1mAWebJAxSuJA4g+j2YkbLjLzkSU1ovKI53uJLcgXFo
3PQbSn72gDcKWS6KY8mSrCH7CVT9d4+gWZXuEIH6G9g/qAKdUTemXqNyXS7SjnrO
3hiSRiOZ6DOARqI7GRvbb7uG5xzAGG6LPSdYbJYFqyaWBsCGH7rOJndNnTTZrUzI
8l++TYehv/J/5xe90YeGHrZKedVjkVvuYzBGWsMMtZLi3AGjbdDRQD+df4oRZIDp
MTENdnAyoxYoC+p0Fu78FuehTdLPRYBB+2bdijyo4c4HbTr/3zmgwlJNFD/qz36p
Fhtt1w8A5VWYC7WF7CgDaZp3fZL5gseVMaNviv/mipzn29EPoCH97993XCFHMqih
ymuFYaxMq4hV3kLRaq7owyNgfyx27a68vt8Qm0QeYtHjIuKYew/+GGNTF04FtMLM
9oDpob/QXoxpZxFdv73+3CBb03HY/ldzQCxCK98yhcjoDOnKa64ZHwdxgEY0ohYX
B4s5C0oitaVfJ6ECzABdIHGdHYBzTy+/QaZCvAul8i/yvo1SKpQKMnUBgSk9ToJW
NzKgNuVe2w65aJLbOBDxdG8FluJinQzg3G28E1ngQz6TgfFat2TUzVAbuqCDSP39
J4qXuIrw1ASTrE0pnLTfGnkybpPiWAMjq/W7MQQ2dn/xOs9D0w9EHrpjbEaEiTRo
cZkvSqpvpazGRC5SPWOgg4N37PD5LPCkbdzLU31SqAayyMr1Za9A4odeQ19eh+At
W87J7go5TRSCjrW79OhjeLaONXvi/WkvXsO/SWpjab1KqNFkzneR9DNNdpa326i/
w63nErJ2LGRvnixuHUjNIhf1/A3TX/yr3kNjT0XqyaZ2o2dnpAJL/h0BNQHTCaAU
u+etE0WRX+YlSCP/bZq+odKwWFA+cPnWn0wJJ8RHAcnYovAJWkoHwf0uX4E+1QqT
YpT2157sCq658Xm9lxWdsiCDhlj0FnKiecH/JP2BQxvE2cZRkcQB1+uchsrjCcdY
bSrieWklmYTXsQkUe80CcFj7bu/PCYJP4Lv7IHLF8T+5KaslugkyG8qaXd1gEETq
PK5JiVfVW2Sm7wm0iAB2fpigOZaTud/px2QTzNi3UcGs8Rn6FXHaJ3o/JYLkwNZk
VcmRoOA3l7rhJFu73v4vI5YXBJ9AF2IUsnzTELCFn3NdjwjkcdF7UPy01bSMa5ta
Lr8RUwEHnZF486GlGiOl8HUOiMqhk5RGoQW3rzPDNHpSGkYNzHtr6i7Is5SKKhzk
H7HnkcX6Zfr+dQAuUfXRosbtkOlDjF8nzt7SNrIbMdxUClaj3sZW//FOOmnrBZQh
xWP8u+w3UGwJ/xwkCktggH8UPhsnav2zyzBIcVanLulFUqTCpU8lAyeGMZwYWC/f
TwVMAj+52Cs7hG9KzhGB+ecqqtDr+aDDlV+k/YILK/j/QCiFaWkKUqUSed7ErjoM
3EzbPtqGO4cI1FulSiUddikDei7nlEcY+hkK4o3VyQKl2ZN48fi3kkreK9s8HgNH
ok4+YUAYeRXuNoNw7fO2D0xPiLXAGPC0iK+C3dyl+XujvtBdP9pTQvb81AAxBtMY
hTTslzMkqjoDJQYa5oG3bINz8J1aMHZahrAmpZks7uuyAcn+9jXojDiUR+M/nbmT
zLZPMCKHLguXwnTxt9BBzNRjSNLm9KkFL1aP+r3yzlK8fnHHGrbTql9jcoN2pt9G
1O4A1Jm3EAWK0Nueq+8cw+D0Noij1zH8LfL9ducmKBAZIatV2PKWN4S6HUiMUb3+
0KVn00Y1iF925hkn/lVapWWCa6VaLV8REr9spJDGvtVWZjpona9ye/qqpbTEjHcJ
GTWoLsbMYcH80jBfBUfAtFyLLF/UDbqCwwEHkibA7GFgI+NmzmGW9Y9sv8n5Tmk2
F+hwWnUlgV4iBAZRDZCwvop4An3l9864DqeNPU8qEp7HGjJ2PR1snLS2nseqf2ig
GtE47O8cPbAx7uPStro4M1ArOES3R+HfqT6B+N7FGEmL1g1b2c0EG/cqzso05wQ7
vvWtrslFfDWuX49oQb8M4txnLAkXm6QpaOLxr3IZeXQ7FWBykhF7PB6ww+15c/Zf
0hn1/B61eMCmmmCLQAhD7VlFVFgAIOmh19L8bsm3N/fgCCr0pSjX6+E++UBCFb1y
K5mOaJYxnMSX8z/J5Pfz+d4P/PTgGql7Z0aQPpdplIO/8Yc45MaquRlnWqrVzAmF
/ufVdG8oClPvhr+557no/9xyq7kOkS4yF64ow8fz9uEV8OyHGA3II+CGSRmy660S
uuaLlLF4OFFXFa8E/pKJoLjKYfQ/MgSrVHeUGc3lzXjKW4Rgoxu75wmUQJMyn4gw
KxJ40cSUIK0j7AYfzm79emlng7k4rqK8Uy694ts6JQC/6HZg28t6Pa7ZBCPFPyLh
RbcUtq/yyOHJZe8dV7pZcsKFwk/QRT0u4G9kSgcnCC30GIrtVT+IoxkT7bI08clk
dAzFSLnBS4akmywylpSNeN9670Moh3rSyAeoBNWQ3OcV+6v+2TXTGRdHhskYgzL3
jHQ+gYttP29k1JouMXvghYRzZAK+s3wG1p9s+fDbUUQ7BT3acZE7nS0EakgftVGM
uOnLLYW0JmaPoz6RGMWsu3lvWcDzfWgSynnLWe1t5lokY81CbJXyTXQV6ETysrBC
iq8bGW2OCNZ/R3ZHGVJrNjF0JDwp1NLrglil+ocXGXZS8EkS4UQnmGnDEttU8qNe
EqqCcVIsCNEJwHEwSXegaYHgltfup3HIQeZjp3Tr5CHqUmctpxYnd3i3TfbbWHw+
WXWoHfoWmYirfRFT09FOgzUd3oRpGXwC2WFCgrET4O7ECDbgLT6LVCgItCFNEaXX
3R3I167Z2BxBvorv/jmDUi5CMNV+teNWlVTSTrSxUmIdxWmPlc+8BOnHNFChJCLq
HXBjKaE5Mc5JAlBZwF4eZlWmKS2NH84THU6hi5cYUumf1/5rD9u9kBBhX15Tn/qD
lulaPul9Lp5Fzkx5IaUmb+oqsvTZaKmqtdeLPYKNU+y7tc/TwkLM5vDrNGygg3xb
+CPZ02BLb8IN9sD4uador8PUOch7nd2GWeS8O6rXW+oGKc8htNnxe8+ehCVyymzO
UH4xHA04GkqX5EM2BzHY7YyoKPfgCBw3jN87DLS20afMk/pbu7szP+tT3lyzXF7E
UtWvAzjSiMRzDEGFFcfj/mXLFyUAw29QOcgX0jKbIw/Va32a6FbWeFyz0tTxug3H
LWwIe/JgoeANsDe86mBiuVK7doDj5tzAmu6t8pNeffc7GrpPGEmIkPE4un/iCU8h
ck9PFgKgPaqgbvNVKDDmgYdwoO8VvDp+vZXbmHAzWOzVx76ZzTxBp/lFKiNxeQpA
jlhxGAVvCyoR620DD1nXdx17IKbdCuV2ITkH0jsSNYwK3zBE78YHW/a2+s20tcpF
tTIx8XmS5nHhdaYFx2qGSg5n0rJg+yMNM+u9658WlBQBiWKvRoRDSeA/VDTNfkCL
zcz2nQe1Zb/pMcrSjTEZOOhaOZ1RtVhuljPtaO9jcVCcTxeD9mpXqEkBDkU8RBfD
X1PopUgtrSzBkchEmuDDrydu/sGMoaycCS1+g18V5L6TrzB0OTsokflRmGyw+2S9
6Z99woB1oqNOGRGxvMpTc2VcvW21KHac/Uu9iDjERK6NaKQ7DUS2KsQqXZTiNG5r
IMobuoL6Iq81EIUaOOo3VcloN8o0g5SVCdBXPNtLl80+r32WfyszZAk1upDi9nnr
/Gp45GCgW/Hqj9llEv7jEnn/ZD16eRnA3ILC/451c/VXlLEL0PVyxinMGdUPWzXZ
MOxfv6VYU5HNBWi3PFh704UJOfICAXIky4lRnPlvzAcuO5npEyIXdyrIjylfomEj
4a3umHwR1BCT2yjVy2LiWYc9b3ziS2ZpEO6kEoQzgZfuJhOtKzdwhRGnQILEddMh
fpvjR/lmh+S2RNaQIlBaCXyKEeFQFa9LW0l4z6sYsq4uZ/HMKA1XGSKt0DYpoCIK
usiiJKtfz/wiEjhLlVgYmSIIyQwZ1DMHU5S2UBwWdR+MWjgE8ofgffGGZ/cRa7ok
j+nEbko6G5Q0nkUWkWx9Nbm8CeS5LJ+0/lHBD0cl6KsP0hJk5grYvvKxwe3t82dk
tdI6efoNZ37HR6QJzZ2DxFtTmQhGOEFbkju9NIwneVqqPFG2Xp6Z9GTmmYOHThGf
BZ9rjNdyLuKIuR1QK4oZOGIvAyEyc8C+ImFgj6R6c6xc6Vv7i5hUZyY9WJOrfW0E
6iEtUFuQDuGzVx2Bht5dbehkSAbll04uld/m8WHOWPlG5Vfmahaz/Mp4B1Q55AS2
nMdpm0TD9IlDfDxCZOmMt15tr6qreGpdFQaNcBsnM95SnJDi7OB5uh/Wx2m22qkT
EGIuQzxJoQ9Y/6VE7pfUIgr8bi9/xbPlQJxkCD/9JkHrhdrG/8ZspVaxNTLYelBh
jp/KxAIeOIXl7UFBK2p9B4DLpSiulUQimMr9uUMdBOeSEadpbr8PFVZlr6YRWBSq
9ggtVPtDYdZ8oZqCeOVIz8TmmJHZox5oSYDlcFXybLLjyJe+aTphS8n9YZLznxQ+
/3+yjN17by9ctqmCgDxK394g2BcUVbJZzPf9hikvwcgx2HOZQN+6pUfDBj4aRiEX
hfXMoZOrtAbOoA+MtuJ/Iy+NsobbuQVC/wRBVKdLRfbTH0I+ED2S54hXuRFfPj8M
Yd9+ts4Fjs+6udgw1OmwOAQQlZDE0K0094ZCQaXulRRKu9KYH/CZo06TYpZqQJdF
PCKkaMVrMOOWg4vQZf4V7wrzHEgVPsjAW5+Rr2britT/TKMtFMJoZUqppBMANNyg
BxKdm0zku3pbKsSn+ksQl9l1FOw5BrJmTd67bBCKWj/qkqehgFYKEp2Afq7bjhuZ
dI+E7BrhKXq0vX+M/0Y+tH0O+sWk8zUWoTBdDb86DCah8CGGDqJsvC3SxOVtdfUf
CarCW8LNe+s4M53FTMxRsmOlY7Dr+c+nWZc0/is1a6+vxMJNk0fHuEGQ4jVjML0M
LgLVpf1EjUqVMBKqlwfLlSUC5mKHoVXIV9mvw34arqkmbIC9qPhs1Vi+teZQ81Pp
2QKuSAs/dsWusH8uW2Qi92SenOVE3v84922KCdBOt8KAVkH2r2v4YnVlBlqa8XK5
8dQRBQC8YZoJmhgDPCYbZvg6Tk8s8qNBZK/hbXgB51ro64A08/d4wMxGpEJK1Jyd
f6Rb+bDZiImGt0W9ynvy8PccU2nfiYf/UuckzUKx9u3bJA+Wys3n5CCRJooBeSM+
ug2uQnUG/21gm2tx+ICbH5NgpINfCPiGYMdpSFlm6m5J8k4jFYoBh8b8TXjE7YiK
reFJMj38vHs+oq7SEBx62lrZWPfpG1UOX0LmFkCG0N0cZjp+nosWnOpR889ijFaa
q8XOwrCvgduK+iZyOAGOh/JXsNOAG6xQP/vWWiA8e4wMZTV+CFREQFxr00Khz0cp
YzMw7uT3io3TwP8HdU/+oP1coeu7xtpnLjpcdS/iqmIhSB/nGc+KOFjSJvsBEBnI
tHoTgiL4G6SpvLSE59DBvf0EO0OQe/sG4i/uyR55u7JJPaMTS1p0K4gg2WSZceN0
Lfg4mbjTeBeIQ9VLV1K9eSCyeH+mf8SL8XPuhaMxlm3BNH3TOOib7t29m1hx4ayn
3pdrpMKP4TEThnUDIvpULNIzF58SMbQYcyWtgcZkBw9HlYyXrrs1pSRUiuzOMkB9
7zkdHauPmJUYhMU76WIkg6YwXCGnxuKuuD4Um4ghErhvgadsL07TnnOHaPMEKrOU
faztY7hYXUQO0lSubRXM2hUoJ2pH+AQh2GnpUAPiB/dA0aCMYrQlQT4Zdky/Uw/M
p5KP0Sb5BIN4RKdKkvLmWPyanjfngnBixr6GnxMrjhHJNDA9MgTYkILbwyNJNZWX
872sieqF71HOWIPzFG/fy9wOZu83MOGTgzVQY6TgzDPcq4IbRmRPCTqFvgmEx0Sv
ENKztyZkgyFSVUCxsgcUAe2ljXhL3QzeATGHzXTcZE1kEugQQURGoo09c9dQ78Ju
+xiwwTttqBEuWv5f03XN9FrJpOiL5PVBXYIt5g/iVM0x1ORCbnz8ar4ye5oOlVeq
6Jt4CTpU+wgROpNELxM+uTGf3Ul6DBtsG+5RjzhdR6xh6BTj2Gf5lsZMOlBW7tvj
RFHKWzyFHW8ZHhNwr6+gZvzvEtrbSoJyNapNiGxLHKk2zAZ+eQiw82Luanz6BOHS
SZODlid/HgHepIfGnjBQQAZgDcDLd18mc8BOWz+fAuZmKQW836WLbQO9B7WcBeVt
G/IfsT0c/gEtnas4XACpz2DC17Te5R4agyFxoN+CONgL225Y1ccJxsrj2l+JIXtC
8M5JSq6/6WR62rLyRVmjdKLpB3br3qVceYYyukD3Sp5f7v8JOeKOuGNszQOF1mru
fi+4MfNjPBuRLMKRuHCMjWKDD9SeG7k595kYh2uFqfp73WUqb3ggayR3YK/eTfZu
tpTkUb9bZphAcsZwUEvhCOU2u6E9ivPS3gf97rqQ5RlmpTnCMQIxoWMUtp7ztCYH
4wb14YZNFgoYqt0wAxwSvhUryAm28ZPVf5lM+awuhmQ2kkIj45gEM367UXulr02p
Zft50xclKAUB77/ipOt4uIUJT5NAnIZy51Ous78RytC8m115hM27sPkvmfBgcoc1
RVTxqhGZe5RhFOGwoASFLUtqS7Z9nb8q6qNAAiJ1uR67dKzQWBqsuQJpTK07lxhX
zVHWLGNCnQnB3mzkfeuBCoO+fppnvncIBiOgopfW84dIYF8HWY9VmN6WXKFSwtpq
YT6NJJbxKdL78KM/p0+OGmr4ykzZKadfmyn79P+RMUw2trlcMCVqNpomcPd3Ln7H
kTx+yXtT1gtlVjzXkx7xe2KRtJ6lD5+TyXmx0ZKa/juNSvecCV52vBOQA9X4+mzH
1MJit12VDKFVl5E36zyFjBXyFlpCW1NpvqX3rm7A+SgyoU5uSPfqJluidjmkMikt
vb6Wvn5E2YEK1YUfOZkGOOsBemwIEpRO3X98I4gHUjG4XYkg0c8OJJzS3ZSL+pql
MeyWYnQdk+4zKFQZ6TtHH/mhjseFvRLMpkgtT4uy+YTYEehixCDN8wRDbFEgCpjX
+e1r2wuDkNDDJ6WCHHYTJNh2Hu8rx2erRDW9maPf1DQug5VbLp75WWNQhSIiWTGz
CBFrjMguy4MN6il8PUZtW4HqECxmj1eivTYe5fMt5pZG/dizKORGmD/wm8OtSZkw
odRF4w+Z4qxB46S1rzpgpHO/8raKiASEdcwtAA22Nobq21n6q6aPx1vLbrkphCsJ
udS1r6cfTKP6iTAPZHPxzBDqFFFcT/G8QRydegxhLfd3qUsY/C9FomlXYwcqTrRW
4y6QjtDpd7JI9xEu55aJTGUmMR1DFvF2XSi5lGvBExMjA30H5TP4FI078glnM87P
Ihdw2YN6DOwaRb0m5cUvLDLnunJ1QhwLbXKmJeJI9giX+KHdug3DczBjU2mJgt7c
u8ab/pK2Bidm0Z6gGAa4n1AiuofvZzbyJS5TM+LyNuhSkXaXPdM96sI6wxj8jwan
cAu3x18EOakXYM34Xr6sDatOC5tGHL7DAgrZiGaens9/Cs9Lnb7+/dKPNWZtFGaf
QpItyQ42CuFkah86bZUiDqGQMOszf85nvvh+xEKPCo++pzbLawJzNeTdd8MNdB7x
3+GXa8Eya3YHxVYqHdjt0rrjVCmKF/YsXRypHAJ0DE0h+J8Hw2c9Y/DXuVWAgu8c
WmliKlRrkItWD+40SSFuMXzYtqXMK7PaLTuyswNAu3quM/Tny+4HXt/1/LWnMSv0
Uxu9fepONcx9QCvQATPlaYeV418kdJYHCAlmnxMB66tM9LPvwcfueTX9quxyXMOL
MoPxiFI/CyxWqeFaK/O2Z+HiqT+UMqcyY3JDKD+3rTyrhP96GBVSLdv7hVdXfzSY
AF5p1JHoplHcdzNlEsGODGwA7LLXdrMv2CTp2WfeWM6lxThpTWUfFVXXjEW75Fm5
ThuLaBdQluW6A1wW2B9V2nJbu/1FpDgma3ABjJJEeHucacVXdm5xOa2jLrxa97f/
hw0bjE/nJ99ulac2hXhbQ3KVELc/sm4ofIA6Y7FYwIa00LHUFrw+tnstWas5TMtv
7hDRbj1wTnHfN6CtcHmdC48szDSl+CfJ3r9kvyWS+wxdJpIbS4RYpBmEbZHVGVbF
50yF22v1ObcXmy4+3+MnUN0lFhAdKYxLcJLP6Mo1MNpUtI4swKtBxzdfqPpm8sDP
hpApHcxYU0kQGBT2Hm97AhCxSw6X/rSAnAG63rLw9/rc+9GhdnmPZ1MEWkuv0XlV
zwwMm0R0n8kHnOanOm+3PCinRh4NBTGaEJE44EjzuVAZJeDcdDiRxM7kD4WL0S8J
8VW+b0WfwyChvycKSQ1NtEMR8hVlsLWeIK3Y2Ke3FzsmNSZXv33D+jSeyxtbax6Q
OjhlTTMHQnkTxbiLGoe8biXoxwRUOJ+5rpNdcCGq7ru5UeZ8kk0HgtDiiR4Yap/e
t0sqXQhdn+qpPSC51/KvMAu84iGz0SnIchM/2TzywrDagCauk6Uokd+g/QYD4JKY
dFq/m1e0LaH/F7/ALvwcgFVhL4s2U3JldFGBhjZ0QLbwkryenVC6NK3QUFuKZpIa
qCc7cylZ1lpMwlUlOZWOnnIs7/5yPiuHwgaRPutQ/y3gYX/52/lmOoNPQ8/0Qx5Q
458w/JDkU1un5X+GOjgUtBVlGopt+G5ISY7Tg5FbGiAHzIh+BVGZMMC5CI4SVPMG
ffUqNkilvrl9dLbr2rDNpc8z2LiT86ymph3mSHVhhdBVM4tWDSIcCq2H2OylIKvZ
2eVn1vBpgKenga/e2TyB3d2wvZT6diHKCIBJL72zg8gsPTFb1BIEag5DKp7RfaUg
3fUVDxBISrIiFbUlVc13pt7QDCA5RqYPARwkTF+F3JptdnmsWO+WO9c6e4c0o71K
h6Urvt264sGqUIFrOUXFv6YwBuf8qpPD4j1cIY06FFDeIjjE78l1B9E60PEyjVNz
O0iSE/0ZtR/JbYvqeVWLfTUVJlRQ093GsME7ohHrYN72Tz8W1hOfSNWG1WJbiTUZ
dtn7nqEBHQbeDMUpGJzI+XQYmyjZZUxMFDbra5/Ovjy44chtB3qHBk1iEcmRzhG5
6M/B9jAn117SF6gf3zOnIsPyrwWx+D5etjrRZ64R7jpLq4iswvGdKNRo3braX/J2
ocbzfNxn8YyvtCqtC4BAypqt1hG6EU8Le3j2PHP2da/lhNeV+JUkZydRfctjodqf
hUE+y8NRtGjkLYrnG4G5ucSCTifa8wfW7inDkIzNU9Ce8D9g2nIU+73zEB7twr+G
iktSvLJcFf2sf0mQwToauO9CcF6IEiGlw5sdtqMl0JVmeQt37WvwHHOsMuaTrBv7
Hd+wsah3x2FKfvCmZgKUodtnS8CeLh5C51/cLKKdSqcjLybgjvAU3K6vlpyy/0SL
Rosr49EdgIA9Vb2toX1dZpnag6RuyXz1Xlf6pT8pKG7fy7guHAMlAZdzAACNRmRJ
dQuLXSFLeLwXxwYPz9s15ILGi2F2MogebbbNkX5kadIqKx1XC7WlB/X9f5u3pIw3
WiiyivLuPtxaEUviy9XVjFfu2jNgrOlkb/X3onjhFnWTKNDrAQG4nZkhYMMV7s+6
HRLRENXcSVp93WU1Je9MWqINk02NLoaVv3VkCcbpif4ChJrx8FwCxI6J9UqVMAfp
s1mlsCGqjoTilHAW8bShsdg9+h49UyzVZ7psVVfq5i0h9gj9sN2CU/s5cOVmqm0n
52/0jcbBqsJu56+a5y7+DAcwquPWDhYbHjYvNOt+K0l+EnWKfrGGzBygKBEgj4wh
mE8sw6raPWQZ10e4a9+9KX01pxsLj7KKYMtK/HsJ3/OJDyw0FWxa9B/dLgaf+kqa
Nx3z5vkXc9STjK0YeTFkGokYe59Kz6/pbX5w+cWh++vxp8YuZmrhBylfBJYskFd1
wroNdVSat48qtqnGxKQR3q6WB2weweePjzsOZVsADoq7EUixSGIUKRlZ+d2vXHIP
D76fbVmYKDKTYCx5lyiGmZDC7td67sJF6yc3urpZ6DBiuNBhEsGSntw9q2+opUYn
CYmhw038GV1pS1s9xrXrTWTpjzajXTLQeRa9pjll3ftbmYAhM0kbDdTBN/WiH9GN
hbJWcHOQnXNSgFXmbGG+Pi8V+L6t9SSh4cAEZtWcZzFQnhTTSurU8mc2Mm8sNRN/
ROqo702AxjW9o9RYphLr3iahr1g/yEVRJ//CVaoIpz0HHkVUYt6WHmcIXwAorl2+
h4vjULK6uGvm35e16FlDtj80H1CHDsGI7H2Mz8mES6w/lau1JLNwsidV7RhIkLbH
yAS3Vu+IM+m8WBUqGjTFQnfi2q9FGNKd+nBeIFkuPH+GikCZIFpVM0LCNhnOpYpv
hBEG7deiIHxDik7r2iWGiNPVxubhIWULwM763OnCf9EjI5fz9MwRrMNIhRbHP6ze
rkRKyMG27Eg7QIH5XjcBDmz/rpV4ngpfTtPx8oMkErZWBJQyiMFXeFk7dW3mbSoc
dQJodizpitleHLt6DwXLaaC9RIb+LknaxcjjBXQs4Dh/R8JXFgrdjerGA03vhiHk
9im0+6QjBie5+nCYxy2jhyEZhypmytF5tCYQ+lcev8n+yU84sr8x2dDwrAFBlu+j
TBUeDptNMqspouccwRHQePQXgK6o7Ymv3CA+o431fnPrZYZvr1olC+Ldku/n8YGz
TTjAXcgXhhcO121vqsgYBF32MbCRmhFc0Dgj9EPF+nqLF8wbZKL80HAnuemeE55O
BFOW2v5SpuObhXuWTRAHo6j/JPwr2GIdNw14ZfX+qi46eza6kjCU+itvgxCB0P9H
vfFh/EdpW2KzM3wcKQO8oV2tBZCcjKE6mNoGMF0Uo4GiCTqyBNf+YQLS+9rHlNck
7TBlLnP0tdaImJCSEB/tAMVJ/eB16vglmKBSkrD9JhRL/X5dpbB17EbjQ7FQYfCf
J7I6KGDbxP58FjFDOcYTODrIYDkuv7DJaFvuP2u0So6Jtqi/LzFPelmkm9a8UB3a
azIDrpp09HM4YB1d9ssn0QCP/UpS79ZEhsU1jtv8DjwZZDvAvSL9oupgqP9QUSCr
flzfzafCtLPMT0zE2wGN1srOIvk6VvuQLqwzcvcbLqJckRgedhMTIyKN5pBAVfBX
1DvWYAgzOQrdXBh2XPHyW2g4m8vN+hynam+trK+bjSc7gCAXF8BLKAGhKlVdXbDW
Bb3ptQKLHwUHTNOSj0Cl8Fu0Yqo6MlyPyIK7mnWtHeHQqD2YjHrMu+E7tW8VHLMV
4fXBx/ItvV3oDohBNKm0YCWH7LSIrTkBsuakmNg/WQH/Xj7tX4torllqpVUsECNt
UCFEiLEA9xD4q7rEeztite92bbD9JpYRKqmXdjKOWjhCUDbL3MXpPiPsjT5/wZhF
k+etOK5y0OPmja+x8a6E5ss9C8bd65nC5oRVrIb7NaTzneb64CUYE8LGEltJroat
lpJURIfiive2bjWy/QFHFO52Jp5iqkxvPsZFozguxqlSheb57yBAvpPIiDOb1LZb
k0j5KLWzxxi+7xq95PfoEb1Fp9UMO5vuc4vEEny1Jb6uqZkmSxWpkLZGOlFWtOCr
CznlEXQXnrdslqQwDbGYAJozq+Oh2HsBnVX9Rh+TDyKlFnPwHDAVV1xuaUSu8JWI
yYJD5lrowS+XztVvaNfBlpbc6qabvGhRdWcToJSDTt8+46CaW2n+pucDKzV4QDX6
UAluwMJdv6VW23LdEgepC4zjnBY7ennEFK9lZLyZnAOfMIZmeVTk6osDT2QNJyN4
zm3bRGrw61nA7hfRayUitlMCynm7pmy5RNVNcxt3snLLMnuqaN0x6ACMuQ6ytYwE
mlOZlvi6hLgs/aAj6n5rcPqjrwsKZiMsaVYX1C6WBqIxSFYKhew6fsc2nfOS95gK
7HQrQJXCj+mLiq7rfTAAOL5Y7A7FtSnEYThuf+asaF5VjQiIzrc/zNwPBVlP2E0S
VXQedGQ5geFvSYP8o5oCqQmZdbahPM2TMkvcSgTkfsPoSWZGjdAlP4ftZwHNsnU0
Zs7ZEngFff9xgl+aHJ5sxZG3iDpvYwcDqTLvviGY5kkVspvoZ/fkAzXtlRq+WHQQ
YVlJDdHMOjUaBnPsLXCcoXcver9mg7Nf5ZegBL/hIa++jgnmA6YbYMFMJGILRvYh
OMVU3trO/DjTT8bpXX7NlQRpH+Kc9H+rLFa0PBS5Ic9qEw3kiW2xE7lqlNKYLuXj
915kFjO67eNsJCaFGy6TagWCqIz0kH/TwyWUmpSDaO0yKhsBlyRw0u5knXG7B6OR
365V3nRCfWe54QY/dQsFCKRZS6pIVaXLVzogd8AXGRtjAYPVyTJ526c+DVQUxuYG
QUCGJHvn12dKXFVBef7k3SHI2KtN1GkYYgSg7rultg7BtN2KSYnqVJc2NT/TPUCf
JLN4+OVvQJJN+yObjyyPBFR3txq3TKeAnUTPCaOK+Nf1TTrzdeDq+qi80X7BOnMi
ahy5/Q3UFyNlo42CthlF+T+0T8/VydopjBpVkAmNKjTTdGiWndnztyKd/tIaoKX/
JXom3L9OkvF7LZNU9BxuflCJgx2rD7bGVAsUDbBLiZd4FOD9ZkIjJoQ5a/jopohJ
5HcmqrTT4AVke7tJrBOZ2Q4NROjFXGyqLZ6TIdM3o4+2d8CU4Kiv+w969KDmv9+s
QthWJQQlwoIKNTaE3xwATvglou2szJQqz/Jj8N8rnYStfEBiMc2D2NEngHdaTrYz
Xmr2+0nm1hDmPCuZyCRvjzvASKgrjggaAffzdiG3VemLXv+8Dj/gSTTbUVI6fsoC
cpEaEnLL4AUh/GkxSjheugTpOt+GcwP1E0Q+IbyZNwvlkTT6AmiQOCkTdgXeon6M
VRpiOCIXPS2jUUOl9e46DsHgI86BIXQ5kQEScMgg+goYejH0FY43Awrfi8mucsNW
974AyLsvtcA+O49f5xdIHb/NPL2r1kxl2erJ1ayppuJjmcVSvhBudhJHraPu4VmD
66CRpq/eJP/3hfeiEzEDH76NU0JesrKmeKaHyoqBBwXBKIA1Tg4MOsHzbupQ7ayR
aH3KHYGQNB0h1uZPjv4mtxRSHcppezoTKF0h5dYiAnj0PH/Fn04wni/s8wHPX19P
mPpt4uCShpUKPS54orfj0J1Ta01RaUrxNiG0ZBXuWqvfb8bvq0LcrdeRdBtVWMRN
MOurb2SscJ9V2YQ+fVq/qDPr9BE4Z54suIm4pMLWS1JVJjRssZv5S9avRJJV2t7F
y/gbWJPA5tTZKvG8cZ86QehZ5MMr4kASkCcNg79Vxlg0tS6Gy6/Cj9nlW/xGMn40
yYB9BVtMCIf+Dvw/mJlVpO9dPXuVEVLLlNminTlPvCkTWxfJakpSYtktGes9VQps
5eFDsE3H2F1dd0ApvZV/m6HqpuCyfSef6SUL5ev7fcmaEi15V4tPfEjZuJ9RwwV/
ysbij/JcTC88YQIN8j2CLwG7EsCJtNsXOk3oLKtPDLdN9tr3zmQtW5Gk5doI+KTw
bvkkkYp7id/9/K9imDBPGxkScKCIW44bsidbZ2HIwDh1mUsS6mDJiZpsXgjCNWNI
2qNL2wEIcvwA9UcYzkIGguHMaUNvKnME/vEbKLAVaPVOJfVXy7j+oIPCYSYdIUsG
69d4xiiIiZoh9xPgrgN+59zjIF1srpWl/GGexzkfKjwk1hMbWsZYh9L3rjA4Mqup
Pph8QSvDO0P7s2YPVTWmC4JtO/yxnfP17HxCEZT+xbGtzxIAgdQRm6h28kmciiJn
xF7k2GWBJg2n55gucm+GpcX1hLMaJyuAEt/kdbMaHm0//1YmF4vy53JeN7bpG/52
U3640W9iYUENH/HAz7dkfAfRPHmhC3tIEbz3KJts1w47I4RWnFNy9cMwbZUNyTWT
z1YRL1xP8TWrTeuiHBZH52EL5ZAcoZdllTFArTCjBjvvFc04wP1dMAaYUaEGbE7E
vYgsk+bPcB88CwoG3K6od6qrXvCQLSo7/8lfr621GtbxeXVv+k1i8e+qamlKmDjA
NoT7wWN8IJy3adZ0MhgFB6CIuSefaXIp20fMvWxdE+rtUBXkQ21CIMyBH4h1O46p
CWXJEbwkqpOwJA/durv/1fXjthrlANRO4tSDdyegSeDkU6QlhOl9psAjfKsZpI0R
WYhrK6+rV96ys2dhdNZNrLm7jEbWdMDO2iZtHw3Zx793WhHM8RxINNet2TGMn35V
p4bvJHmuqBu+uONF1lyrl9Xs1wZilX6Q3U0mbwNujPKvf5tco6VlqVDI8S4llQEu
cdtKpuTbOVjnPmNFFBArpdoa40jsU8FZ5OGK7558fJo3a2G+Wc+Lz4oC6wD1sT9g
SnOgM0Z/SzFZEx9ewugWGZ64hMkoNU19tnl/CT8xKC0iDhQOSZa7wb0Hf0UchZrJ
AWtoXn2I6X325V5C0DYxoRzF55S+7+iGASirUTOrnunwzrqnHzZqpxVMTOf7WdwE
j3cvVCphqXEsAS5SuwnmUAZwqxxuym15mPZz0VpEZmQm2xZlt63yA8X8u4Lm2kHg
TxnRUIyzQEFjvMgNmyBVAsj2UWszxaIePSDTorzTWCRrk53CAUnQn4byvkyn5VWa
Oy2NpkzUnRGe8nW+3e1+vhY8u2cJqOs7hxdByzEsCAc078BYwAozvPuckF78QFo8
uUv7XnKI8D/gjiIdUaRo0pomQWUhj9bKXZD0zYRwj1uv+ntPZKdqfZQ0QwGIVQgp
WKhv1/Ac7BdWYMIyalilqaJ9+c+KD7jRkvWTSjlemR0m8uDaraFMKDq0ZC2qK9/m
W/sE6oy7isd2ql8I2YugC3KDthRa1QXOLJ1mzDmM0wnSQCTerm7KX+gnEeCnPZWH
xaHr3LqmIrM/yXXTuR0pQvrHVZOrk1igRkktuPgZTSZZa591EQQiFRR+lcpm2CFD
pWMd/gRzK7in/c3FMywUXRjvQr10nbTBVjC47SqpzvGqfFTvyn0fdE5o1NhFJpp7
ObZRdWNHnHnKgiS0ak4hsqMypux8svh82Ho1UcnPAr4XdzrGNoyjxSPJEr0W6Tgi
VGXpAE2AEDar+FaYSsRL9j8ieCGw6yK14jSH3PV/r1bya7ze6ITeKkfDtRpcTLxe
wqJ0T/xcH/Su5t28z9sLqZ6Me49SjiLseFaewHZ0RhrfsfeQAKwhzWw+25+8M4sB
QCZcfcz6ViXB++Ou38NbnMATZhAMbC1PjCmpiBJTAxouSmXiLTcPLl6EjpYNTrXJ
npEqde+FY5+zWs4zQA/ovt6iqiscA3ITZ8JNcqTRb7Chv/vYsCFuyU5P/qa2q5/P
tyZ6v+VtwYsiaktCSTH68WlacY/8SpXFr85tafoeXGqbqVYXx3XXL3g6ggB/zFaB
FkutcDN95XLxC4WkaCzXim5cfMdNyBRwBlRi4I6StsAZRuY+HlnzoPRbLwSv6bv8
Nmxc+PR8r/bys1B7/4PVKt0LdYz9IAugxR+3rLI7HQt1jEipBs3/CY8OzGhiSNRs
DH0IUO46Wny/oIUbXY204ZGf99CfMKzKTZ6jmJkCjSO6mqBLBlNqEePgTm8b1/HH
Z0Vs1Vc84uKLxLtDSx+S1U8IvWxW/Xd/afi3EXFrFHA5T7XzrVfNf9J3sgII5bpV
LFRpRKHcmqk6wwsH30WF1onc8gEzY613FtMUTlo5sPpmK5EXSg4FX/YJnG/WmMVF
Dk8B08WdH2eQtXSCfvLkA0B/xU7WssJpye5MadVDoa5ln2z5ZvTlfraKkOHcxVS4
V2Y2y3I6P9E9madFxwnXOBXJW0qWN/SqOQKrlIHxzddoQ5XzLipfnAQRoBwtNnc6
/cZS/WqyFeTODfahkJzynGQRl1FqixK8J9X959Nu8WX1g6ClHONWkbHLHTXUm3uI
CzGvVR+L0FDJziYHmGajnyBVudh70nVJ+ixJiJd1kqLZcJ2zW0ocEo/z2NE/a20Z
vzSamd2aNOXRFyVJvYkRsjui+JWQSH7A7oEb03cuxsDM6FrktpcnNpzigDXwwkHH
wsUaprSC3mHRyBqlZei06uPkgsIMErCrudpkcrpmk36LftOnsUMiMF5tSPmTduJQ
xGmcsT4EJPmnhM3Zz6H69uSBocJjl0cK3YMf+YqlEWQUKsfNB5YAo3dvfqXnPH9W
eB44GvL0nUHwL1s5A6iyMexYTEP6p1OnMWqq9b1z4OtF3Mqxmw+7prcupyODltBV
yWQtXV75QSRc5WRretVMrQ0D4mclaPtoqC6R+r10LJRnw8nT4yr6kUp10Uscg/2B
herLKEjL+m0ChqaieCI7reT5Etf22vjdDIawk3kusPo27vV84mBrb/CyXjUgDTSC
myJsJlP0OKr6QfdBkXdAhQh+e2WvE3GePdXsXs5j3jXX0l3KaBQ2ZHlln5H9zZfn
WrruZl+RHoKQNNYxaAaHS7l0YXiDDjWEvHmpjfYeEIxgk4N7O49Bt9ZlbzO4DASd
rd12tjFSAzVQE3MOp1F95AT6DNuCcF3VvgWFqgem6ZIAb0TxSsdYDmVlzU/7fzEr
LTl3qvdMLTPHYsKInS/l3w6RcS/Fg7LQv/f0QmoRTfFfcDiLYFe+qmdtFNPaba+J
Y+dHQxyoYwyXU6iZajEnD6jynTX67QtgmXjeDSD+5sSdJv10w63y4QoOqMNYVthz
mGHjkENCUNAfB9KNcspq4cRUZc+idiENjiBIxlT8jTcc25uymjy1xvwfFmKEUxnd
QEalLVF+3yV26mWQVRBlpJ6OZsfSEWxgPhBN7nVAUvjqvugWY3h1BAzKWqYPBPJS
LIx+ROllSv+d6Kd10Y00ouNk0oqaCjV8bCfSIAsr7qZWpK0oolV89tWuA5krShF8
OQPYQ94oGb5XTDVInSOuFrMR3r8vAj+zvlf47AkcOhdJFlqxLkuuP9dcLw6iZw8R
vps3NrKyUP+Lz69GlEXRbh9dKGlHSSaQsW/GXpDnAdyptH04Mv2uR5TqbURg97B7
dQFXRxLaEBl8lFgLKT3f3Bb+IJXcVmEzewJepaN1GRqOBbiMQa/tD/AM/OsfXHgx
N1sdWGA/x/eYF/8bTxtwn6o+T8XEhInKyczzVtFcSfFMFjN5T8FsxrrrtvrzE7s7
bSvw5vQP2GI9HBjTGU3qhumxrug6SRutW0mvHzH1bydIZRdHGy8l+JwVLdkOkW9U
PKe4QNWFRsdTqzKjrQjNVIeEhCo+d3NQdOplZZ6J2PaFkvoAbigiLV4nYq62BQpw
0VlXxg4XaycIhL/4KSf293oDbUXVhtX3DPuH7c/4bgY2x13xWBJVxQcx1FfM1AEe
cbrqT5SXd9emzRbZYMUira1NUjzdjPtAc9KHYP3GR7xMd6jh3IPj4+O0KD9bCG0c
MrcAxM9Z9cpQPmrkbbrneyC3gzqAX41wc+uH3O5LVJLt94TMMi3YtVUlPbunFAE9
ciLyC7lfdmY9qkFgHHvA/WvWTFsOTs1zVwSCXyI3SWwoIF2Bbpj2Ooz2ehncKRnk
whBDABic/BdH0wur6LdeQ8HpcIjpO3biOh1LwD6NqZiaXjM5HUGvNrD8Zmw4cRqk
3/voKfvbK9aTfU/1itftgel61XFdWFCz1y2VibTPvhG6Z/yoSJGkalkOXiuVlz+F
zEgrpjqmCcLOPettCaFYctb2TNol9b7PSjDBx8yyne5R1TnBWzJIvLKE1JmV5vn0
/D2NYTkV8YNbM9RIL+gPq4LL73Su9HN2HrS0B03VArFuvsCGSDl/Qn7wUfdjkwpA
xUSYdHdzgXBSBM+Dc3rxxCfIB7uxJhRMkOF9q6DTDhMMhHSeWt6sKZfN7fhyhCVp
hTriPDqYh2wtZhD6CGxX6cdkSwkvS0ShMY2nY2ObQSt0pq/Uh0OmE0WE0qNpUrZ3
osT+hV+4+3xCC54jxCSmAS3BtNAgJkEcJloou678YgXPMRGUfm9qf1gM9sUZ54iZ
OVH82R6dVHAK80vJu8RTmeG9elPqw3LXvDoKdB6oAX8HIXzpWsaMnS/NSI1FI/sY
ndcZjFNBGTX/rDwbISl8uqomcauTZofNKhukTUUEL7BTcn/0t9U4LccXPisE5Ryc
muqfctWCi7Y5VselX0NOzHavWugu63T3knk97kEbxLkTdbm2tyft/mC8X402bb79
QX7w/NVuXrUWAb/ad40Lyc/0u0sdMWDrJycy5BdzLA1NgbL9O/WidUAs/nMBO1C9
Ox0CT/el4t1Yz5WgQELamBgm/deV6ewnROsI8NT0GnQZ8SDtOBp23r9bUtJ++wi2
b2LE+/ZX5EpyKwXP8pZl3PmawTLmoHZwwMXhULgOkIIL0LoRm6RMK6mjiivUXuu1
VtNlaur+j6VXspm2dbcD528slYavisoAzfvS1qp7dhiv6eIupgBwOwkuf99kYjLO
GpXADAEFqg7HUM1ULfI3CJDqnm3MJNzNbhHrsWcFCJikLBOAJehP9fXFWTT5a14s
ilb9cjL7DKpeK5Zb9fTZcAM5BschKYjpJn8UGsdmZjDQcEu9tA1muhVDWjNxtGDL
acoT3i/4gyprc2a5L5hJSLq/JkaXChrYRrMjFYhMwZrTQb0mUkbE/se8oALNkGYL
QpRDsy+DtM02EoH5mLGAelOug1IfitGJmBN50mFJVfhQqT7Y/RCuL9vTXUbuc1kK
7Gq1MpZqp8w6an/t4jiNRuH28IFvVlBzY96emkM0oIOPReaUDKtOFrZqtxzgvuhu
I1qY6O45jlus3A/0XuTlDhLf0dq8756H9tgYg51oeOqXypYp14MtxBcTh4KRvH2Z
C5Pl526rAR2XIldcdN8wtVDw/Nz40YZ8zKZAm7Oe2s48fdyRCYACGqAKZi+6RDlu
twziFpZwjpnjWfwKCpOCnAfkgvECzONfZbAZvh9ys7HxlEk5NKDbNN5ejXVzMDZR
h+uRRsZFCBSzjFTU0srK0nz1lXV8DeBspEzPCnPr9ARWUCgnHdecg9h9HnJk1O+D
3SWNela1iNEaN7IAw1kSYIM5mvNb+4FL8P2rdCCLQPW6bRvqbv8sgHotREhd516L
QSGpsyEVgh1mbjwZhCGPxJnqupi3Li1xP8TbSLiIilQ6+FA6sfosDgXiBKpoKMoL
K94EpOhSiPdoWuv5lQlzKtAz2okycD2WnwoYJOXOs9ACQEJGNiseQ875zqRbojU9
okvRYH9AMBC8yqxtFVtYVtUa7X578ZA7o6uYC2/UU5Bl+GjPDiRYVdZDyKk9znZS
rBbQacKzSFf99+uu6sC7RvBtnH2FlAAUwfNzN1bw0D9gZ2zNgo9i35VARUNbdXor
Zz0I/Q8sgE6Fvam9nbdseUXKvKZY7DB5IwHfEHPCduxi8jJG9BQdi8kWJBNHqjVX
xP0jtmttY3y/BrcLuHrKIhsRokrcD08lz0PH0JhhASrAPO1r2Y6kGRwLjvnnkimT
EUOHEO7fc/WKr6Ioc1XULuGELcu4Tdt44DG80XqlUqu9FWXhPoENSzdjx1I0OJFk
tIprbYqYqcYrQ8gkCZlX1OiMbxjiNOFbmZM1Q8EIFHzD1Ewuh9HWJyrNwkWb30HG
ZPFoUwWvxl+l0Wqh4o8SFVn/1cTgRy4jalCxhxKzrymXJraC5KHGMl27QkCoTUBX
j08JD4wvmFaFn9G2XOpElIboCIq9o2CGsJriBUl86yfrtPNV5b7LiuDzDBRj9tpS
Ooh/9+Ne/yaWs8X0bcWbYBudQ50TdRo8+mnwVjo15HlnBAD+Yv6rv5JXAI4VaNMF
FI08DxABuRKawL46Kk2wGrAleHLjRu1KjtowNWBNiVlYi70osEUqSoqru73wvIp0
lvWwtXtNUedPIghIr/QvmUOW2jhzhyhA03liKThVJ07z8I9PWHAGnPSSVzgon2Kh
gK0BJYpelTy99kI9qK67J8/3bwFxDsNbJHyoiP2Oe5R2hgjDPzgjIbxKiv071xp8
MIN7fTaNoG/iG26UD/dLoHtl7VQvW4GHz3Ia0zzPbu+F0BNKDf9BPTBhHPUAXt2O
rGjM/gEHLrAwWWveppYUFuJSq2hxbEqcnkL9/DE0lyudtTs1sQQqH1E+brf8+mkg
OrRIHljMyfoJ5gPsNVJqlfChnISRtf7rDNiHHBQdG9yxFG9ILBD8KW6WJ4u4fizc
HzidAekYYaA0R4dVT6fVmfkGNcrmZhWSzmR0I76Bbprkel2pG2qqyWejUADtD760
xZ9W1FSj81gAKFlYZZLOS3E3U4oy8PvN7880q8jPWOaCm/4UxhnlhX+2ydTzmLy1
V77EJPdlrIahEnqTZMIUpWv06BZQNDBd8L9wMj9nMS2JPN9BFPmHwJH4wazXkSSf
qFF1Kt68Z5NBpqW4M9q1nigkUK9pEHznt5eqI6DAa9gIewJ+fxrboEYNdfGF4k6T
NJqzn1Zwob30iGihavwM3YwKvBMCafclOjI5fY7lgH/kZrxGgQ198+Q7Qyi6GiVN
pgAzevhK4pCnlcFe9yck3cwbCL6J+Pxrn6aWmO9N4d6IRcQrnd0NNtMhFj4WmJl8
rA4svlyBRZvApR6unhdGqygfBs7gD1v/xydhZwX5q5LQqng3kzvtvQ3r1ek/TXov
wVPyvlfr7PbCWN8zycySNoy1VsDZ03LrlXhToyQPMNJ6E0fV/1mwwJVbHCHmiiqJ
r0pgPsrKLXdRn68iOEVX6qXsc/+giM5fpNEUsQsx2z8yJ74nKriMquJEjG53fTTM
WNZR6BwxnDujm42alGxPpGDAoqbp/mfsZxV+D/v8fHoJ7UlBgq/Uh0kCCtA6UcHj
7bo+4ba4xPXmY224lp0IaW187kyyri8Pngq5LptM7Mu4AzytsJKomt0+hy68QvJX
soi6y4hgSTj845L5btlqX+d7sq7VfR7zP3dL4+ovo1SFW7lJqc0S0I8P+QzP0kD+
rYHfyqWhx1U/qy9qWs/EAShghBCx5vS/X+gamzozEVdYvM50qZ3YOytr8moopAUv
JwsNIl2EjCp+KpHYEnfisXrwiKomreyRlQ+TuzXhIl9LTmjYhccbEm3dnr1FIu8v
kRtm+xsw0y1yMWh8i8KEgUuTkKkGz3ZaXfn+QMP2tGoUVNlsUOCsGNFJhXLdKNWW
ZWYEf7KhgtEOUXUx6hHfeq7rOVmKTFZmOVgAFI0Nvh+9YbhpTNkowkw5y7N24pl5
GZ3mmGZx6wLUHgOoGo0hTQo9/ZOQzyITb5TGooWEFX6tqjJgIPpYhMOT85NyS9RD
3n2uZM4OJyMwBm7L9VR+qN9onRh6q6RAbss9aLywyNPuuDsS5ywsqvme4wyNlJck
G3dAfHxDe0RBaJaXJtS0/r047hSU/gJHjf/nU9BfumJMzBymu/Jz1X1lBS/s2lny
gdIL/6X/wECGpyKDf20T8/XScesJ+2Kcu+6Zt6bwqbG0vE/c1QJVyjj0GxxhKZwE
UFddVF4pfwITgpi1MNPBBLnum3VWcb6GcLNtdO2RcawF+0lOaJp1tjJ7zzi9y96N
l5oVTZfZw8/kREPwLcSNl4JtLLQ1pb5zZjyyWklZ9B2qxkPkCSozTwND80Lzc0JF
VCiub/r/y8/va0H7r8blk7HseGyerQJ14RmlSijErNUl6sxzv+oBW5m9M5W9Bna6
tuYxqenBJsiPwWU5Yl403CgY7vIHtKp9SHkhAqbxfCidd0vOTttUKS3soB11EMjH
7L+3uTx2gdoobkAwfNOeKE8R42xDgG3lVLBoi982+hxOvbRFY7izYcw9lqA6vLKa
19Ua2m24OUEJrXSt9op5RFmdYMYb+V7h2A69l4shSaNbtIr4VKlumTArf+OFcsg0
n7yMCnmxEWnwJjAGy51gJeLV1m7L2r9/uUT7OLnXVZv2zFzIu3mLas8Vquz0KS7P
wq1E9Fr/0+DqE6GC4mwx+7VyDMCADzIxY5U4Y2LuVUp9wuy/ETXAocVnBqoAbPTe
tk+Pg1sMo6P3+e8YeO1s67+kiLNTycDMmEXlJimd0WQusa4rAaUPMZKeER7PRwRU
V43Sl4V6KxijRgAOqgA6cFrQ8em2nrf1x3UosgWrYcBDQ6iiYJdeeP4B08ut7u7o
lnbwCsH7w2pCDITPpC2g5u7++dgs31/ltzsVxi7APBXR6wLMro/bbTB3fYbyM+uW
p413J65B22IHCf6Wt5MEQw8upu0vNMyLlX2ZRhvdDthw/HuE4SacZEP0tRd9B2+v
l11gakiEDe4mn6JSX5BZd9n/Zb0iiagmJ3hUfSD6qpcIUzoQtIBpftwjgf/N01r/
+GrTydZv9dEY3oaFJrkids5kbeZX03uJLsNwS+2Zlw2ksApEANuTvggUbHuXYzTD
1zNilMx+G13OcsEyJ8us0nQxC9Ler6PiXywWVeaIMdoues9k3zTgvK34w7LTTB1K
vXlhyyDqJPn91THOLwcAi2FdDjwTrGWySr66zO7VJe/GZvBND7O9eOQL98nwKED7
J0pGyl0jKYupXUrTvTnosQ9iDkgDpzyEJjOiMefmWNtwiYqCMGOpNCYHafA3hLG7
BcYBm0m91Cn+bgEFtOlIgsVh4+G34TpfsQi72ub5ujwdEJ600tbqqyu0GmteLdfR
NNoTiUoanNmg6Z0VzdsrqJ9RDfU6sKoT12GvTxP8YUG3igPmam3Qr+fgE66HfX6z
GRm1xGmWPq17v4smN62Izupv99WEh4RG6NTOOQLi0lMNolGJd1FMUbuCW7vnPS+1
1LZQfuqhOeZuYoSEIfeLV15V8vU6A26+0l7QJe9xQ+jRWUmoqHswvfG4WVOMCNJY
2F2LVnq5WSmPMLA0wLKwoMuIs9l383nLPhawOSQwUP4ATJhsDHuI5q3casgqdfsY
SCkjV02NPtTixvx0wvAWjAg+3GS3fdabbNsQcY+45gZAOXcfNXPTJvUeQcPMlL+B
tagS0oTPNDFOWu70SXg3ovR8rqSs0gFVVPLBbXCihNTpr0vuJdTJcjwNmeQgrppM
j91Xky97XUGdrMJP6QOMBiukzVcrusnYjVD2U7gG85Na1CNo8vRShLu+GJ+v0SdS
AHWY9q5GOmY+ueDo0CmUN3txUeZc3NHz78QZRUVdcr5gsuG0x9/QYG+gDYk9Tbi7
886QFvt8BbQgC6XpMhi0DydZ8a298uNXFAWF/183T92aFpUFx/roBOA/KpiuJZTt
1U9VgHMvDFMAlMVnvFPetmC8aifuCe1Lyt6THluZlm6XxPxbeq0/0TVa9XK6I3gU
Xm2Z6q2fw2g7+K0qSbKuPVoAz6R97g0rnKZ2BfXirt2f/z9Ws4fJ4PgLVQeiP1lI
A3a4scw1pn74MBUoB7yuWF3ZdoXNPeZmwjNz6GprpijBD/xksqdJAeWsOQkcF/RM
52miYlF1CZngtMNTQkUHyTC45acgogCH1dWVxSaCVwP3TrIz8m9TrsPxxy9NYGNk
vV0pPtqqlsqBmq53RUPzUHT1dRmC0a1uCOuVawC8NXtH18+vBZX89W74R7+MJgri
4NAZEDp7PKyPpDt3vXTcFZhSDu8pC56mucXULRtzoEObuEGaU8ebXO04qOitHuDA
HoiIiDdhEkfE3aQK9sY35op/hlIvcnU8WsEum0HsRt3rFc0gqVa9rl6KzzJHDZGD
TvfcmZ29qB43J7Lw12w32tb5zDQH7wMM3Y5kpGoAaYa4WiPo1hAO7wvg60BB0k7s
zEgcxDYado0Wg+XKYYsTlXu6OX9/mn3TVbxsUngE6COjO6oOtnL9oREj81jFa0cv
eJ7mjNXB3xQdYoQIBwtiIPzuE6SU/JT6SrXmR0CuSLaDKsOe9vnO8muSyw1ClQNp
t6VzQ0Kg0DKE8Y2aAit2zWSc4qAeqPzQYo4ZZLyJE1L699EnvjjkJyVPOEYpR8Xi
R1ksh9OzTaHEGY/IKEuwMdDf+7M9L0G3y3TlMRURwE+cX2v7CQFWZVv+muzFz6IW
Q0MKMxHfT3mJ0CxOAXqV4q3XA9JScor6vUb6U8AeGg+bFVTBHGDfjTDD6p7e2tZo
6MJhx9gk2eGVY3XI5rEHy4Zjc5qMYbNHiAsoAJ+HhzXT4BgK2v1pSb2bI6DuTlAr
8Rf+W/jXL+ZmA0LNvGkt2PDZy9OrYE5NGzr47pnn3oNKKKlkm4OzhQt4OS7M+OH2
JpbqGlxE+L+JdWniGxn2jnHK7ldrMkm7w/tbefIKFMUG0sy1KkGz4uAFi62YkMFr
DUiZbkC6MDx13qzmtwkKSIyh9CHDB76y3JWqUnNG6v8GgflXMtUfZWWh21x+dNP1
Wk1eRVNdC+XzFCVhPykdL6Q2ATS9i9Gvcle3wvSAJobGhWolj8PGhRm7/HBdBhaE
kXZOglGd9+tRXWxpqOgPbRMzQMhp8GvzinPTVYAUgTujPVPaWLgD2a0fmZISOWMp
LfDfB0VxAbnohuAf+OnsJZKxgN0ClztjvGBPZ0gqkxjJcNwtEueSdUzcfhPqMBRZ
qQTZX+9cfubArfIv5vG9dME8elGt9leohw3qNdaXTSzfMQatwiFFiWQQukgjx37E
9f9VbMgoD+jDvVsUa2s8AFIRTY/8/n8T5c3xIOhKMenRf4TNt+QmwVb0Ef7RoRLw
qjEWQ/ab+eApxuIT/kIe1YZM/5Q+gB7Shtlg8ZBR7C/D/BMAsxStHhef+EglYtRc
iBASEgUVeOwVLxUspKZOjQvZJPOnMBm+0k2Xv2mukCpaGcVEpdWtoMJD0SurD8E+
WqXGXyUpyzkBODuzPrTz80GL+9TBHYRvvHFC6YI13r1TlEQ/IcwK6mFqIuNiwcoA
HOSlm7XZtgBdXHFdBvA8EN+IzGsSKZIyx/+ZKomuBSrfidQ6y1IiOTXna1ffs3Us
/FHiXT2A5Lp0Mp6QwDcqAnMkuohwoi/bHoSphxVoTVlpYqP3cxSMMQC8rXBYPZTW
CAn8v2cXJB+VHMWLYKHfDtUacTdXR5qq0h8vEpAMp4GvGI6pXcjh6y/BsOKKsaa+
lGChat5SHf7xpO0qNObOoCV2g3t6KVGZXeJ+oSLXikzeKhVtqTn8yWD1a4Uzs05e
bHHimSCgcJL45+ifSZT2Z0/rkFzh5+EMo7pYQWgfxFupuT6qTd9rzNR2wyCilzqS
TZmW4IgBPagSViGe+K2TrUegB2/hO9+1NvMdwWyyB+X1jpwTpCV+6+TYwKfCm6vu
GI0NfLhDN6OrlWAWbmHRKXOzBqg8UcsdkYass+t6eE9+/6+YJOjE98sEpZigwPZA
7CTb+YAO/9Zifw6MkHNjtpFkiczKv0qwp5MMTG0T6BaLFT5PMYcm5vG6HdK/CdZV
syq8pPJJpkcNa5nzwyIpP1X3Pqza7r1jcMgIxAEuW6vn9/pSZpP/ID0w/gfUUJnn
WfPd+1wtxuy2XxVkSwpjR3ayrBFn/89t7/74HNKFCrvNTjxNDlUgzOeMQf85VdE8
MLRFm7UbENu4LHX1SjMwBK4NglfTuG79nDShD+6ZINepuy641UKtqwJbPyuMte9+
Ma3aaP9tfXog+wzO9NcpajG+P4x/RZvJk+wY49AvQUyRxc8v785sbjH2ELPJdC6F
ushJ9SkSX8FbPQbA5AkvUbRA1tADblRgT3C3eoAndGNHFnuph/gygQbWqUPm0n7M
dS7gXDVDyMQjgKZ9jatFLLMAED8/JrR1Mh7WNhR9/80YIWdIZU6sT53gjXk4CUN7
fUkKtu2/eR5/UtMC22OMmNVEmAjXPP6FzSNOaDv2Q+o6myesgK77EQnfyxTaQZsb
E1dfWJZEw0if6jMGJV9z4dVd2hX0h7FRyaTAKkgdlz0LQo70e2wii0A1n4rtgGtN
7UbJcN03nGRwG0D7PVqmXDw361UOW8k3AoShySIFpluE6YkulqRli6psOc4SJY0U
Qc773wwX89MWdrlzDcyS9PYo1gkAMV6L8s3UC//r9T1+kWDvjhqsGfft11D+YXG1
lHNJFg78H9/j/Bx5r5UijNqyBrbX7MCgsFFo32GY9v73GzUXu46/BMNQ8aoosPtB
jAWrsazV22HiuWOekkR9QoBBusqL4mGEmhvepu/0iWAL8/uUyVqlR49IQ7CP3mOj
dJ7Gjms1H7QqqD4ifHk/wxm47fRqnpM+X0x9kh+h/GGpyEaOEccYTX393RxLG/Vc
mwNSMrW2gmrCQujoxzBh/cB2SujLBa7eT05CIm8AfbDJY6Q8hf44aEadlvj6m6dp
NfkyAX1kyUVoRZ0nJScVrdzfHl8td3PW6LhBuw3h0TH0z5JIwU8C7hsN5cA6pgzt
a+1YUkubnI4i0QLxYWIQZnvTZCpu3cwd9KKFlGmaFGRquwqC7MG9fmIs70gfb5Gz
AUZHkfeLbeLFezNM6uRHMCufAot45+F+v7i/p0HqMcoPcU8j+E3jyS4+CG+AJKbU
DmH/SThZXzPcglhbSiBWRTG8T+44SfmNv7prZd7dcmlI/+NCGLyw4FTDUS+deYpv
LvvD3vJRGZouhojrQGxBDn2YkHb9vW0tqjDAPPkg8QWiRAd9oSuGx6X6DTbuBAiM
yi3UqNrHVTtZmmghyRIchW/OUNNSBWRVkizRDdqXl9uCb+BKdWVKCHY87USI7l0t
8T/PERs1Exd+nX4VSuYezAbymQ169YRj+P6lCGPwxziT3wggUSOO2OI32kc6maIk
qoP6HXwx/XlnVZI6y1uZUvLj/r6fJCZeAR7JWSIph4M4zFjM2lwUurX92ZdJZpKU
3bD0mzZdY7k5y0mDL0JHFt8zPpHooKd+5dr6Pl3bcjN7tg5qj3i0Y+jPBgPVAGoh
u1nDc/iueQy8BQzNNEZgwqmiDuHwBw+7GaSyQNoIuU9EaGZiCSLmOx6fPH1QPtx+
fLJI5cLB9Cwk1t5OFI4n7H+h7HNe19erH/iSkH50mi77oP3DKRa2TfrC1sPCiKAf
FRQZAguJSm0xtADS5PfKY+h1ONlYpRx/SbP4sUtE6RRp1GQAzu+LN3x/9+wMZKOQ
sUPqQlLiMhfOU7U9A0HNcxw4fIn2JfByYCvhY0UnqFf4kwFbsd7lEWnVicxCgWrt
L2gjp9HllYJGMSkCuI2H8el5exaGfTZulQcEjIP48B9OjDmP6tGm7hnBNT8Zugsp
UlF9C/f1rEGkOvi58lXln332sWAMEsSMVcw42EJ3LvX7OtXgaGY5ycdhAaj0/qSW
ay1eupaS6sIHER0zRoEREnk1Bx9O5vFVFIcH8Ya31jNAuHzEh8KjPv4e+u9RX206
NdHLMCoqdFFaqstZwEcnH9RzDw/1CpaDxcKuF6CaaLujXvjW8FcvA5TtQOfi3xvP
P5SaH1jINLeYuvTj6n1BJ2R2hdDJ9gvHX3UXGB9NXUqZWzieVWVoG53VOBLD51fn
ZaHEpb8+qMPh73lb99V6CahFzrU5gfGv+VHg+D+wkGKGIQrQowdw+RxvE0g803Rw
28uRhe1ZDxTFMbQ9vXlC/W5wTgR8KSxzFy3yvpCPWYc5JLugYxHfapAoo4Ye2UPx
u9EYyUI2ubLy8f6JR2mXfNosI/rSicWoActs9MjxX3Vr4jKCAb/dhq9Ng/xj8ePT
Ufzu0wM0sPvG6qIC0Yg0XaHtJlz8BdIifMc+LH4GKKmMbkK6iMxN9syGkWdlR0ml
SOpnuovRzxI+1snIN72U+ViV4AcZ9KbWMkF/yQV/1VKR3hUGEw17U+Hx0MiLfwWF
yQ1v4igeN+ah6NqfnSZhnVDnrJuTewo9TqpgBujjKnwRBwFTC4wMZJcdyB574ViF
5oqOKHqKuRUEspo0xpEYIrtBFaTEFiS6+hrgcMY37B17IuXPXohm4Ss3nJJO8Dbw
aGDHtF5EVB17OlBRMdoUj8VvlX4wOPcTVBSomRvuMPS9SN3jSSuhvv+g20yd4uhk
hC6jkJ+Dj+HC5/hmyhJmNqyJ2aXELgC1a2o2/0YMzjRSJUFdts/9Krn+Yne/0zdw
EIQRN4aS0BqRS+DdtN0JS15tL+tkGLyfJjCeglC4tj8WyNFvOa+AFhid2gv4+7ie
L7eFscKrnF+SoS8DZU+p3WIm5LmHIgpy9uImsfd7gUEJ3fJh9bF/0S5pHi3cjuEm
81v8qkbjrDxQv46IKZHnGw2Kql8RJgotcYMN1Wb3splDQy4hYqmY3fjaoq66k0hi
otrg+renmogRYKSwGZkyJHSjyjMxGRaCLRVciaq/QYt0OpMbND33HAm9Hnn+HVFr
HEXZ9ATQVG1i85kydH1PY/5SUmtlwE+p7h0X1mCHhyOk9bGTo3owXPnX9FI8RPFW
9UW4ZJj8OSXJEI+Vz6eSh44YGi1pCItsUOjQJuWzdIbEiUvWrY0szuBCRzcD1KIE
6KT7PEEOYR0iwOjAG2U8xsnA2vgp706N4X7OaIfUXddtnZ6umBjKKZvOMotnG32S
9jmMgeLoOzGcJjcrUe9slhd8Y0HqngMAch/nWzSCInQiY58Tzn9B4XeLNwJj0YKB
8wVPGqeYUkyEzryeekSw11kswYHoQAGoMtRQDSTxc1LjSTnGH4BCfNoOZrnd8KXs
V+PA8zZdVTbN0pMPzRn6P7l+YkcZtvS3gRsICduGsKwEh2roi2e42LMvF3R62X9X
LhCDv9KvrcBlb7iOWMaEAjAet6kjyx//FUi53nlSKjcrUQjKQteYj5JliLOvjIlj
WqkKzDP9csuHpe0MOLAeKxnrdraWeioA5Rtix297UZPiwRCQ3Eptzy90VDbIyHH4
letZH8B/LVz3ZODsieJ4Mz+COojnHDTWAk6SeyhTpjIkrRBL7febFhsbSFYqXcFJ
CGCW8I7eqllkjWxhqarAkEeMsjbHMVKHD5P9dDB3Jijw01qoaAOc+7mx4HVZUuzs
er9iX9zlcWPt7fxdW9n78LLZFb8kucpsOpnnjoN9Mswng1jU6LG3jImiG53iIz9d
ZoRBLLCWIn6F4kCC1ztOwipw8pYxdYlrLLI2gbeTiHBtiz9wCytPXCb4kPWuo3/d
TEnqmAfNYo+TufioYbNHgP5GPpShJrTLfO3CKx+JFfqQVqrVDqBq7kLu0VNNV611
PlaiIkccVwysBGhywVoqOji+JF/aLXlxZOOzExNzWI4oMl5s0MnR9VOrSv/CkPC6
OrZY2wklASE6AJcvxismrmTqRtKzLqQBBDSAcT0ShgQK58g7XGeQ/xFzU7ek7sdP
sPtqmM1AJsI7CxSX1ndmjTggwbAzuZ/jrzPwnS5vrutPNvrXngmtX3Vbw9UHLLRJ
PMH04/8oBw+kxyF/HqB0sUIVxHg29C4g4kWL9J+ecwOSDjF76UbXU2Bddb8Vduo/
CM2aKBZhf9+YDqpEWR9fJlrqMEDph8oyKW9EOpfjI7tojQTHuYmuWsdgLtgpf2vR
BcIEdn5gprOsSXRRCvR74cCjxcg+urRGLky4uuhn9Ke/t50M8MBHabhM/Uq+1WBW
MOa6cYmB6GOzLb7LHpk10A6PS8nFsppEZunnQU1VCG/UHcxhnu9FUG+XOs8mpiyK
DGlTM1eKt9g71c5UgG14i5nHVBWZfccUkUrLB43CemD+x6mvgzV5AAveNrWoXBcz
Jp+Ifly4XlquQXNMNm26OPRqO0tMEwu8Kf8dmWSAbid7SDdUr+Dn3rUKd8U6tel4
c2uyD1Lb39ueIeQpWDNdx1YXXTXwtyZZ5tb+8LtuFXVVh7AVxffCpHKJaR1lSrTy
NlLSaI7MtPhqYzWemro60sSdW1GlMzByuYnrfBq4DLoTc/AGrcZIhQUMOR0ujD4b
BwBZtirumShYTWrSD6TN5UAc6p1uJ+Tqg+oNlTerUOKLXwyu2dqbHKOLUdcBpnn/
ZizJ3FKMo4Xc7f83q8n3nGJ5Mhdd7tGLiXFOyTWh2rw0fI7Ggnki8QwG6HaEttJL
M5qtR4LbX2uxA4E5uT3o0ZmrRVW/MmSb9na8klq5JWm8SPnkhw64khrmj6XnRf98
1PK2LcKyUmrA7qkf/DP81mwFWDedpK6qwXGmRhZmpvVzkuhvjVatxfaA7KDM+MN/
G6v6XnPkna5ssl7JS2kys575RmcUljOzrn1dFxk3vOjSV7uUd0/W3OJBjvjg+Tqc
of0ZoeOE0usGNKXAizybT8A0NdXez8CikzzY8YY/GbztxLAHRrUFG9Rq9Ha0a0cy
XAZ+lJzxFX+CU5zs1J4LG8+keBRuM6hXCz76Z93MGNLQfpGcZGT7fT8U77YjJCiW
+2uJ7Ha1lJoUZ1LxB+sSpho5RB7B7jSd8AWqTTOCnzLDbasCVr5gd1G3Ebnzkg9i
lMvnuIZo1dnRNe6hK2upP1mR4/B7T2Lcnqlz/U2ux0T+ZMNz1noCXlh6MoC0y3lo
/QCiL1O/peGaQ6MY0hbJRhyjK27h707ppAvpPlVv1LagBQf3tUEZz3lw8fzXj7EP
1+0Z/YX3/hIDQY0HNRtccSX19Y1l4hcgE1sD0u4kvK3vcZTD6vqCOAFLTplcpGf8
BDyW4yt0U/SlldkbYkKJdkDyXqgbYKqc562I13vez6MVaavQ5Sgwz1moYpU1QfZj
xcvTJIs2Z/vNxqMFaPTRa54z61o9Vq35tmUSOfM1Yo+mLS21otKnxykFLtQisKcS
yvQ6gqWCkBZQFZT2dSIphr+Yye7BHp5wWii1U6oyg6DI2KuVXLz319igJJJYrWjN
yrxnOTRNFmA8WUeLPyDGPqX9h6H+CfSMN7TAnzvWtoXQM5SFkLtNJx7ZtmMkr0tw
79stdzmBKQM4BMotlnd4rhK/RRI7jDvswAlGq2/VPr53T4KlVxOxiNHiDBckNLUa
THpK/uKMjc9gNGSSi7SIdEZrbZ3NnRjNT1LblQA28nNP3ebHCp8Bm0oHeLzIczEW
cLeN+quNDxqgPyLNOlIlP4T6xe4/XDcnZgDrwOiafBe9ozCm2dIqRl8f32e1Mh4k
21bPGQXr7HIobVXzgfjYHGc5snu7v4PCWV1xrsXdw8L9DdQFpHkGdP7IGuJ8sxDM
SYuSr1ey8pZbODOtvALDgQp+XI3grdcBXHRKkBc7To9Fb/lnmoT7omxR/2d6C1eC
sW6ktKeZvC4u3VnctPEQVr148VgKegKoa9LO9Aai6fqCwtjMQ7CdR3tzWeQ9W/4q
ddbbri9od4gUyfYTffkgy5uzPoHI/W0/4MprGrkoBcr6ihKYphwno1GSIP3XAwpT
fKrxmNudaRy2E9WayRdqaDt7X/5AkPTvDCTiTwJ2pJvRDlCuAct1s/bbGpOMlf0K
H8R06I6uIOAMGxGGAp08x3YXRhtxuADXQj8D2Iy5XkBqfvX06fdYjwz5jUKP8Zqd
HxyeOK6nZmwk6pV6lIO00jk97JAy64wXlExAgfpPa4/oBfDsECirAKjQYl9LmcJP
aWgTsYHh+uAOFLnBIcbkFQO//BCnVhdl2y2YHIM0kKXPcJoCwhPKHsCkOE7THlC6
uSLS3pL4dDEe5yWgBjSLiXutLd/QHQBqFFqhPaa2IdsTG6NgsAdIA+MylCv8qiNA
e4JWoZuNscssHq/Kr+NoVtctvM0NcaAwrVNUIX7nWTfZQgDVNSkeHYkbxCAIeHmF
+NaNZ/SQRL3S1IY8G+Ubcgahj0wIl6yIr/TSlskBBLQEKPHPeSuSZqvMybd4fm1M
wL8XEP8JlEtogtcj9GFvvpwgWshf6sazBYiMr4di+q/6Fm1uiJm0HUHI35tNNA7q
uYxlqNmE9d+E2LadiqYAivPon5xXFoqBQEPZIQgPJPiULQAcIEeBAToL2g7ftJA7
LDGIoL9CqibajRgCBwiZ9v/umk4rcQjgusqrRyo7+dhmwQWOZL5IZkKwgTVBjvT+
MDzgeFMfzHQzMHOuNkp8v3k9A63l4ghRK7yj7h3tfVbZkOtsajEj/Nd3JBjHFyGu
yAltX6Tu+zj9jV/VmVq8oKjqR3bSAweHYGw99w/RlAgFs1+yQzvsfMsm10LtMBcp
UYFcHdooaetuJvAbYHjgmcY7X16za4qWaFne49xNAgA8jQ9HuGpIrmG7yBwIC1uf
BWvVPWtP11CdY5h1v66K6qQf8VZNz0nMbweFmYFfdoYu/YLTGskzEeIX4guJppXu
xAufYH2jEJKAb3iZGdlJekc5Q4kdGvWov6Ov1tdOEaopfm11afjyxJti7IiMr6Od
/WtYNl6EwJRuxJ1F6yqKdlP+j7ijrAIiJ7/bDRUebjEnLrVkz8tOdhDNVXVIvubx
bfKYADdYS1CJxyCMcvFj1UG2ROuJAvgmqFuSB1p2GsXTttV64IeGk2TmE82PY4OV
54f7/z+Ucl34xS3QK8+WovpHyXr+rSXcG/oI6vTxk75DC1PNCrZJlPhc1cOslTCx
hNSOOPf1aSwvSsP6JnRy53NjIEJHzvNAvFHrA/keiV+rfysTEjR+LSOgoFyQ9fsN
TS5RCkPVCtt/itUznqjbQa8tNIFMpjkFcNrEiu/HjiINuSzS7aR9ZxblhAONEtn/
duz8gRBT0eWorRJwpYRawZAUaGcT50xIEGDVHhtiJg28WgjYIAGFV1tG47HeHrKf
S3qQdev6oQWKgNzmFO+c5H+ZVUF4tULMay8uz2L9ZVeZNTFUXikonuMnDYHO+/8O
sKad3DAUKZWI5462ecrgmxTBBiiSNV5VW/nvcW6lCFzq6ndd/Mp+Zt7pzKJxNhKG
xVFRfjUHj6p5vAaKP+5/LkTuenBcPTaphaIH/FXw4h/XO68uq8/5ZW0MS4W/5ODN
89B+vUMPyLmZxhav26JCB6sanlTKslz8kvN37V1dy88ywYMVbpGLJ9dt2pOcOiI6
7wMh7/OH7EF+diCbbCmbbcgtSya2f0RUQ7y8XaM7fkgym2DxCRIx42DfjRaYpi2Z
ly60hkdoo/dUsn44bWIeX9KxuJPaQ2V1lmRU9PpzwWPspab1IvgIe7iKAr3kqw9x
W1TP6GEN3MbfFYGRSZ9pKP0ejXDoCqx0Faf+e/vj9tsaTS5LazHRhRX1zw/jA4Mn
QltfbLDMa1xXQ3E4XwVZE9YlRiFuNg45+zLi38/CYhGXkglHoCNwVmFHcEvMQFu+
oYzUe3l/++XyvbdFHv7HaZRLRTr+FHNnvz+cNgiQi+rWgVb9kGsPUIh62PLhJ8YK
ZXdlPZyZH7dBQNBXiW04JJI0CkD8vveOVbFmnRgSzVGM1G4HtQxcgitx44H2dyHX
vSTgeXpyqPZ9FNF5ypd+ghzy+8Q2Lt/H3A0gr8s5qv4+Dx+wffVTO+QvCu98QHAT
TP0Ujq0O1wRQGnRLw3R0sPUoJN2ueBbDoq4jz3HcMtJKbmTDDOjodg8wLcJ7+KEL
rpOl/8GJqRYE7mftswgEeBKiwBnX6OM6hqCLL1RG/4em9or3cLESe8rd6cXC+jNE
s+z3a7hQP/c2hEL7iIXNIzhin8cs+P5DrScp4yFzwXRmdfS37GbGftqLSKe/qM8Y
oa7v6IdjubxQHG2KVZJKTkWACrp2ZGZ0wLgMmhsG6x0ezJ0diTm2cU7CrIVXItmn
wfI5Gq0uG6yBb3OatPIBsTN6fLNwQUOYPzGKHbJxJRfxcLzRKae6Bl7y+vncEsiM
pOAZBD3rjtQwhSVrmlWgfUgw5A5/kswHqruz3W9AjZu0Boy40XP4F8ZnqbY2T8Tz
yJFSlDyGDUH3/vlSm58UgBD3QfN1JKr2AcIYyFVz/3Da8E15XYcNGxOjNT137bcP
vS50ATyzRjnl3VScRe8RBERxPkbmRITeMBY4lgjRKYloxse1itBXJWbO6ftt7eKF
3OtHKPUyWqvP1fdkq6axaQRy5n0ul2K0EXEuItn4h2fYDbOlzIVqZC+CjMa9/fYt
qdvxp8olUFBXtbitR+jfKCF6gIXJ/i72+KfLWGcx+3kYJw5YwE+1SuElECvCGowM
1bsKtEzLGesgSAiwHT7C10j4QqKvSQMRe6PjMYQ+x4xSLYwUKxq3m2W1WJTobV53
5XWol1H4I5IxKxAlBAVdXyHRrw7pOJskwMWqqF3NcGL/8gMRg9UPGZs1BocRZuZZ
0uK0AMImKDv3lt96nKvysNN8YWPht7g23h56JFLQ1CaIODL6byJ4FGVNOfg7H6GJ
35l5IUk6pTpZHEbALjS+tDzYKnsAPXuSoxMXmkM8WMXbO6tqvm6AiOyyqhbRj/VI
XCMwj9ujA0yqEG75r0KmdSF3l0S09PjQLfvhps0e4H+tEa31syCCF/XYcx/ITICZ
pFE/wn3hNmkFlH2FRsum3dI++9Rm1uiQXzxR4929CiPnv7rETInYci34Ut47g1pI
4npya5KvplZtzhv5pvTgoUIeTH2gA0kFSCRrIVflISCvdP5/T3eDkUVRnMioBdFf
fHJ+8ImR885Gc0s9vkhb04erkFF7VJS6jW5DIDeAdCy6mym+3KkVApgb1yGGdvqu
BU+iYtn/3Au4nvJmStUVaXcVmzGNmdC+vgfZ46jxjkQS7cbRIYGtqU4unXovkUXg
5exsB/kOSqXR6+7xSwsoiLji5vQQd7fkFC7q+IwAsQkYfC+zV4dHuQXC7QXRmOqZ
V7HYldPx3joGKdh9mt5eeVfU5oTZSJvYi1S4pStCtgiQShRMnKnOMfE1JleLvUa9
ydSWIM9EaJbKuk08buGcUMwN0kyyftBovBxRMQlSGy47JQ8hYgnXAK+i26ou45UP
TC4vMstUPonLPSTzpMPs9dlg04t1C0y+doMrVriE1xLx5L+Zwsx//Uq12Bsth75q
C0jatPQWvFODj5JnvPvQ2taXheIrwFjyexT0raqm9jShmUlSgoGFETM6sRY80Dw8
BOQxDIEhlfHxqw06kzO9+iurtWw4jXICXycKbtSyptBRBvz3Z5ZtZqqrYoukF7/f
2QwO3RhPqO2Gwtydb+RgLPPwFCGHIw0slKVTsUYelKFBzK+WlxpkeDnJlOx9S7Wf
f85VgdRGf0dNa6bRzsou/qZOk0Mz4X9S7f6VLQk1ihldHumRiYwkouaog3jz7pDG
8xv6cmX3eDvSyfl/B4EG2HepRH1hFSIihIOjGC0HbVv44NO4vGcIaxeu/L93GD41
nuqS8TQV9+x8/LmQX86B7VkOOzW7oEqAi8/lu1jmYoqUR8Qan1e4zpFyGJEWbVhW
46fHvoi5popVGcULlSnLaizNJzLqy3sEvRILMm1QVYO8pyucifk4j6ySlW47hUJV
DLzY6v1suCThWbxw3R4DILWxHYcEW7ghkF0TzXH8MMgylA3C/qTmplJmC2Yiv2nM
q2LjjWn80VBX3VTq3tBW965dy+aiylWeUmyWpZSp7D/vK7cHngWPgBSP4ESAyDJN
+CTnbrupnb3iVj4/ExfbZ5MJb7LoV7P0nnTpWD/CSUtPYCmpwduSgb7pcTprNjlC
OwAalHZcsacJwMlpPpWMVBG4f2zQtvLhg25H1+BtCfhQ5tKDkldUaY9sMwhHoTls
BOslvTXDBbG+HHghtdWUGzumWlk6t8nfh/RRV1XUxrSGZeRlbVHyprIIIFeRNfQ4
oqWk+NnUzmcXWN6FkCOQolVtN1od3mnmfqPhES2WQfX11drsaYOWj8zsxQ4j7HlW
4DecTElSJeUVmHDovXNk6tn4A0ZEW9V60ISp+3FBmoMNzaMFUx6XSbBMuRvPJQuD
uVKqE/6l53v3y3JIIPzVF7YMXAXOBx3BNIDalxl0RP94MvkzXmq2/nwuZ8Ibp+iC
duK9PEm8/6WXGJJFbTYJoG8TOA/C5EYv0eetWScdrt6gfp83POA4HPYk8g+2MZFu
kB3E0FVkeUT+oiLyQ87viosXLczlfdLZYwqXcETbmZRbUGiCFxm0FJmHlT9zTypH
UYOq1b4gs7HZNsvTAPDE792ZgdAoi0FX1D4faZFxVgwNHKzmQNv2unstE1DxcHIs
ZI9wnQ+CFOq9S8BRmPMlU8Loh5wKercLMqTpEE2hEq/FN6Cxw/l7/GGeBal+sKrv
tkYJ+S4/xAx3spS8LZpbDXhAVBmsINGeSCsG5YlLs6zBbjLr1KXobrjoie4YIJSu
Fs0CPpSe3iYLGSgg++BRXTipJBBu7WwddXDeFW5xzEqQ3H1xSSpaF+fit0McA3uA
0bGavQ+QRAbWkYjSok9ZpEdgR96BSL5lbp9BBGvxhHCgkhOSFMbbAP4iQ7qp9NNY
kgjX42HmWjy5wEe2H1Vt3pnw9MZ+EnqnPlIhVxUB/98snaSHVL1anlKuHtt/sr3c
YgVz9xHpKjoWuQhZQDn/yZATdr8tyKlP5mzY9MJ4cWLxcXJJ3v0VsNfCtbgmj10k
5utqlD+XXCcEsecyBtFNxnwSwYMDou6Besu+1w1WUqDUvgAXOsdCqHNne4Q0RtDE
0dFdxXFKetokxE5meC6qukk4FA6ZS+Gm2b34PyAkXWtZNxRCdVLdy2EQApVmUB47
NgqOMTEE6BmrFz/jZb9n21+rGOe+nDtwnkLtDKQ5RkSvu0MP3Hvil5LKp6kmIrZK
Uml6t/dN8ETdnj3w630xubzEiwMmfJnXfhbGmmhTON9uFUJBpohwtDPNlYNj4J8+
iKEBtNLalY6q3UD4gdq8oVjNfC4Yh57DpYNUJolWUeV3VbuDTl/gUGx4kFScTDWJ
uvyH85piVW888hPS+Bf6UOIL1vKHBnxNZQJniqFsU+v9z0tYA2EpYorPhP9vT+fR
r80HDNzhzY+5AP57wcYpTJKd9fi14VSiK/J2fWkD9SW4ss+Xq6HhLOPpbMhBucqL
O+DU+BgIwtAH3dhPK1bsJMJdwB1xwRGPGkkXyeScyqYSyjxJ567GRBmTYapk7N6O
b2cd0ibHN6IrqrL/WcLXdFKoxrL+IDOnQkXg82ei6TvtXpPcPuuv9MeVyMCrRPDy
Apx1UNTY17F61PYh2q/cNiIxOWK0Oy1pyBG+nc5YQzEhXugIYm5f0sS3+nDOYkr7
q5BZTEpRreTYjYGm7+CO/7JjzpetvkkniXPW7bgjvHcmCr/z/mysq3GjDjOfvXMc
gCKPAsGWX9BaOA9OXmc2/lYDmkvVkSdaFhR51uGpTrPhVnA8RN67wKT2DtAJ17ce
5Yoomu42vDyQlA9HA0HpJU22Fql1X37hyiEL8u4Ceqwh+6KqhLRP49gP+rBGhpqn
Ny1j+kTu4x5T8CkOEyooL7K+aVYVpfXBdW2szgnSPdYhFqdEhRo421y/5Vv7Ecz7
AgGKIBpQ1l6hIco9B/6KQLyx1/ESgz1wVM6ho73tcz3EVeOEVc6h8SRfjq7kL3NU
PH/mEa/2y5LLtXKZAZbIbD81bEm390hPI8fhoHQM9QjxncGs6vOG1wnmEoJtbgTz
6lT9ZtksF9JkK8PjuiHZZ7rZRmqTqnL8g6IW7uECej1KhXbhbGScWbgn1suHv27n
s3NMEXWNgAuw7Fc5bubXX3LCGYAJp50tFrx3kaRR9n5k01atfw+1qz3lrE9kAByX
shfZwdZMBsHcJs7blpxd2VnfJ8h3zVrf5MC65idBuKYzdQEsG62uWOpPaDUlD4W4
hWZkO7dN5R67YHNiHpYtriH3VjnakAfIK0x0PSuEP/RYLZrNMNffYi3cP6zSSMeE
CZlXoMtN35ou3uss8+Fqo1bk1ihiUv7hSDJccbW27irKpLXHktZK42zN9cdCaS4O
wfzoxc/aHn1FNhqzUr0Ut3S9glzk5osPsrWs3UbTc0/599FtnO6BXC9bG8YefL40
8blA6UR1zs8NXPmh4pz1lMlYqPL34pK4ZNCsjFOMJKxF6KhEIFHxmSDE4gV8MS6f
3AlZ5nM+oBCXd6woQt2CuW5B1bsyXcXRCvi+FPGdBE4AYHFEmFKHem67xtJ4x1hp
DB85ehdwXFuvqUtjOjZYMvRhAA5cbu0CAr5JB2JNK74765IrbuXOZ4fpVL5yUy5/
//JQ8zVWBRkZk5W+V9UdCoXK/Huw404txnuMQ1eTMPS9D8JTAHuN4KTGijtLNi+P
17kOzwJCA5cBHO6vpTQipfe2NKLqF0Ha4JMpvNX4lO/QOGgR2dLsyRS/AUEVygBR
QPw4+2FHETZEtPNOKLAPuX6w73q03vrygALCHa2/djxX20xisgM5bwsI4DDiSwFS
0cGUZ/JVnHqE18dtOSSvdRHDxDELvXESd9hESVIGxf7NePVvAxFz2zhS4DG9bewL
7YkqzY22htdokgJewe7ZLK58AxPRULcSoAgptzy2CrKUWFbRrFi1OGnK/ZfEeczC
aWXqxQ8Y0d/FEmePvQZpyArn/P9A8+o/yXtlZiErUsCVVogGMfQ8Hr4J59xLEq+4
azGyFOnISyO2/wQa3b1cbomdWlNXRliAPp3k7XYTBe5Mnv0/nF0yYt31oJyShWCG
NzBf0tQ5bu6lCdKfDgAMoQNqIZcsqbW5liFRY9rBkKy3PYOVXq/KvdmTk+E+VkMi
OICmFjhgUTSP9AX06FB8gKP2GdBDO0n+APcxy5x5DBMJmKngfk3NoCPWuaWb2EO9
yq5rHkOTCVf86ihTQAox8JFVNBod6SPDYsyiyzJEdrqpuLA/659sYDz1LLYuZxm0
93MntabJEPBWHWszOT3AXn4twhdAUq8XttdwjIAuR4j9DlyogxZ+o2zNAOFfw+tn
Qq2GcdnXDJEVjnZ9z+h49SjmERnu7lzM6c+7ZDnVImfoX4/JWXNuO/2Kk3lWmigK
FhC3iRtTQrssdrzFZibgE2zRvZvzGo3zKoeq8bV8yChCteItchbYd+TvkjjypJbx
WZ3mIgw4tK/GNUpy8EF7Xa9e4sdgUhZdmMYUnkPC1xZk3Ei31hhhQy6CSSCWq98R
M+4YPm3M8XoT2IB8gLGdIZVVrjuMqyLdupjUa0c96d0EOZOPa58ZFbkBCUa5QKsg
YMfYA63Q+8EPl+g9hVvSS2ZQLEQX67aSrDL09+NtiINScMMBwOXsEWWhgS2sEPaT
PVfqbv80tnqzb6QGdaLFOFrmpN19XtxB3f3jVYAIvOm1nNb29HF6LTNomH7L05Yo
ZNArXtO4LGxoufYdnvyxJkOF5J66uiQMSIXlikufYr9be7jL0qCtCMH4DrAsM3T7
/OvA9HIpK/m/c9Wu6wsVoAJWTzAlCI4dU5pvnWVYSkMwSEIyQrICEOacCSzWJdXp
VuiCx76fT8TYGeEfKgGK4nmxPhqV2UJNgnzsFTJ2isyuyKL04aOn3u0nQOsTotsU
ZWbCWsjv3FCzHY1FzoJNIwIdjXh+KGca/oaDQJ0Ia00WaccCYDiHLdo2It1J24iS
2qW9PApdGpyqlAojPn2HxwFom5hWFlVc4Y/VT9LFObZHKbXQUI2ebN42KsVah7dF
8Lpn1CBSmJ1kIf8Ewm9Lk5aq82HTNjfVNxJPlHjlHsu0p4KKyhdu8Yf/hCmqQ2Cj
OwZ1Zt0VHV72y0cv3zR9Mbt+400aminrSEzgXxm3UDVJikZH3mPOQZpCM/3YJ4zl
kcXII+eDW2yabE2ULsHETVeScKajPECeYzBpoZ65SQPcqpBznZdmnDnVQy3mrabl
7NWIwzhNUQqZOyiOrdfPtr3i6BCwrm6vfTNBWrv2BVx6OUhYX1j+Sht6pOTeKIN3
AwjmcQIBuFAf6AEfVp/NWMKzzJ+EqPY89lRVeXjFQs+Lod8n3b5tMm6WYvuWVICT
9BqLpxg/fOCUrneJWWGdpkx/P1BIIiP4jCJlA3S5HmL0o6+pGY764zY5nCs0gAhC
fCnBQl21uqfmbanCbsZccr2AvscvWwENL9EWJDgVSiGncQUtS85Dzi4eN/Q+azbf
speXOsmgTaCmPhjryU8Z+BRi/o23DflGLOZ2gBguiM+mKDSirs2oeU5R2iTSgrVH
VK3+Qy6R7FvrnaygjrD34DV4Y42ccvpTbCyA4dd7kUSE3tkRUvEoEyeCCx+c457B
q3m5yMqSHFHyXcPZIPKgNKaukWGBV/sXrVQCfLOataHa6BFvQf9DIyWm90q/Zm7s
B4R2ETSS8eT2Ql/RhhYVOCSGvtkanyMWlu036FO7st+/Sf4DPLmXSnXnpwak/9WU
nqgiojEZXEF07GLglfBiK42279KIcudMVlSqb1rpvRkNOQ81LNezGsHPoENtiya4
2W19UJ7VCK4YYHfkcbYti70r/rAEyr0ox1JB52L/prg4Nb16cfmVi/t9CaziuWUl
jezaBLWqUYRJvZOCnITDAS296AkM7lEPQjMHSzFlWYS+vPvE8HSe8phtFnKwNYmn
uIRNGsUXhs14aIzdgBTOGobzeUTUKut6dFwX96WWOc2zSw8F8nN7GsULg+kZ6OlG
JdT832Xs3bOOzbm0Q1d86VOjFLqCf6pfkXSiBHMdRUarbJ+bB2j0yJITor7j5jkL
HuNBxvRBhQmm7qZg4+vCcZ0k4BdFDF/Kq15q3rhYGtvWTxrnxuO40qFSxHNRNbkg
ESMrHuPHxFWUcrYaut/al2LTJFKE+GaclUIFGaHMh3QfpYpEkV7sE/cLLNHG3orN
c2VM3idcc0qa+j51cs16jzuXodYT17ENI5+HBu/67u6ziuhjiMHda+1T5ehXZOUs
LysNA1r/71DSjMVYAl4b4Wy3UHScIFkbQXPBO3VGvu9OKYT26qO18S9Iim1ROAe9
OeEC27aL8BmCakoAK6bPPBPtdX9JroJ3x7fK5+FKos6AHGHZPI/dR/6v3It03IKa
exRhPGGexTH0Sp6JMq+XGjKzpviRCKwhr5Cy5yzq+BRAXH9gGAoksRp0+m0jbrFh
/n5xU+FU3ZbZRJPNYZqx11vRSTbSFuQj/7Hjvgz4Ehb5vxB/uuegXFX6YnUzc9tD
Cd+V3QksmAGX7CxACmp5LuEaaYtzpbHs3O3bNRjt+Qb4ns3TEyLIK++BRozMG/B4
6GdL3GERfE7PxnU3D3kGsv2F4r5xqLHJzb+BJ9zubs7EhofYrHCSIrSt7/MHXvCY
Sj/CY6oTc3yu/tvZSrA+VfwPRj3jr9zrpFfiq7sY3ne0r2pVGa4FSqOBsKz4GEZw
GmoOHGS1IKlp26Zoh4STgMwpT8tDEjdJJbtexPqqDKeT5FoT0cL8Pf3opT+wH4pB
akyQUx+CMUx0Xzlc7fVMamPC1xKOH1S4JHeJ3c0pGTnfxB4gPL4ev7yL4y4BXjJ4
R2C+pSKmyapl71FQguO+8pbLYVjITHUM7rxjMVTlVYWqGdcZrjKiqUWuiCcvV2en
//2OS7PI/FLuVd4zYnIl5CJBcQddzJVcd4Cxq25TWGzedalDXbuhoHFiXli8m1EN
g4Q4ZfyrNYnbKbui52/I/Tjg4PboY6XUeY3vdnJj0itKk7xCufeZYq3oobYHDsYE
dXYKg4kMa0bqc+9k4SYaw7RO+g2vdwkhMD5jPZo7AzNhvkeUkP99SvqT8vcY8JuT
Lpq+lK74ikmG1fVZHcAoJIkPmsdsuCqzsJgfGexJH1p3g7MCvQ6ws5dYLQxnzpS+
CgxaRg7vWaLvhUf6O5xZeChQIwEOXPR72ssXJgKURhmGyYw4mBhfIMSSL/OCbfCP
KszXA8mBnfRtfZg3PEmkh+TJWDNG7Fp2LNCJjtwv/LAjXSz21jCsZJ/HOj1GTEij
Ug0O+KgOrD/y4cudUr+J8ldn6+jGV/lAKwMZO5DYJtgb7tCRtbcv40SHIuIvJSj7
4DtCjtjPQMuNDeWKHj/JC9KVuUNBHQiM6imY1e52OE6osmQNVsJRf4RmDxODckKm
uAAivGV/LWofIlBobhoLacIXk99C+1963+J22vArgDIn2vbiHBVHd8oebdqJup8+
AXrmnTft9X8W1cdhL8STtQjZ5jtk9x8S/tbrElX3hfUy/F1fQDLd2H7l+HrdKwIJ
EWGotWSB28jWhvnDxMIHs47m5dL37qbwg1JBXdx61KUv+iP4hrfdyxnmkTLcEZ3x
1qi4tRZ+tXBwd7mhtMPiC/spQrZ688Fmb4eVSYtjSpPummPESROkA+MyEzOrjnld
l5g0MqXJY+lMc0WE6L7yv9/LbWVLhqjJTESMAiQW3hgQf6Bd1jfAM2hF+EAz8gMa
HLgZah5zvkxaDOYmvqxQrEbBjI6XS5YCbOYHQYdUmLMAqfJs1tIN5iCinLmgEHDG
9ulCDFQZB1DEfxB6QmajGpkK4u+iT9Czc8/Yzf6hV4pgdPbUdnv08f3PPtoitfy9
sY6IT8QOZXP4fHSvTPP68lTbv1n3NKWhZgUMUtSQ2FNxvPMKGCm8781ero4cc25I
hOQ35NAgvAxRKwVVB7rblmyB+vMHTLmmn3DWVQDKmsNZgUZEbSwvtNx/POiDURU4
+GPPVHUEL8Gmd0/3bRrlcIPOvTjJlzSEU0w0vLp8EAhms3229hUWSE6JSgG2lgBw
/4gqfWLelztI+74NEL7KTtIlQzhH+GBgGNWqZue0M/7xiCZw2i94sVocXuevuDLR
u+FCjCzPMMiMAylArZLve3UxFwUb9c3JV0gAlbA/h8Sm7bx0QcNFxOuQOPoCFPK0
LjGcIocroO2UepHENEYEVyP0ZphtAGtIRtuiYAvtfvLnPBDDALVmCK97dSyKC4UT
+QxuH9T3Hro3jq/4t/xwxWH0fWF/quPz+XILDsA1/244BYVnE6DPBUUUQuruWdv8
cRMI02gs1Ckn3TMBZ1+OJuRTPtgOf2Q/zdswh9Q5gKobUO/PgcEqt7ak0Sw7+CtF
hbtDAFvAPbVT/Hyefnqu+a3a9q4HToz/4cm8+vDwOfWMpL6iEIPml0MXIVQFBefX
oHbobrDNyJeNowkmm2nPS2ypGfSEJaehEPD+MBAoU8NcuDVVfIzfMWsprnoniMxE
HqrhkcSIZuIXQmWC3CBarW2QTkSSQUPG3YjBmUvrW8ZMrfZ9d9DupF9tN+Y4XhBj
rCf51gXNlnbZ7auJKsg1ZsFzuLLJkL4xjSUXizwOPSK6ySGIui/fxdUER6wn1Rk5
IHkPJB4mw6yJUMoUvaxnb9lHSv1Ki9mgHCW4sPVbDJannOOAMF7DQFi9hHlbJm5l
aVa8YHZprAXW1SzggPOcymgS4JGbcmDh+BJRhLYUqICOrzjyBvrqfEo5ykXPAanG
rUcT/DzvZGr8Ce1e+82ELF7J6vx2pFGqFLiAGykt2IDUaEBWxq4krMAyk6jBZgu5
+YFiPDPU0HAOPjQwsSteuAkwJNmbYPIKq2Y9ZCbzUdiwQXc+svkyBlp3shvN/mqm
/1tWXSKMxG0cRgjbyiJ0RHh+Zs/Kuu3oU0sDx+p6Ii297xiBj6N4fcb5rFTPwlNd
WLjI9ioRTpMeYN4qIFj3kp5VpgikXh3UZ18idtNJRG8C7+Ixmha+QCdiLQJjheCh
OYaUyupe+HC9eHQdk5bbZWScGHHBBK7AyJwNkM2oFDXK3/vOGMXR8Zn68fiDhwCM
3Snw5kdX58fODo1m6OJfENPhsw5Nl8YTKyjoRaBD5LFMFWTEgLo+37r+K/iP1nwu
7GNtDfVxitFgNVZMS+NhlAqWc/U+q22zYFRtAC/LzAfg/WvTRMXxm6hPUm1TGMok
Qf/xjTo3YkcWlKKEMCMK4wWJXDMzJ3M34dz+hpT2F9SL7QHK4Lz5qAtCbMIcpROz
ogUp404Zp61LvEXFglh/RIW8SnQq4t8xtkkVyH8msPtQhwjWrEsv/We1z2lOZOGV
lM5x3luGizd92tmH2bXHzTCxqjgXoA0lQZRLJJWZlGawlfEGmHfpAzjEr7ymH1EL
JTOOEDwnSM8grJ6z6G75xb2YDzDFuifIpDNubj/LY87Zg1UlIHl1y7RbRAeXHKaq
cwuXnTUzcJGE5wcjApxN+Hbylv1+b8w1e+JMvV+1dYHZT4xk3s0zvSI5VuLYOT0W
G24gd9rXZzJYa+j16VOzdd+b8STMH2z+C9QgHRRD5phx7z4+CRQWVvctIEZyot8m
w2qp/Y2r8Hwh4oIhAGS2Kegjv9vmuCYk8CXKmyMRWwIz65vB8bMb+ZuxS/LgrlJu
lT+qy45J3d7ckfLwMZcLx827Lp2LdG3XMvC56x+HkGA7LO9J89gmrRjSEIstr9lC
xi3w7mi/Y2MLc8qXR4O82CsWLx0WhV2J4Bq71VCQtClaDvgETIZ+XdCfnPaP9po6
QKlJjORl+8grUYx2UZ1l+pXWam9pl7HZyiL9+C/NDQ3GN98VDKjakglFtP16x9XX
ubZKBUycXuL7oBdpQEu9jR1yKag6WkX9dZ1//Y89NhFOHNndzknCclIawI3MeZcM
Bjs2dGZ4akXGIlneWYG3gQsF5KP+Mvn9Im1YPMHNR6qK6PS+kBQs01jw9JuxMB4o
lj9quvLGn3+s+Wi5Nx3sXVVMT6ep2R+LHcLbJ1ycyIuTyWMAtGQdOrjTf1tCAmf1
FDw9u4uHAhkwYaNC01paliOtY1+AYn+rZQYbaaaPA3Og4CaYsckgn5nYmE95yWgd
PURmK8JX8j66zqkE1dEqRSkqeV5J/0f795T2e8aCuTm2EbCokBLyUkuKlpzY4dYg
tSuGzgdbei1cbyw6i6Li32ZojLzRHXd1D6YM/sgjT/nwlxysDRRwqtM4oAoLJf6t
mNggc7i0BvP4nJeeHvfOUxSAN/mYbL3F0TKlNR2pPVJk07PVMYeDYnl3DNQDAakj
BsFaBldxugyQw9RDTbXYyDQF3MwH6ltQk3yTvS4fnnby5td/Q2+rREcGwg5l8xKm
hMxssc5+vOIN0GDmsCZ3ojx6wnCdMaf35j4ji4DZZ0chCBn2S+LUsqxT4ck842IM
RKYr+a7Fo1IXT/gaJ94uhFfXs0SLO75bn9/8dTx4a95fXds070pQ9VXrZ0sxm1K1
Qr34+pepsCosEIqzSzyoscKoYa0ni1PFUI0/wVFI4wvPgOY5XEgzPzGTnG7kpJ/8
qKLvfb5LIVN6PEyhSAKyHF2zufgCJautxBp8W5UTVpu/fdexPBjRfu7VKzSgi925
JgxG8P9ZzHPVTv4IzWEAd8FDS1nWr8LCrFa2pBKd07Q0iLd5mTTV/I+9S7th5Fzi
CnyCa8l1yXqWe6KtWiUNL7Mx3RitOU4I1Ll7pS50IUYs8Zzw9fhiwTqnYmEIvu3+
pJ/Vc6iTgomrCcv2DZnzWObHKSUI3zzLLIBltj5x31PYDGWs9CD/W1nbU9TRmuN2
M5SV6twdlNbnXnMzpkQUknQifLjQySJxmScxI/4lgp340hxtC+7Pe8sZ9ndLC696
PQHJpBB/sJmhFkCy5KQSnJhbyLOBLRJXrxWQiObE+9LbUTiw4ir33oDAstbt/cMo
O2IH73KmK9OUptXEOgta1Xc/GNcVVO6PSenN3wfIiQ/4xP+52R5uZ3/cdKLI+xwg
cIJozXdJlH45PEwVnWMPeRvMRStPwD9cPgpaEFkvxOIJP7RY/FgG0NcW89xjxS+z
b2Lq9xyrE8g3PcANkPSq8CydcDi4stRMvYVSGFI7yEBP2RZ6fhEO0G7Xcc2GJ/eq
ilEENGpL+x6qwHIXi5eYCAUtpExf1dfN4qMu2bMBsHODRdhSuUp18yMBIyzU0o/a
RsRpQ4kmhNhpOVLOR1hv5iQazl+fyzIVkAtb7CPwBUNzI5IS+f3EQPn6O3/LmSm0
clWibdBjxZh+h59MZe7QiZj1vbI4ahWiFSUQwjAirAVGU39Qa1YDPpy/6/zXVqtt
tX8BMNvX55gQHXvBreSj1kMSrEkxTJZhDKrU0GrMKwvmeOUdmCiEJSRKu4V4ZOsu
xXSpWxhVg4KRR5siyMgF2ItB9vIQi/h2TwCf4Am7nWFs5L2l6LA00h+yweP0NsIR
xJ+hgOHOHmkYI8yPCJVGzzDWLJGbBoPp86dT3XzwVkNWZHauiSSCYrL0cVMlUN8A
jKI39pGq63yAKo7U4+hcMXexcveAUiLOOULGSDWIKE6tTVBb0CkYeQeatNjTQqSG
ms2mS9tXHBgWgqynihm46sJ+/xfdyE95RXjBKnyHT1/zU4SdDGHQO0mQZQgYEwLm
1SlShEkf/9rW45McT42a9BI13sRjn9llHz47S+WBpdhk9RM/P39PAcZaRe2xQWEi
DT9XaPn0JelEy9PEwot4jSAkHPkg6Hjxp3ixG/JCChLwp9CPpi5kyw7VcAuPG4iG
pboSOHLGc76vvUiTkJYR1cUHy0T6M1JatFWgs71H5Jzr4vfe1hSmszi/TGjwvJt8
mOrpwQhcnY8UpVP1udZef3qCf0tQMkhCbY5/53szPnmpszvFgzpcJM+NyAFh6BZS
Ei5RNUHfM8xqu+OAqP7z4sMkRcgq3REtPsV84b/RkQNKqDn1Rt+BOpu5VeyZinpf
lFm2clq/Jg5ykqX3fipty3FlyoiGSPmsJG8tEhPRcIa0/sdjNGE0vsQmsQqIMapy
gAQTEHVY/UFtg4/OND5LXhHGAiw5Rw0yto0RqVQUWfSDLHALwegGlqW+ssQdzFj9
MV6PuI9C1bdOBN02BUq4tCWaWkwv4c0tp/vvOg+ad2CiJzAU78kpU83dENsLCown
OZGWUjsEWx5UiKgpHd4OhKn6RjJ7BL2bZC61IOav0HaJ457hIoAW72cdyCKzHshR
994wSZqubbqIIZOQX3UKwkUfHkbRSivO4nPCnZKeJ9LBuCjGqtKUyndRadZ6o191
EDYhscO/1+76GbgmJO7Liclq4mfyEFvzTTvNfPN+01J6F9rmX5K/0xerXlXucdGQ
z1+UGbyIF15ZSJ++jZlWoM57sPou7ytv/6eUs6jxMmHEjYZ7ws5lzMlvujsI4189
sKQWqIU3LY4RylJmYfrEq4LmdmgpthZSZh+MRK4zAZxE7+vTJizFE+VWWKmcxeBM
RGMZUHw0FegBg6m4d2qu2I6XAOnRfVs+iHmia8dSoxNq6xfzQqm8K7uP87trKiA5
fuII7l8ur75v1bzNjCgJN9XDSRInufWREL8SQBxdo303P8RNKnGzucjQ9Uw5aT2v
fRgGtT2yNLeww1AP/7PH7n4WjvTg8+1LgWDUYOw6gSMhMV6YfoFHQ0K7uQ06r3jD
irNY0NvyOmCrnkew6lDlap7F+joQB1EK3wEss88SUMco+p8QtuQyjII+xOG/whuu
IVVJCqV2r+yJ1m00NvxBbDde9eAHxAag8t325WkxlHSOFfAcJVVSNAZaU9TBnvYQ
C5VEJsYJ/9x6uIpRDXzr2ftJ6BzcTI7khRtTzRfHR/bOtP911IeuXTSF8FUp7CLB
zv6faRGGY6XyNIZBO3sTtqv9Yz+r5k1nMxawDIXYEfsLHP6yDVUgdbjE+JUd7Yhe
0+3nscA6GizG2mn8+SuAFiG/31TBA0fMKT0kiv+KTOLf51CcodZGLaLBtksAg5Vn
iO4A2EHEWiOZivToCNnyyWtaTBdK/L2I1mwPTAka1h1twCYaAUKMn+xXsOC2LB7G
98lwPNcLMFZOzAMkfBV7CzgV+97NncHiTCTlpjwFcxYnKvLbFruhGKDVsZe7o4wY
g/2VL5Pls8P58tOhPvk7cvvgM6T02B7f2qH6lXigIu7z9frPk+ljIN8DpXjrnsqL
lJ+C7Fg6tA+QIa98dN1DQIwjp5cwCoEbCf71iZwD7V5HHKGYBC8yngi6hDo1TkLM
k+73D5Gcc+XwxE52fWuCrXDjkd9K9VrCMeDkmIPthI2gKm2pVI03zVgwK4BwWZ4K
oOGkf0x6U4pfq6vPYy1lVMnf0h5UUT93AuK7lU/3nOa1ZHUSitiaCvOy9rUnjnY6
AFrIjrtN0B9OHzqpFcKW3R/mwJJ+Vs87yz59ydpe4AsGJZBDOPxchtjqgy+LySXW
jPvwEcFZ7OSZbQ2zkHksI2UZwhfJHBC+hp4j2XucMeLGCxsm6GdG6ahBoHjUJup1
+AoAzgH1BZA7FFz9zuaD2Yc/GA8rIaZecrWmIaqCPgWhDYToxZK7+e4CHCs6klih
plZtoWX5pzbBD0duamd5T6F6xsPOzcMz/S8KRYcVdVKDF04jmfUUy3bUZ7Lunt8Q
Thn8iitS+8N7EeelrpwGe7kVfoGh1TvM2GX2qsgp1MRJgut6YMz1Ab+tr82dm7Qj
B/0SkNpcuBf0mLrLqVF8p502xwrgJExsr/kWCmzJJkn89sU2Jh+Ns2SYDNpzguJJ
UPjvHHLJEHjDL/dArj8lNjFp4B++8hc0m2jFmz/XdSlpV+Y6bKEcrMdi1ZB3b3oh
yOdMAjFxkv1mHUqk+E9Va5N3G5DtmzSe+sy4CS/6JNDDNQ2K2I9keOBMM237LjyU
ntLYDnPaDPnadYqpLXfxdrtgUZYx3H/pqUxujgtj9aQgWB6TrggGEBqrbwDkJAYH
uKfx6nz2hNiG1DcpTlvRRRBB5FLF2jmG9Hkrv/cAm+L2rRcs5rDfmiFupKs/QSEj
bb+guu+Um1QjDGbFg6o60CFenP+U5K4RlNrclal2qd+OwXM10hXGH81YU9FAFvZX
DlLJo24Fx9PCs2L8mFVbcTvWxZJJewlbLpTY5ycpG8ez+rf0PW0833tdvS0emnYg
3+EFiIn6guomqv8mw1ZBXH3lLAbiDpuw6SL+HwiFyOCgedwrCIUfZnUzKg7ufUA1
clv5Tx4FSCHww1sxzkw42uP3EuQBsezp+vJryXSWuMvvRFrK7nY9YksAbXmSLPiF
VtnBrJQRP2iNjAlvzOs6sb3EJxnS0R+0w/qi6/RGpJkqySJYPFc8jJ/lomvdLwH4
m4/dV1xxVlFg5EjKxGCKEbr82aRPSl2ZaVZhGhwlafM/lyrZF6aIRszjQq2aVhs5
OVY6WG7sAv5K/zMSSxLwGcyyf2W9lz+NCphFX59oKRQsrW6pGWCGf3fQIk9gHU6a
CZXmqZDqlyx4aIUiVGc1djVsdsM67xqi7pdIhyFosTJwGC6g2VkKyF7AMt8M1Kj2
FTLDKi8i7zRgAuHYnf5GAx7p2BY7o4CUq9PLCmtggLFNm5DmYmbR0bVYqfiEoAHF
4HJXyUyOdeiljea96x6tMak7OlezMv0zPi50C1BkKu7nJJIb+79wexoC8zNE1GEF
hxFULdIpLu2QrNHshl1nwbjd9pOHCX7pVkAVjh6SR8vY5oI7fRDTgU40LFDVuOPy
EuEVnqKeyZ0/ND58KlDvNhn3Ke63RebXeSDZBlbgj8ag2LDEtCjleYAT6vfTo6h5
g05d0r+c8GKkM4GGGXsHQc2yyQYVfvgQ8fr5f6tt3u554OxTCq9v2n5bDdwTD1H4
skm6slzqzWH669y9flx/NjIMzwb4uWn1BjiqqeVnheAt70nj/1OPUpW2ypFpsPX/
MzQ9Ysf+jC7p67V1ocxDO2wExHsoM6IcmGgwHWr/JoW2lh2SYsXB2nHXFqVXfiaJ
fs5dx2DhrfByvBCtcFGcoQBGOZYqMQu5FQvw3BCSwbazts2SkWnVyqzvaO+mwpix
ZqBzYwAsPQ0UBFx6qiFNTgQAPcm4DbmKKAPFhvdsBQbPQT6SCFJ+Vk2TI01FX9Mh
I2LbiuftIfSOtzlw50SZM5XzjKnC/iTTrkaP6AktsAsSnCAWoH1LQNy5clmOlba1
WCkFZsqGWXTBm+ox9EzpXhK9jc/zb0FVFovYjHPnGsOlN/QgvqhFGN67Nsu7Z0so
6CEfKdqLRkn92VX/iwvrVXkXTPCwRS+fuE49pNEY8TnwvIu3GaDuRsrV1Ps0Ku9z
7qY3ImfT9OUzJDMww8orD9uV7uqVY144kch6JC2NXzDZ72wZNO/9LwBhY6nAph1M
4jRCdQ8+t7wv37gztIxylsKNRraniRUwwax7TkAJ49rBcQlgDakWORRzocbdI19d
258gxl67OHShHX8dWogLpmz6+ahGD9p4Pu/0SHnGFCg9hpUTWCfFmlfv47pGDeSe
uhfxI+KeYGzOMjDUMuEK8pC7I9zyEreAXgTmNWdleptSOO90GEY/hGbGqL1ns0pe
idjUmuA/Paw60YWMfTsMUlyBZGLqf+sZCbstflTd9tA5yfStj/6oRCGDgS4lMcQE
oSFaa/LzJNHM83dvzZ9yYLVDpvKdKQ4rx4SJuv3gsbkTClrBgGFKJmUbdF7HfseX
ah2StDt3dwyNUjpWusJHl/E93UCoKLWNEQ75jHLQnUq0NH0u6f6rOhV34rv5WGk4
x/ojd36gKjI5ExOPTgEzGwoRMdVDFHhkw9q0V857iO5ANM1x6GLKUpl0qXMSDroZ
KOIe2b3T79/yaBmkukZKAXPAt2SnLEAT5IWKOf86vduoIW5qzicF0W2C/ratffDr
lvwKs+ihcNluv3Px3n7fY8/JW3ZRCiVZE5L9JnK9e+rvDB1XtuPM72HMxAiCx+zL
LacS93zvVcOOMLXqrx1fUzgtXCmT4TdeBv8hzVq0vwptUzkaIcMYAPYc9hlpxb8j
2mrNmPnrZlav/29owvdnkJHUkjhH4mIlnJSu63MI6UQueGJN1UhpcVlsmc9YpC3U
s8LC+6xcAYVVddkmlRmhAAQAfJc89ILQh3uTsQeloLRZQbxwtp3JorKIhyVOf+ZC
/8xiXEgBgFuUHGRRsx5qk8phkWr63drvRRUqNdV1BNdqYBZJ2JmotZqibRy8U4DV
aJGGTsHY1RYGF0znVmvT6w5WpajxttWgo0pyYClICxk6gXuqxKK0AaBR8XlZRHlR
2U3bcgpU5afxp7g28RG2/POAHf5yFxhJTZ/SxwbQ9xpgXr+mdrbAH17ToPaqGw3/
G6EfcYTrzK7vW+d46G6r22lFuClTVENRNc5nrEGHb1RUqjD57Z5YhtkoiOAKTa8d
cqgFeKZSHyaC7EtDPJV1b7upOVFwh65czGcnrm6U76ZIAwogjo0GSA9c3joTFoMO
Xc+4HcP/Fswe39WrKI056tA7r6oy0GSzUz2GYPqSsdPeCaWxpW5RJu1VOn/5Zy0Z
gz4pJXFlrpvL6VnXISXB2C+60RMU4/41oKVoovXJC+do75ik+/8wSkPR4PvZaRDQ
CcTfNv1t7j4Lz7eI09i8wY+6jl7m/i083JEbN/Mqu4k30EDTS0Lpn1me2shibjHy
D2y6XGYLWar076LRZwyFFaWmDIqwM9GQHBOmVeUQIZt9Lc5cIszuu4JNvkCW1iVB
5o8odngAdNqCg4GPw2Y/cDIg+r+EdZe/yKi9diwQaRMrORGwu1BoxTSlD7eThAnP
8odrcI5EA2Lfqpt024xw3eZfG7SLXXI94Afc91yq1QGclhsewwACVCLH92zWas9D
B8n4Gk86jBU38Gx+A9+UC+3ME8PgX7U2Drw3uHHKieV9LM+YTIkA0jwRNHLVji/E
dROTgbR2VZFhS2FXC2eWD7/Qwas4ZJPhJKT9vE1m4jLFkVxN6ZXFrB64JaZ4WMdw
xfyCglS9p4zsWeycgZOpI+T63n7MrZpOY4Bqzp+tQaPj7q5F0RYji5W9tN3ihMvq
qM3vf2AtK6pTxEZlR3kp5pI8c5fYHeWIbZFrPdAgzJ7tqxaZW1IyaIrMAIMFt6a5
ExT19TkZqJXlwWAAql3qvgC4D66YquLBKdexH9NinsiDrYLYFMGJuIY8sn6QK+xL
99YV0wj/AvPUeELVyCKENX5aDIEDsJEi398tqk7rB1A6BDUljPnVpYvtkuhm4l4E
Dzz/rfZYkJsXbg2bL4JlCyBZuKOQh6o8ChEiTsVhUOPVWP/6BfiJoKH42EQV82jv
ChBdlFEdiB25t1Ai47MTxTiJzg/fnkq3aSflQ3LRvJbaHAlpNg76VHm9cRzSzYdG
TKnP+N4a0L0PNkNokagYsAdv2Ht/DIPljRF8npMLAH0Qe//a0wEn2yEsqSSUrpl2
0qI59eFe+D/SyskdYrVo3RxuPUx6XamSI0XAsHlrRC9PLc2X3Nu/D2Gqbj37Q/Ng
CeY8OfglVlzBeetsX1veETgJZAIoTbMrzfPWkkuvjE1io+7V/Vtb04lVxprdNSqY
S3ZiyH/O1gsE/Y/wvLBwMMGgOCX+6BwmCwX7FweIUZ6p1VZD1RjOeT2uKBbSJl2z
xya4aD/nJCQzISC5Hv9awY1jaX5svkaf+GSzzlF00LC1q8Y7l2hQIEBznD4Yo/43
Fxh5s+NWgKCcvpL/zjC2vZrDKEeHfh208bG1bkgm4g+dWknHa3stgG40TpUue7dG
GyOSYc4kdAdsz6kwuJBMbUrmMGu4Xc7l9v3EVno5kMRzIFIo8gNBebtjAbffTuPg
+K/RYgl9zFpcWBn8iQeBRsgoyXIQgD9vPfSfjgF7Q+SxakEtvnBRqpuBiaNBWJ6Q
IJ/1ulHvHulPPOFHhZEjAQxPagDnw+oWn99XBZjDpj1YbEmLkxOxuXP9QarWWjxY
grfgYiNZ74xc0+MJVRiRYvvJhheeahQamR6n1BDrRVZJMLdljlZ7pNq9ae5gFp1X
czyTW4F2m7F4b4In9kcgSfv2YskHcCQOixcLQwuBSRaVYiKHhmJ/2s1AZcOZk4sM
/q4PPXmc7+gS1JCkozAwc5g5D54axw5hyyy/d/pp7hoaDfWyTUHk5/IU2Zke9msv
H+wAcdba8laFOGAVsZG4fvsbyDP48A4w1FG3FjZpr5jAM8QGzgqaahAiuCXLG/q0
91HeCvjeI6be9dRM3Nv1mbWpPvClgfVTwxrWeczZ0dAtkv3j/snC4t1l1MwbD3sg
m7h2jVWOGrjoYiSa2jA8DD5EWikVI6+hVeXHG4c4ZDIuKHkFcSB+7JJp2oPCAAXM
iVRPAv8GSI7fL9lfslPFFlLBbVDEjmT9M6ppWI/Oyv/j0zAfkdXcDCh/gE6q3VtB
5KAO7Mr6Aebb8qJLie6j93aiRhJPsoZ2dRWjhCWc3S/detzU8oexhGOwcCRTnlJ8
wOFGznv3GJ/rvXVYoUCBVWbgaCjbJuSJw6X8+Jm5ktwajsyzvJcLN+Fjm5B6Rcb4
HdeoIZzS0yLKK1XXh4kp6buUx/sQxmnujEeXf67bHyEb8cE5nl8MkVTIgSivkT5c
vQL4PMTLX6ah612kRTY9W2TXA0oQTDNw/MMTfHPclwju/XggyxTT7nZxu8AoPOFR
K8grF14PQj9iPyrTzK/b9+a+/rWU+l63hXVVXXE5jcka8A7qwSghL4al5+1Ap5aE
TT1wooDeS5Dn1HIqM5H7LFhmbopB+dDfwMphmld5RFUlCIrq4COXCIEkGTwhwS0C
IwxQ/waqvDhZSDM8JEbOtS3WCwhX5tTXXQYZQSfJIpJAbC97NPTPcyrRq7aZlwBG
n5Olz8RiGBbPxeYoBNVH5TTmyq5SS8Vpj51OHu6oJTa9xQt3WN/OBuiGrPEMdZcm
n/CfuHyxSFIZW7dL0EAgNpbQ4zAb77R8+I0HNG0ZkZ3FnFcTje9d8EDw/JpjNSPL
O6HHcIguYI+1mFnpo2MnC/hD6SYeklnY4Jx2sL3/b5K10vAMQ0u2U4icGWGkolrN
rsb77/7VDLqNbkvIVl48Xoqqr96DUetnb7XIpXghkpslmwDBpymOwJLZWEQbxy3N
Nbvn+UnUhYFWkgZ4UT367xm54JY5Cbld44WnRbVQxojXif/J57Dg3l0DUZl3lWxG
/VIit5eURIfCfgdiIwmqnTs0fsR8XnmL947lacsZPw+0LoIpaOPXMSTMeKR6+Wsu
3ewRXy8iANPb4ej95BZC7s4DM+nMkr+bMT5qPhSio3bI7kcGccp6UrHQdYtKi8K0
zobMxOxZ4LAuKjH3KE1y1ADPVoKmI+wScI0KqfGdbHmFXKNR+aa8mZ+tgsuI/THJ
44yymhQmk01AXZ4N1J+Acml+ywBqfMJ1qturdLEG08s1kqdx8hsQkxJIaN8TKRsu
ZWT3PWJRyqrRYjTRPd2YXfCg6Q4TFH0kZ2qbxUmYmy2o8sQiTKsDfvw0+beQx1Jm
USu8ZY3Uq3iB2ghY7NKYC05GLAJE8KAko/s8JmqSs7D18RNF5SdcXFjebPV/yYU/
Zl3+37K+XZhVQETzvQvkak6jz/BVrQmP43zN8VqEQMr4UGLUa2A94cLCCjiUDq+e
6WBa38tQw6deFx7UB/Ie+dqP8ERKuBL3t2dyecTzupoViOdtgflsvgJRYhx7dWx7
7spTFSltQcnEOtM21mj/bNSpp/FCxVieY0XhniFZjEp2r0AFECdGncur5JQdk6JH
9GX0i5jNjeHcTMjPrUYpWfYaTyFrmXnVo0jNEHTTeqfTxEaOJYTqJEvBlQMP0oot
cF8o+boU/6B91wNKxlLk7qiBBUb7WTds3HBfyP0Ogn5qWxPlq9/X2Ordsvcq61X0
9yqNcCdBakh4p6p+grsPNWZ7bwx6XY9tnzI7AmydZ2TOsb59wNRw3TVKxGVu1xx6
vAX8V4944rkxeqqJMK0Q3YzadYZFl6+mPOJ2s7SCB42i2KhR5RBuywh/y/SwLzq5
qgsseT/2bS54iExAO26433Xtsd9aorrXtngNomujrYLDQcbWdTJIJxYjK6VZ+0Qi
z5xJbEFwuhF1tH1QAfsEnhQX7AXzlKPaqhw5KSdAIFRKHNLV0d4gmDoVYcuqAGTn
hTbZ8mWeeYlRDDHAnLAb89XonaW6LtO6hVNkQvvb2rtTLINY8H5XsgE/chWAG2R6
zzEgho9/ihFmUuCgoCkd6MuYXNCSIu4I+FLq3KhpfQdH0mzfFCRC171xS6fZGWgB
jJ/nPM97UjQEf8e6jfD6LIy+BPma1MIVZJonWHgUsDrRXFGgu3B7IBSFbrNFAu+p
75/0BFORWO7o2h2OPgNYcHDceipJMf4t3JDQ4PtD4oTOnLvlZ06JNtuEqrBGgNVq
YbU/Tp+hhH1r0N8Gle0iP3kMJfGYMgt2wRIKehuP9vFka7QUw4zttWVpBD0YExUB
rAVVqXkyHZuLI7/JAvzYwYq3A1jBKUeuGVUb24rwQ383AgVqVZJlmYwdjTsjwc4g
vF29oJblxlbhDzVS8VFX9Kk8YYj3JhdUBbiLE29ioj03FyoIgQTNCW696TMuL2dt
FJ9otH6V3YIpmEYW/pYwcY1yH7C5dLqenP4IyOgRNfhnTfV8dtui4GzC7DzsS4Em
o3YHG3bv+7zdV7/ZKNtJp9cPKjQdJH63MDMJjzmfn54mwfcmxRs78NOuH4JPMnwS
Y09ot3G/860mpQCw/2+30p5LEv1stf3qBv0amTaMEJclUs77Q4VavpHZTwhkkfbZ
I3UeNjBriG+CVuLMLaN+Mr8146TitcaUsmE/6IpQFV4hsmZt8qMXh/snx0DQI06l
JJSnWu/2zp+neJ9nR0IPry3Mt6VFTpPVtiu8u9NWsZ7qaupYdmcK3nm0ZDY0aVYr
+NN/LUenQJhMTyWu2MJ3UZ8EKCyt3GZrkJPvOqZ+eHWe0A5j88u18XP2nAtECIbg
WDwVCIKsP4JdYSM9Mp0vMgrb58tBlfr/Dhj4CZGQkvZMmRdz0Fxo5udYziAt0WjD
Aay/3GTDkx3fIXVKSubqPyb0GXmbVS4Asi2UVgthnf6aSyFHhwgSlllBz1xxjflK
KPRnMoD2CIuuZoSSnNvgH9caPgKY6B4s/c9TcNHgN3NlbQXsS0HDAtzHt6lb/Y0Q
wtSG4NR581ijhh6Q0MUGdsFO3yS5DcM90+I3klgJ9U10HopWnirGJPaf93KMpV69
kl/ABExq+W7dgU1WZCc0N5Wg6tfGxOhDdlXm/LcRo67dWx6qa0Z47tkGRWLndIak
WZfsCeKbH5Q2cp85Y/dtw2jttMZ9THTSRoO88Zdb9toCWa4M3Bu2Li8Ma1Rd5Dfi
z94VZNXmhcLQq/o7B5EaP0wk3EsdC6pJmwI8tI16TKk1Kx7SxhnQ0Abhmbm7oxaI
roRxRXg+yNkhO+gHI8jECOUX2w1zQsC9Nt8JK1+5bYUwUnwyBi/HZdGOaS181/M1
YmiLFhidj95H92SiTFfRFbxDo4QcP19/H8rddCYr1YT5JVFE/59au2UmtN1MLtz6
FPDDj0zbRS10942ecVBlv6s0HgiaG9Twh0H5uuBOXZugh7eVWRc9M7RJEUquNECz
zV6yQFhsxJjc8LpAxDxUQ/+qxrGXK8IA9DYoD+34NZOvv8XLsBD+NTDspsqaLvlY
ccs4dtJ5Bb2mAnWHLcZ7Ns6D6ZEYB5m9zxTQZMF8kB0N6to2mWm/rsw0cmiyIzYp
18KD1dlGk6eoWO1b4GhlrZeuY/UmlB9oQUBtexqKfuZLnHBXXvOhGBJaXsovzD9e
ZYXsKT5i0zf77pkVyczKmie3i3Yf0/NtNsIVin7rfnFE8LtG4vMs1lEj4kZ4Zci5
1JL18tnsAU8/7Cmfn5M4XZ+On5cFToEwhYdRwtLeu+0XBXA/ocYwP4K3YbhRk7wT
pJ5uiQDLmj8tGp02YTWuib4GR4A1Rcr7oUOJiA7UnGPQEt6LCvEgvJt1kG49plaR
pBPMMBG7sP/zoojzDfzyGZINX4kL5kmNbmcXzOrYQNjbhBkj2ARntpHvJXuv96yD
Ae1ekQFdMlmI1PUKyGJi/tJ1GMZRZrjsOG22CyaRwTUW9SjL+P8/NiAjerYzq9Rh
0u6RCnr4kj1dKlLpys91RHnMZED3DqrYfZcYrr3oPzlZxzqGysWFxIQQfN5p4CdT
lKidSk5lNOudTxlkGrqiYs5usDKqzfgaq5c7rkXPq7CPFsImp6FpojeIGB1eVuPJ
mpnWAJfz18PQ2dEGrfLAaNbpHpuzYIb6AvapLj/5S5pyo3X22kCZEwMXQvDRQHcj
kSuY9mRsj86cCzri5ys6ijUHdP5kVVHPqKhihwxoBAhosMCYEwMWfkWR6+5AHZBI
o1ml8xuRjfDJkxiJ5DB5UJIcDrWriGUGk+tW5rcbvMovc/NGD4eekkiK/7WY8ccy
gYHkOG0uM6ywbITcxofEiq51CHyn0xu7ibVeSi9B4cQnu/+WeORG4RbeIDDSvVQa
h+BI2VFY1oOMlC6h6OHAp/VwJS2+bShJRzrzB4RBY2HfKI6j7chHFo4LyaEk1l4H
SqFwNNKdv+4debosHLnS2zbGln8cFSa3fMRX2JveDnH8B4Wi1uBxxP2+SX5bTi0R
vVW2tts/i5A2Br8cx5u5hT5i6XnOOUBO9CS1tND0HdZEL1dzoXtpkgLsItMQXwiz
XFzSaUisdINBSbowz/kPRJxSIXCvGRnhMjpg8GA9nbiCHbeq90WPb1iSIOLwllJI
M+AsESveji1AHjtj6fCOURTmtmLBl2U9atKtA+z4TB1lGYuLSOyh90r20CsQhtUD
jmhDUVHJToNjfUCxyiIOq3y4tYdm0/eXAsmPgyb7+6FWa34hY+hXOohXQvGXqnrP
ayN2/E+rGm63YN0gc6JgTArMOOKL+6PPxI52NV/77kSn46VcAujA0U9JedJ7c3SF
TRgKQARdWtfb8BUExgXIvBlLy+eOLgKiCl4MQ3FB33UnmW25ojFtKrqFI6YN5TgD
FyE/RspxZUKJtdkKxH2ii5zqM/v2k2BnIywxFJc/QTCW8ukGdqfMwcLDt0akvd+b
4qJrSYIQLHqGDKL02lJoJlRjZo5yZL49rl23HdGyQVI1CW2hxGrniHA/KwZh0kpJ
AvYf6w/WOLF3gpi8rUWViQO6LrWpVKTmNj2Sh3wJuPR4eUWwrHZBBBzfaMnVVLt+
kKSjVF83MYkB90uqqK0tkON54sj6NvpxSRX0ZNUd0Zdk7S6RXv5b2KgCpGD4Gq1F
JJourhkSTBfV1Zogkd0MND1zFgBwmEtC+8teFWcMAqydwc5MOuH7DtphR8wHaxrB
OHVOHpQlCxt+0MlhSB62uAncEgAWSKcJBwmjnBJMosln9C7QSLkJKRsM+sXFQ0AL
qNBZ4oK6QMm1mM0z8+Od7vctwAn5wGvZe4lmcowm+wZ9/Rpv4vFTd2zjrxHFfjTg
K8L7g5LH+54DTbkJt+lxuUwwTC1DkwbXx+XR10+ffv0kREo2mDtccT5alQPSgH/M
iIW5rWMJyLen8q/F99p/9xjbG6K0acGREJIP8SPWPlALdtu5WnRvYNTFnGI05rFV
QjKqP6O7KpU99bqv5RLRgh2vJZeyGiNasdrLOT8jUuOez92QFnXKDBQtOR9J1MUC
MOdiQ8cUfMgaRI9hJFopgSoSZEM6Z652UjlZk7KKMvPQy4vhrwJpDBqJwrLryZAE
y1r0R2vkY4Cly+zGTfcvJfrj8XcF6WTv/xXRirOAB+6jdY3p9IP1SjCH5wDI3B47
/5wNwqu6beasWHw7n+H75M9XvkWRkCLNuuldfG/tKkzWgUYKJDdhfsDEOOIf39yX
p98gNGZh5mBECCg+2FTKuzUl+ajRaRM/koKzbtEiVT8e6dKNFgQcHe7OyVip0nl6
4Ef1hCVzpgur9BVyi1TUbNE/4Cqfn1vD70SkWWUCX99SRKJ3Yd1ivyVTad/nlTN6
zDX7G6xJTBDEn+9QDmOZEOYevRAMDULj/2316Jdsp3TNaNk8P2nWTLqDMF4QEeyT
LidZOMa8Y1XWBNGuuwhzbVSyPr/RfozbeKGCWFgNAT2TFi0QET5CdFOhv7l7tUNq
jROTuUhHkl8NFCkcsLd7eXxDfX/w8NbGQIBohR80iWJb2PfH9bKjkoRzlPd7DXY/
dZQ4cTfPCrnlyxBrRHkGSUZagdKTNuTBHNy3wR123rOAOv0m9ZfWQWLNgpOXpXyt
JgvHGFEJliEvd6D7fn+gm4OFm9uGasTtWG2pIj22emotSoYcfg6TrfjJ+I1jjL6l
TLCIhp3y9v+ky8e30Qwy6ulAUTfls+WxZbTsv29D9q7ypwDF2lIZ55Ixm/cmQsNp
T1dtNy+ZkaZBNeuBg6l7udr8e/d0JrzuhG9WVoRZU3C4tKImVA9Py2BqbIKKP6pZ
Gb3+TQDMr0A1ZYNoH9GuDanlFOcLAheneJn8Wz2FOXZYcN1FvGuNzUK6fAaWlc9d
0hELKmGBhhaPm6Mh0OvcD2GzEQUikWicN1Zsu5xlIm65prwr7AzfE6qtPV5ln1xr
lyJgkF8vw2b5PDuvz6vkhSlriJDbrOyo2j5FKZIMM+Gn3bOylTNFo8Z2MOOJvbZn
2RBHopvtfbZJu9GhDDOOLqqQGzndAPiL0rzOve4bBsH94KN4ZJoGf99yoV2PbvmV
gh4cv105KGWYhvHyq9KfEpJZcPJfnjP6dG0DsyBDdaP7amxO9sSnqGP+9ExBVmoo
4VCjYD78+0HDcvJO7pUp+vb+qY88fATtQoRS3aGOmnpFG8dl3H90/1NoOYvpdtPL
KYURYoQZhhW8BPQp4nWpDFv0DCVEECvFaBD2o5lO/c8CbeqG1BrSPAiLtSU49ZVe
yaCQF+t5g4H3WxZ6H09K7VS7xUQxhgFNs/0AT+fY2pK4SLBcxnWUPtOhAKSziBfL
mAKPNINZUuu1x/WZt6rMJ3LZE7XojF81VUWB76H9VZ4MyGWtLq9K7VXTiEC98Xey
xFb/RRwyP2AuS4fzAtC4KXWPPs+BHny2ChNtq8Lv0xTQYVHKwHqHqwAARnl1rrzr
N8lTw5OWYAxhp4PiPAuckMzubcYNApSnUHUE6fzLNmQv4LCozAY++o5Avwn7+Jd9
MFIiZij11sRM3gIlxGc74C8+l4bGScle7/9P+iMefpHcgZQg4BGaiPNMhPz7Lf3j
2eVB5IwtQ8Ufk1kKO5weiYFYMfnq/TWHT0d8GYilAnI9bi9KQcVnJFZfk5jlZu00
/an3rjvBDRBTCgrm9S8zMkATRwoiXuxAwVKKasYN6kvwMRbUC1R5SsYBEoAqc8nc
amDMhtKLDQdb72nj/PQWYmXn+uLWbgYmfr2LIEj+MxEnaHSHVAJXdr2i/d4cLyaS
i3mYd1g9p50pjpLFrsd9J4iooK+YYUAL8lgognXB0IXwrDfRvNdVgvwD2i1kRq2y
hTNW06YNPHdnXvCgzd6q2y13Qa5qEk6AU/vwa4VYcbkTa5Ihv66zCoCNgT64PsU2
yk48PexwpImwcbu7hACC6ghbwQdLbuB4xIzn6UsuEEx8gTwgARmvvWhBOzTScedm
s+QW6ip/kyxQ3MN0+lu6WY0kRtc1Mxwia+XRrQrREq1USTigya1rDwTTTIKZMMPB
RdDBAyYVkgeSgYsWJGmarlR8UIawUYgHQbCMIeVHrtqQixsupBWTM6lp0RNtkj/Z
WhhBJjTIlzM1x4+CxOWi80RRH+qJx/wD/Vkdj/IlArqudT1V51EYmw4Ooa0IxdXA
g9LQWp5w/8zOujqy+Jzx0Q5rMY/M7op2QLSZxxlufpun+Q0xWRrQ/TRTAza938dc
baE2k/WfskbVuy46fzBrR1pR+4m8HIhLUksUD8Cu+qdZM4w+Xoh4i7rcltFOBflM
TZ9PlxhawT2AyRdIQOvmXUFUEk5axgULDcshvNDajt2/tmySm6MvUqLV9kzHWRfQ
t9JxiGY17euHw7lgAbdbQZx41F/Vaf4bBEzGzlSQ0kKY2ohXwb5tA2ZyzOlcTIZV
E4ae87BD9dDoS23hA84MJ4uXmnJ0WGPZyEt3Kds0thiylp7kV9X9gmTaO4XlhDx3
OjkFlMjr0sUZMrU1cHHKW5UR1CiYSaGwilukodQHsK7nMep7xAJ6AwDT0nhVdTcQ
uYiyN13nE6aHdTaRUkOjE/nT6YCSQ70rFLhlrySgJMsZfqFQvOYeFJSYGYpKiDW8
OLjy5D2AWc1LyhCL2g5ztLQet2hwLM7UgNrWO8YbQkSZHrC1icvbXpv5L+g6u36n
Un+SSFjtwnwNSOj9ELIX7DlhjpQQQVNRMyIkrvFtmgCKYGhaasyCSHqUm19kEq5b
L18/Hokd7z17ebaLoZkXpfgGSJumMEQioHSB+sjXQJlf/UROXxAUP41o3R/lxTWV
Sl4X9QUaJP7b4Zk0R8iBpWQu+Kvn2Y6YFLjcWyAm8Hun8W96PzxGtCnf3H+TorS5
3EYPJ+vTZWMyaImZ2BDcquzIvpVL20MmfJ+qx0aog7WWYs8dIkH4TxCGO1xCbHZX
uYiQaWpdAGfREktchTCTxjz2FQa+75aqzOLkthGGnXklkxxL7WFf9CGFui2lkram
vT2pIDi+cprH/plQVPdnyXIGTgx0n9C96J7xw/Y3lUQ+MV74yvQYgIVnNU/owAYD
3LKf+TDVA36oUwnzV5Q58bZ8f6WI5HMGnUl1dG42JBAPO4Dlkk/o918Al+DTF47m
IOuagPEkkkNWWQHCmOuO6b7FtsBgDGGrLpIJ72jauMQRYZlcH9UBjBBbVF30qbIs
h4UAeQJO1elfKr1eN+Kka5WNBukextJKjM98ZiyYzrJ2eocYJge3+tjb0O9t3Xdf
vSKFNie5891bcPDFhdzl2fowqGAnu2DLIN/sozwhLByw+LBY+s8fKheCrLzrziW4
zfJOPCAcPtsjlNx7a6g8fEMpl/s5fTv544hByIw0+w4HjgyRbs35X4BSblNwSrOY
Wah7HnP5DrlfYl8HKzGwevj0KsMxWy5xHUQw0A4q7avcyAg+sxp4m0rsFGqVxqQP
p0+qDHKvY9aqaPEfBfFb1pIm29/VsjTM0lRf9NH3K1u6VAzL6i3fWv1XOrlBTYGf
Fx+cY/VKa0T4cXc8jwC2KZqkSoOuCkNE5R2lScXHAk3QMoHAZk0670LUC2QpgzZQ
l5mEkz/qoE5ftHef29RAUvc4+GBQtAKunCL2QU1i5F2y/Myx338vhhF+qKn8M2hx
xAlwFbxkEXPi8GIopT/EQ4owAla9lspyd6QswEnDFDXvvCb1j5sJaHfrvaBsYjzF
NwXo3sfkTQiFri50XJEwk3LKHstt4uO43wNnbat6dk9bynmjboSfBvZF2/glTqw0
OH9CT5DacLgK/wgbLV2qQa94oO4nDgNrEb9dUbbkMzWJgIR/9RTmi+vJn5frw9b5
a9fPn6H3PvDUW4hky2N8d1AZ8q4Ept+F/glB4ZvHBzx8Ceg8SLnwnCBzH6cjgcNA
2aDH4koII1jxBG+EL/tlY4R2GBZ2u1mUxPNoaYjSaFJqL+vTop4lpjfahBiVrDHY
yLl7dLm6e4KSRHpVjwosPcGiuFwWNfD7e04FlsN2oFja46+BBeK4qPbq3Q1YMw5q
RqDi6CCll+0YUmRtINaCspM7ZkI8eAW4phh6LrjkrfDmZdDW1Nuik84u7n/BJchI
yCIv+f77LUD6aNekg3HCZQgPXEG312OTk1QDoNZ2vYstjzOLnN3a61OtKB9EZ5rH
pEiKQ3iLZLdbN0MSkcqDYKkEqXkUUtbN+BuD+nHZ9l8GI7LTze5ntaQg88b0GGRK
pLC0KnfTIlJb5ySgIfo7QffQcdKBewMsAG5Zmf042VuS2VotnLA/kAgFeFe4Vih/
1vPZ3dFVsPySPu/nj6ZIPwFijYMCnaF1KRcBXxm4oxRAe+E06YY7+zaRMSz7wZ9D
QqqUipb9WxJCqV5RaPPVJ4WAtz5hr49Su+VL1tXMwMsraL0eUbOovh2KxtgFhJ20
YS3PFLZpWncfuT56mxecfK610uGL8is6kYawjIyKujEbsYjX7wvTwVbqxsG6CLu9
RVO1r04N6vOYkCwiG+4FfxIAPDs3EwMWYL/j8PLn3UIXJ1Esk7MrSqSXi+FoWxB6
Wn1pxh0Uwu08dqXUUSW7rksFnVvsCEct6KH4yzM8OOwcJlipP2ydGcx+2MpAwk7q
P8/x9fBnYXpIg2pqzSxGO6JpZHG10i2Glhw4jfaWS7OQZb7xYK4wLVq/jN8mzj9v
QzeeMxRUDfUtCJpwtdZqLQyUNxHi7UM1a5nKdjBraBTo8NFSQpVbwltaEpPAKEMR
00RMnWXfpI9K4aHEFE1DjoTSbRjuss0VdFhp1B72T8j0FQuslkpOgVyzMZRmyhTh
xDl+IBY/3lW/PoMq8KLkgMxkPLW6kaYLvtU76bps82TD/xa57y2mSCDJXlO0YD8J
RYogr59arUXZVtbmSzr6+M7Lo9+X3HJlGRtQ7AZR+J26wLMr8B7JoDp1Orno1g85
F8ZO3aaITumPWKDHLIRJnoMmgR2Ie2kONATjmPDB/uvUs+3BrDK9RAA2QE27q7N9
jLMo5pCEELKiqDuZwKEGXXAimx+sIt3JjLu1jZ3GcVYQBX9VYnGbo2n7/ywShQt7
SbMy9+eU2wuuAV4tb5polOBIem4aIYtU5y2wYhCZxmulmWgqakTzy0D8l8UHFc91
r4dL2u4f4T8g/B2QlbPavA9gHyabi3myyJxK9gpV4frcZKaRq50w1G2+7PxM1Y0U
ga7UmqIboCAs6Oi4ODagFYN2SgcUKgK0Ax5vZyJisofElhaXR4NUn7wlLUnAtBGI
uHBw0AQH8sVUJ8lZlfjJzgucgAvOh8hrf/GsiZE75hg8A1vZGytBPKQ8/O7/qWo9
9KlbAd4+0rkhVuvYbd+of+kO1kdQa3Czif0TdeAClDW3Yj5qCjDQ0pvfnJQCV+qB
XM4Skkv0qnuh/I5kYE9x4SwzIdv30iTuLQF1EL5pKhHdLfFM8Zt2/oHCLhBAOM/Q
+R9L42DspaHoMMmVPzxWlGvET3LmwIlh4sA5SNtAvNPtq0M9T1TOJ04Mflcj9QhU
orLd6+l1I7kcYNlV8kPMui5Ipzw1zdGqjm1baljtEew+v94lpDJhLFJGrLtRKfPv
eaWE/isB1ly9Zr2dVcWaXbKainyrBUBiKmf/L9an3EyKP143dv8QNFX5gWk0FPF+
LYPqUf5oGDPxPOy3kuAdniadxYdu/NARjfKyZWArwVX9cnhULjJQQTAfv8s+RfGl
i3koZX1CTconAd/J7/mUuLEcGkneokGDr/UJv5HRCYxXuCV9KP5BhZyeaT8AmH9Z
nRZEoeUksE4Cr2dX1ylxOqj45iowJugjErOlChBbt2WDMAQwegH7azEcsKjCAYSd
0OVSMxq4hq4VeEbYH2b6XQtF7ZoKPdDva/AEZe+T2hOUDjBDQFuqHqprrJ8Upqcb
tn46s7Axs2zRIusILcxBIQMUVrl3Hi7o9kkrNPf80aFsoWVtYKNmH+7ei1K2ukfA
BgwLZmnIkvnONjm5hkN15oFGfuNYOY2qAFJx4kSbLZhD4wgqHco7l+9ovkFcH+el
MZPTxNj2TpibruJl8YV9qTOoLju+duhmDocQg9Xdgc1YDxqAQhTaKDatDsjyqxNG
+D8FWSTZq+Cn6C1sfp83i+xf6/GcSujs2RKzEy5y8RwW3Fdwn3+vgLETnN0bs1/R
LNIEmwKloQtfmmLiKp1XgknXEj14a3anzWNpb8QvinszCplipPt/u+K3GCuSsavl
F/+hesUWVx8VchrnxkSbRKokLpsqJqDvOkHV5see2tD7kBHVaf+egjBTCxtcS0Nv
k8MBU4/6/TOvDTVm3rkpd2RREnrzKqRP43gfk/+xxwVJB5fXZOBXIrQB/VOdI6E+
QbFzHfc0V2BrvPjNjfD6fMEclwbh1nuNDEJ2XALGNR/fvhw2HyRiTcGakKQrGyry
Q8F2ULYYYmAKhc0JiK8ZCpY3YIJmSEAE2QT18aW9Qv2rC/jv/OX+9915O58gHIF+
zv/IrXviURVpRpoKQ/x/ZoBLwtxCtM0nTpiWlo9221kpJH9zoSdgPA9ugqeMDj0W
5fdYsKBEEehPGuYR7N2HfnNRK4fBUpQPpoKR58IEVYdw5tXyPpD8Dsh88qqwfbLM
QZYPezgBPKk87FLjzwVzd42nr0f5lUe6F+PlK6AsQiQ2+ND5JtuvTrUauSDDFipA
atKk1HuqdXtRQZOpcFmvSRVe9NMzOHIVb11lVVFAe1+haZArfLqYRRkIhCLAImn0
BPyrQgc+3EQ/Jbzx/Aqre1rXw0h4WXwoOtIrqbXGoVOWcHVpebTMEwJ+Ob+gWIBT
RkGwpuW0lDPcQGS64ms+nMxh5X/V2N7zERUl/ebSicdctjI7SEddtWj2gM5cJ7X2
+6AFYUpsHlKsaavwpYyGDGP0tYLga4aLzaTiIxbcqd0CBzQhujAdwplzxt7tFqpF
as/A1XJ9NCXi826spCi62V1xObtS0Ekp352uvAnlqBxyzdt0QbkYvOVdgyrmeKGe
bDdD2qJT7OAAFCPdcUvnZm1qi0OnSnW/Qn5y7JaaXi/GzUtFyOJKsZa2NQEnB4s9
PYrpJT+m3RgQdw1Yn/pQv9O/Jl4BtNGqTsKwBjWH7mw5l0oMvE8mqKsrTyJeuZS6
LVlwZhUWJ6EFxKYtYjZ+em96eJmpgEQgtT6GdjWNdgElI4NHz5wAvuoO6naEvs4Z
QgQ/4XOPB+M07jx5TZpejrA8JRv6ogfmwHT9KDn5d4jetBDnrBkQ7Q6gSHLPRrvz
ornqhy+9xHSezIF/j2BV2DoUDpj9wwzrDbT6uxzZGSxLoXLvpNBuD/scCtMXU52R
UGQduw0BsmuWNjBlYjcWXIpsDYexFjbW6/rl4OrReNFgsyWBu+I7dc7Uj6ucjHQY
CX8CrCNFBOozuYmGm9pwDVu6tWWwaIFsHzkNHeNH07U2+s/kDh3WN6sMhLlXopuA
KRq6mlZQbCATN2fIIwkP1jmReFVihOLLt2KGVEMw0VIMRBG/IUgef6DnZTb6DiZI
+CNofpEYrFwg4KGzkm+KDJZ4QJpqZewlfhgkUtCSI6US/MRzoYKhiv73ZsOnixXW
IJa2Nig0b6rs2ak08eHpZc1AfS+mvl3y/yzSczrMvG5FpXEPSTyEJqBhvYRkkE9K
9d0JjaAtgy4KSR0vGcsWtF7zS41lvAjmIZVpUOaAhGjo9Pg29hzNsemherjj9N6s
Kyt/wux/gOE5Eq2ApTTTUKTJWCJ7U92gbKKPS1cyKA65IiOEmYbUebVvEm4tcA7i
67ti16Crh2dn5c0RZE0qOf4BPwHlvd0qFOf7gSbRNnUUccztG0cyejQUVMLlFdUK
TantGfjC/jy2+pNDyW1DSTsgMjWrFsalE8irgyQnnmwm9VB2fZlEY48H8V4VBZxz
ezpWsx4zgAAdh0xI51xbQBR/hoQyXERdERbEr76jGkZ4lesi5yL3dD8YTPc3UxQ/
vGvAK9z9Prm/nhy98Uc7IhGa0I1p1hN7bx9Is+SA7WSgs3E/jCkfBP/TmqY0ckLN
Ob4w7+ZYi/d8FjXe+uG9WAw7oDzfGcCvoPYABavoJB/e1w97yHDKYcOP0TzsC4H2
7UQRcpfyj9U740u+4sfFWZ8humjmI4GNN0E3ITstBjQORD4Bw5rUfNy1OHYAIZL+
0IqKVqYbW57IAhhUTKQ5n/RBeNujk3y2TZ4uPRfx+a0MTXKaaYWbwZK93RFOdWsS
WwHe/n/fl7ElhQqCeejKAFlY+eztM3y1FyjETCbzEJNtbpmDiHJKjoDn51vgK8s+
gd/DJj2q529SyO+tBzvTDsA0RJZ+4H8MEYxp05RVA1LVKaLHm/GP3MpxrARLROm1
Q0mV6ROKzv7JgdXz6CuF1OMDVISbBsBj9ZpXXosHEm8I9yoEZ0Jk3jkGMVVyENKQ
dLRz/0lEzd+jcRh1OtVOwUr8QUq7ftLq7p7urIUf8sR76bY+e6JdC8rJJ+37Pzzj
HAkoO6Wxcxgot7tMNRdq2eB28pkvb90UI+zCufTc7hHSdTnr+/mVnsSA1q67e0L0
wrt7Kphd/I7BU97LfN2mOfa4k5shlllj6MDrfMDc3h/cnaiIqH3souJUUPPTLCOA
MD03b5yzCidD3POoQ7iUIP7JhMzwaoZiFUO30VsFsU2rmL0YaxGitEMXMeV+vZ3M
D81s/XpmPle9h+3KvKn+HKjB2JqKFEhDnhT2GfEOcOp1hKWm5D7lF6DGZC4nIN1G
rLGgywOe+GUrjgp5XlPTQKOGYeyyteL7aEq0i6bRmfoycHH0G/IkB+FLpIbNuGup
eeH3nJoVSyOHGVfxygMTow3sGmxWZsz23+jsM3kmfmRHx4A/zYzQ39aVev6KCL51
l9P2ScLQNhuKhO86XgCv/Fd4A1UhIULYP/KRoqQ1ChTRcolr6fS9ON6Yl8LsU1Bq
NR6yh10BW9GaUeMSQ9mU2fi88MEZeOUrTO5AxsjFZ/419ipfYjoeRKFjorI/Cxw3
tMqmVvpX9UJZfKiw+4MOAVR0hdNrTutbbKvo8kn0yQVfc/Pxihtzk8hZZAxv3DVz
3rkAdwuXSR8fCNRETsmXyiTLsU+6L9HllxuGZMcGmTfo7vwdbYsBadN609eQDM8n
bK0UAzq5UQDvTQQqA8n/VQUpmYys/VS9qKgayQBL+OEBAArU64yTsFdlduzCGkHP
6uJ5tI3bp6Qm154tlGS+YFywvVU7MeSlYud8PfZToGxi88d9srBrTfpnIAzEWWbG
UeW19ODIIrS8TDJHydaRdnOcLqIsAwV8lVQCnyyAbGaNz1tQvIYdX0yhp4VzhSGJ
fuFIeWK/wlXkOcT2vTdVSrA+OuKGRV5fWrwQFk634AYo9NXUWjDPqKWlBn+kIBtU
Uw718j2FdRn1NGi0PN1BLRJ2v8xepT1wyB2aBVBCZYinhV1rxjsGAwxFvmJAmpNk
ovcibrmw2DW0nIry+09pvsv6sJNVQNnqluurttKZV8kXMr7HAZpQCuLuNAcbEiWB
TSWEN7U00/M64bWsMBIU+sA5OoK4aKKnfnApMoUlPeQ9XCdP5XpoBmxCRFM9I9kJ
gblbn36e1NwOQpTRcxlTFiKhtQWTW4AVLRblLvEMzU9hoNyOyjx4X+nkCXmH8ySV
gbRLN6K8OQBZZUozaddwuXkRnq2H14svaBKia6uy7SRCKFoh7q2/qQ92f7zLRTNY
IbQnx+uF9EiFonqGYbFEEDyPMlxNekUv1El3lTO1n99EnYr9V4/6wvrWoG6eFc4w
4lakoZOQUdd4HN+xNXCL6u6tsBwB+tzzjBCtAdElC3q9nM6dYnM+2ptjPWLy9aeU
6Vaa9+QMnNr9vmOF9Iw7vD/KaSDrKaNNzpzJm80VDvNR86BRa5Jd/k/1GcOrEu/r
YgbDdyb3URKHt/lNVzT/so8XSuUHakbjvwsgqVu8PBdkzz6/8FwlkQaJMKAA2hNW
7qi36h6aPpk6yboPreHRK0FOnsS4KkaoCwBd1eZvx6lCSPOFpLuBmJTHbECnz755
gy6XJ0t+2uRco0CdMybsG2FFh80xf52MhtRycwZtBXDgVxNjBAELZOX6fu54/a1S
dp6bcFbRQ9HY2cfd6y3gC2qRdRYfIobmSiUC9i2JcXXv1WB7x+cNnkOZmFdnkarn
4a/yJtxr9Wc9luB55R9xIZQ5AMAZ0Va0XSX+2hz1KVuBSl5SitBCV8ap1mRsecMc
jw9fr0Cqy8TK2km8Uvy/mf376RroS58T0TvnZE8U6k2/YGTfJYm0MHoR3x89WMwR
jPGoWLCc42P+ZGnUCmBP+A8Dh5U7HDCLa7kx1QxmGY7CgLw8RfYI7reN5yzW+6y3
FzoMkEUymfOI/HDWcZPkXwjX35F58q6Ix62NI6vhtXCUA1r7grO6IOJfsM6i5M2/
D7rFJEzkgwT20AtX402jBNDSHLlPyf6gFM6ljhaejWPxIMPpkhvePz3jPNPktHYI
FVteCRIaZAW9Ld7U+o81Q8bXi9wH3YAG5ZJ8yA2DSvFaM5b/q7zu0LjiwEmpwMXT
2sH+LV9mcIkhso2vYPuB5KzZ7743mQMOlGMEwg9PfiX2KJgQM/6VQQdkaLwBabg5
mbKkasZ6FoVq+J3hladqD8MTg6xXQMUqLhD70mQB8t086PmYShjLSd9X6OEClTTn
Gk71WPpmW2jnqaY6lzK5qcnY2C7Ppxt6oWM4B0EOjIi7Ft8U5aghBDhHYeALJxVA
agjc9iCGyYqDrYyBf8n0p6s3333ucz6gPH5Sll03mq4BU14c5EtJoaAm2EbeA5pw
5Q699YAgEZf0Zst8p+Nwp5hzbDhOK4Yxc2vyH/t6bnRGc9FeKIKa6S+id6konzNh
AlrPy6KpVkCj4lym9psokzkr//jiGMchgXZNATGy2ZEgKJYVDR54DGA/nw/Weov0
58pLjQnpBKoB0GqJXTBv0PuTYZGTUktUC8P4+DTfqgvk0PSP4E596DyiZxm9LRM6
zi0X+NDavobO25+GflwJwuiWffxo0DxF1bS8VA7ri26YGFcJTjBOYER1kGUC5Sop
lqGwf5upgnKklHf9fGPylG8NhsvQwZV/MO45UraMzPVtzgnXRkXTlQBn8gJzgmpm
qT2m3MO30CoIr8LEDkXfajKO7KZofeAGxFcLuUvibyR3NOYp/OkNfsBPvv0yx6Q1
FRdFVF0pRz6GZZzLJ2ooS0QMOnByCHk/y336xvcx2ayXMQYP0JgT+Wr7nCiR3l3J
JSo8tYVTsu4poIl+xJgswfZx+ipHzj3banNWocRB2Xu1A+gOVKzTIs8O6Nd65yWf
s1cztgCpYQAIevDHrfh9gxX6W5JrUfN1TEFSNVcyuTe7jYvlrzMZBfsdMVZ+5z1N
GftMrplUqKPKYI9LWTMUFMrEhx+3BoJsCC8LLPREN/EzEAJVF+mp4nmn0erbwTrK
pwpSj10ruHFMxo/CxDlMF7/bep0w5nTvMToFWsEmwLmk6Zrv7YlvaPyUQvQqEdhY
/7BAhZW5Xs6EmuJq05xrJEokw7ITWDatD4hnHgPeWmnhRgo5M4tnYDJveMormh4Q
RdGKp1wrwYNen6NCTqN5yqKF1T8YKMVNc4mcUyB3BYxMq1kgkB7rH5biBEZJfA5B
vBeuOxAcC+e5YZNr4TQoI2Ack/Rv/qmFIslUbSXho+mUXBZeux4SFYRmtKIA9u+9
51sxW/VADTFi1k87FGuaDTWWoc81+ZyoJYIBth2udlDX2ozYCQlhUq6/iRBdCEao
IjX2e2GR3YMuyho7qno0ieC+f8xCofm1YIbWFG7WR0FJhcltIZn5Chp39w8OyKx7
dioDIk3fCuFCUH7GQDxGsw54jl+QR2moAagJZltL4cWsE9c7P0/zAYlIpghnOOlq
Yyqr6wcoZ/FqDa9X4MkrMPr/CIakNq2KiBCOp4Cq2MLtFOh2MCITzJ4f+hPb69K8
DQm5l8Mi3l6HcFaDqPopUpIHmsTRsJW9rlePzBnDTbwLWGoIwTC0p/gU6kwxvo13
4eqA+9LcuzuMTe4Gip5CcEXqfPAlxNKc/z077uhbr4T3/GZ0fT3+xkWJh7Rirlpc
Hmky4mNCZok+p7GBOqeBNLZqPgNd+s8qVb9VF/KdCxCV35HJAE6dC6pfD0gpKPsp
sA+SRTQuZ28G9+g9st52yyFwXsQdwv6nIHevUOF3iCOuz/20D0bsCPOdLSjl4WbL
rHNQjGVbUW3+l7dEMx2K22uBtS1/41fZFGM25BywImXR9wuBqvaV7LhB9AyXs5vb
uQ9t3bj5wvT2DlXMVCJgIwEtNWTf2r+peQKIHOt6Xx6J86YZb4bQJ+TqgtBFfZji
pNOZaCFC0+JlyDjuF8sVKZRnLmN6ZwQ7Os2RGNqz179hj46KFHHREWMO87TC/1Z2
AGjFocwdweBXo9SnSAxY7xxcsDYYSO0Fk4zjQ9FunKEPFwtwDDvTXPuzzrvjNAFC
2D9ndSS8zudLl+py7oNLaGo2MSYX+oJkya2wp+g5sBcskOkPaKJWCl0KLmINxiv/
fhoSRzYZLvPkwdLiUSdrMIVK+WwJBc46vIiVaoyI9Qs+B7sFGw5cY4s5JvBT1y2D
PCMCns1gQyuyBxKLAiHuRBdI/Jameeyegeuxuo0KEeslwsodva9jNu0bC4DYa7/v
kHTLuyF6CrbMxiuyt4Z5+WrefLqW64Cdk14bW31yCG8rEFmkdTIki3McoE+5SLgj
HBHufFZdlvmOR4EvG4QnM/EEcqqo40nRsy8pz3w6hmpfTVpXQ7RjjMXBV27uwxiS
ylhCym2wtrXjccu81toWV5jmeJ+4WTeKWjOE2pEDoAVu0ZLvi4DMIBX1nvRhG0EF
N+djSPfPP+E7Jx8X0R69EMkOO5xHz9j5OK3UfzqUF6EvXpOqybNGOh2cXPGA57IY
QnEE3lfaV1fP8BvwOOoTbwzKTamE+QZzI4vFv7TyA1Ha5bM7iJhB836DODoa1UYQ
yB0CoUE6uyNjxrjWoxAGrNbvpnECgdhrw5KV2FFrt+lWhtx8Jmm8rL9kTw1Edste
ocu3Q70LOcz5W2WBed8pP41WzQBak2XLmGmiwATZBGe+PbTaYUDJOTmMoijM3wfw
PvkNjYlPJB2u3omIOUf3bWEOcQzde1NFYrRfI4fDvAW1CRJt6lDmzt532WVNKoGe
gIejm6SYhQ0Z0jAwD8yJygQOF6Jd+PBdFUOuVOTJr7IUwFUCV7aRK+EdY4haWEbr
n4feUBC94Dmw5T2kNcu9Wu2OcuZwbVjIk1+4junDRw/se2YsmuST3kIs2FTk5wP1
71iD+IuZvz1aYtr1ev5pD1TFqU8KWPNzcNMScu5smVJxLok8PQ0Q/oFesUGFWeEB
heBjrKmNPx5V+sPI2PPD3A6QjcvQ5SChDGpsbv7fJqW5OmfwDWrU5yr2RRkuSkfS
Y7BOiBUxibGhEdHH/ZI7a0A2emka12PNAbGrNJu+1YWNNMgCiktFgXynhBm+NkNU
fsHAugu2f8eDYI7gdbYX5qOUTkpWUdl0box5+nFPHBffQUEfTu4evYZRsSesWbJC
wXiB3PGItEnIUsXU7JAbDz74yAsfp4dJ63vQxM3RhjsyD8xX8q9CrKSuBp5xj29d
jLZmCqoE9GV1nUT4aJnDKPGmYMjcYqcUHd28L1uqUTbxV+KrznNXWhs7tN9HCvRW
OKy+kXgo0Zm3y8ls+AZAlsBC/nw4CXGXhZgbTQWUCJm/vjSezgK/8mLP0m5/daie
VZ8mqDSOwEN4Ac/43dizi7ESUBiviLftTDxP75lFez5xEl15W2ws5KOosB7k0s14
n+KZ0O/w/iwlgfEY+cq4ejcJM0w5l8ZSVvS59hyser2ZT3fzJh8PGGLIwvNg/niM
J9Cd4Am3ymecdl1Wj4WNcf0S52SVLmhZaS1RduFiis6q2pY4ZERZJw4O9ahzL7t4
5+bgZ5T1OAOqcNfUM3E/gJj4ZzB33/yttCFBsO9dZ2mt6730qpM/5WXyApfqdMr0
2FkX3yo+dAIq5EmDPRJL5egpSJpz+jg7TkZrq3GiyBtyVgWTWRoDIBRX4C3fnJaR
xbJ/nzcan1jVSC4eTF20Cxe+XQHDPBEkknDais4p2aJ0SBwthoioWWKhQX5tXzSy
wFp4gkkoDsPFJdsIcSIzmTXGt9D0Jz8o/hEvlmQOON2CUW0ov9tILztCZlh33iRw
aH/tLuX9ubMAHTIauU81h+WPFm/2rvvQ+1TRfo1yYhpbwzOd1wDIEOt2f9+HWeYG
+hoHF78RZOxDWyx3065zsQkfnrVP2v/zRWT7N+NdW/Njtit/AiMmJ7zUSjGE9r/6
AjjZ+SD5fLoBKbyhExTf3uc3s7qA/JpDEKykQET9mPaUeRMb81bPq4DhWWef5S0f
ZULdzMxeuiKCgsBVUBYLxWbeMjDy8U0aGt7IVelhA71Pp4qeonAoMO+l1Rv5KkiR
Qj24pWZ4Av/3jhwXa1sZyBqZT6231+OL5Pw1tfpa2bAXW0uJx74bZbSMv14wNoV6
neDXJv9JUKCR0ygSJecvWZcwjBEHhGs/MP+6XYWPXjQ3NHwysEt6j8RcJGmRrk0m
B0y+dT1nqT0pqp00z1nuYWuF+1HiyV29eBceOg0PsH/NGthXmE5ezvzugbhSqyCe
a3P4yUMFrT+Ei7sUZqai5tG5hg4vYe9EqRJkOQaQ/B8lFebJJXANapkSqjkcbaHv
0TLC1PlKVKp0dBzPv9RgkyG89BLv5w43BSBuhsS9v5L9THgtd/Whr9NpE+oK3nOF
qrmH+K05gpVz+mcboQyL8Lj2igV9inYYfSBH+YGvkVyRV+uzysjjgPxpbta58gv0
KkaOs1ev37EWqGeCEuwCgyQVTXsU0lUOCXQ7ouAtMaTycuDuaHxlroR330JfIrk4
GuALgaxSDnAHkvW9ZE68QAAC0ozk+Oz7jTN4O/51JF9zL4IR4Q9B/j7Szgw6CfD6
yF5dCO6SK9qMZgSixsJ8SupyhbvB8uxgscf+a3V7gGQANdBQjmBXOPt5PJfdxHOP
csKqw78MONxhpqcQTtzMnEEoh53hNKPwfq1Xx0NL9BqiIiwU9ht22xGL/AhrXaYA
pr7cGZPxGpdrHxQ8iP71OIChPrCeHFg5NYm8YGWCgzfUBaBZQmvkpV605rvaUNwP
QdttDnvhyiG4knLG6Z/qkHl9HwJX05X6X52LBpoTIuSbn7Ujgg0KUJ7kaqJsywGI
8ZFIj/21Wtw+Pf/vvCHHcmbUuAp3Uz8PDxnpRuoyG4Z5eWjkuP9jdyocgDF+PTG6
IJO+prZaDZh4bHKP7YHQXkGDgjkF8ybWeNGNwu59rq61PlhxeVJlSUDznQKdCtfz
NTD3qLHLHCE/XCBczLduCu1DIPRn68wusSNTMn/+dnpp9GjrftfqE+IHRQoxXAmA
kslaOBAy2GjOBozmzqJzuyCpXSc38ai3xBkCEnZZTqVc1WvqtYG5TRUES/fFWEeY
URN7gvI2J34CjKGsIMflzTMCz8Q1aQ4U+hF+tM1MSzlAeNFEHa+DUd5YDCKvBb+s
uNZFzwyGpAHcF3nBFpN8n60AOk0sNEtIodnuBfkZH6wehvntn/frJgmT5+z7MXct
ttjXHLD4UyBn0qEtTgnfE4nLHRICkfXDLgXnS6Zf1vZM8oZ16aThhVStEb/q5IPQ
8o5lbFL42ee86eIk5FF2vUjW2n2glb+8gY+mAOs6306emVJCY6brYGRUUmqbDd13
FktpHiSD27K0OokfTXjbSQgNUVSwstKqkViaxllMhb/KHGbGQX5/ocLv55XQcF09
xXVDnZZ0vsYt59g1CRLxbpolGtJNDUW+SE/PnMyuyZOPsCNbTDqZ93M8LcHODv2H
uYGEvCmWvnyzBD7fNv0e36uVQI0fKSVNKFUFJqQMInlEtXPTN4TIeQexY9TbFyfS
zxgg1Fwd9ICRaAFpFRDldEnQvzE8BeEWRMtJK/YLyFc+yyaZwzGwQBq/49Ed1jSC
Qz+3VUfNhKtC2mUIP+DiTjyflbbSUDqiYgzGQHYIzPAGexbEC74vp7vtLQ6Lmgn4
gyA+kABXanhT2t9nHGE6xtH1woxgcMuMDeJUF4q2x0RYNAeCbm5GhcRSeyJT3zVC
nnSGmOh7Z+c+6LJmgSYuGZpZdBkeIrtYTx7bJI160XkKhq1bzbWxbl1ta/zVQlFj
p2CWCdxJ/rt52G3ydUNdJoa0TGUnq6Xa3ODPNa/JlXMSJ8Pd7iYMsqz+JBIuKzOJ
P4F4TMRPFNwfEj/YQ2t1yz5P5jEwVgmp0qwjq9vpuXAqiLS+vyxwCcxGlGUFYaSf
qAJKVN0Q1zFPjV+6lrAAMfK3kN4mx/BhcA1+00t6bCEM20ym0dH7Xb64WxXa0qJL
Bt6w6+YHXTDzbsDjnhZOs8BtcOfYpDuHZAEuePsAwR4GtVz1gg+Fti3BSN2FjVJl
8NIrlN58gMb1q82hsVmHlSCxakMN6OaOZNfhIuE3miBbVuENQgeALUzwjsanEpMj
QsbZZLHTXglinbG89tJckUbxh/vNZkD5Lc9iAY6sOb87nzgDa2t4A0i4Kw02P0e0
VHgtMp++skrQ9aIIuWTFdl69mWpIJtqRDE+obNNLhsEnkWTzi/KB9/RLe4H/nc0C
XhpUXHaNbrgg2Z0o3UMASAA5c5198NU+9/ZgtnVgH5hzTqr4i3H2p3JxUTxrFDjR
hFdRCwqP6OIDDTGRfqIFa7nt8wvutIvck5ZzPGVC6mtm5PvH6uaFY0Yp8rnPM8U+
ThvrVvwG6htRL6NUYSrdc6OB3an0VslqQEjKbcoWW6ObJxA9IoUl0i1gKw6b6ENg
n1m4eZrtEmzNCLd8lGaoDG2q2w3plLtGHRx2NlFTNYEJPD33e+OmjVi/P0A6JF6w
Xrq9F5/XOqt1FEwRbZVLMAe+k93xZBL9RuhFr8KoIYs2rKJ/8zbq3nOWYPfBueRf
5lFM0mzzpQyb3trpEEoNADNtWt+fyapvnVwmJwb/ZT4Qwq0gyKc3jhbeb5WOaYJM
aeuLXe3lf34VrfZPGY9oJSz4j+zLKKb2U43FsH8q5UmHfOE4e4Ga8J+6K7E16iF1
ENRunTchpKZ8h2E+SleOtPldWWnp+4MSkRFXZb0lLVFdhgmBFr4UFC91SQbCndu0
3atNrKAjgeYPdxdWvyRtbVCldnBKytLf+SiJqJp9bZq81VSsKVlWYxQzDpA/g0YF
+Lu/ThIYrELKz1tIK3+11fOuxmvcVutinpgZcDony2gB8hgCdpOPVvjdsnKkU+5y
FCQaQoDUoX68qq/EHpI/sBQcqOvRrxLN9mHyrDt0MjHGs5AY1yCEWY7Ps8W74/3g
4edV/bKrFgAhTNf7yuAD1H6OyPMP9vF+CQLYD01mlcV8HWERP1hfbW9MfLwp8GQA
4tWFLZeqZJCHu0nZbrvxkteaAkItivwwYEx89ZOE4fmbBrrCdEgKM2lZ++Eoeuzs
76icBVrxpuIb4PEKOLeEQvn+h3q21TF/zU+979aGt5xaMZaWmz63BoQKRnulc+I5
PS1cOVNG/KuvF5LlNn9/t+dFQc3OL9P3bB+XYXtCm7jm/ujNIJECzinvxjh9fknY
hxdIp29ndxwwavy3bk+wBmxy7GidO1boH7moYBkZ3h9QQ9teG9EYKvTSUPvg1Mld
A98hTwhmr9Yiqj75mJ79i87tA9fsI2ot6nBMuO5CgcGlSfTEn9s75OXlFgFc2C9Z
SOVZcvW7k82TbwY7WzcTpH8/hsA6xi8SDK+Inq8vunHusPOgC5GGx49PnUlnCSol
3UczM0tL9e6VPg9obQ8UJYdhshUVq2f/R1ZZ6XAdCAzhauNEpXBav3sqa9Wbtdki
TUXinKlpISNlXkFEE0938ak+hcN0WOlB7gwfgIcZPrcr3zzl3JfacGX+RNKOysAu
eKwiNFbF/biRM+uq09HqBchXP1JAUXNDLtlBGK4FsPgOhnGIdS6cHAyzKIYD7oJL
J+3WfsCI8b3ni8i45lYllPhjCYWSrMvMd4aDEZ7p3WGV94URv6HJv6X00I022EN7
NSXiWXbv+qkuAloIyOEdj5nMa/Ggpiqpr+VHxojS/NhwhucvTr91KTIaE57xjvxq
JecazlOlCZsm5bx+rnRWqZIOp7vK5lAWnEL8VdJkTQFFCEot7gs2ESDOy7ySintJ
ryeiYQsqKYNgUAWy+OlZlC5QSRpR05fUzIIET8pkPv6oMxg6h5zOcY2crD8+784N
pA0d7v6jeZE28aulwTlr/+brxTFpNoeFzXi0PpFvPeCSnM70D5A9gXmNJFduX45Y
0l+aoT+1WS3797c/escT5yCLgdgpBmU2hu9n59WbVTBcj4RPXAgzjqj4eVqoG1gz
1ZDGHDNBXwhufgZYU0mPH4RE8apcdX1/NyGNBWFffmLag/CLsf9oUfY3qwwS1Hrn
EpkcLbZmKCM+jKP9sO4ROru0+f643T9eBMoQmMpGTkv1gUF1kXIRvotDr/d4Zddk
EzdUleP4O7ni67N17q7umPvKOg3jZ8YRlPY+7KIkhXvPL7DstrXwxsYuc/quPG4e
O+/Vz5YJcYIRgUwttGPIt4H9vhHU5dgfKZzjBR3BQnAwOK61+GeKKscJbifu1cYy
lN1racziZZgPcMKUgA1j2svg4JsHVFA7TQs6JFdS8pB5K8qasMHUAv9ALzZCMIS0
4Wt8NgnA7iRWGxQQ9ISYGdntqmecMGqac5H3iY4TqaSL6AAsIO7QlAMO+d8CZGXx
MniuztTvWsbcLH7eJtGoIaHuvD66xLcmz9wdRs/m45BS3yJjXcYzEBc6gcxKyRjv
fjB+LT1EPAbKkWArxxUaLOTrda+ZMMbaKOsrG7teIGApTc8HGRy/jVd7lA4WdcTO
rcUt8J9hRS5wA/nXUtEGMejnqkP1Gosmtz9mk8Oo6dZHEoGsQp0Y8DcKUoq9ujtQ
XklT99GgUIw3/8tcGvatWCKMBJQttZoEfozkLMAxCgDPWOL7i32Scdmzyzd6YbsP
VSct8ryeRsnsaFlprqbPcYkV5dQQLGeKLAIssi49+dKDGBdIKetW9wNPDvCGsrGy
nys+uxUz+t6yk2vsMTl/U1thXHFnvZZguqt9liMKD8RuuhguwvevsUVUKPlZOHA4
jbB27nPE18Pkqo3NdT1T5pl5SN8pgvABUFwljYV2hzKkvHhmeDCrv7A/Z6lLQjsV
cbDtlVVKLMckltFwgDJg66wCegGj4MQKqmQVqv9LD9d4jyPP0DV48lo1H3jvuuVN
SNBLmlAlMN8aL7oFu2kMZa7tr4zs70djOJEVSTukDRCVQXv6uqVZ5XyJZCnb6EeJ
LuIIjtiSL4IUUpGZZMTfnwvDajcw57byFUU+lLSKYjv4XbBJsL77TUfQP9l1zEsl
75zvscWxBiRKCw4CuF6QGiQXKNiDwzHTmbcnT3uPanFMDeY34ZFmn08YLz0c+6lh
8WBEAYOg1RPtQFcJQNXJoF/fb3lOgqksNis3B0TB2HY54AnG2Hy2rP2QckN2Lr2m
xDshpANWVV49LY7Etgowx8CRP2dlvoV9KNkQseFDR3X9ziDERC0M5+erAJbijjo9
sC+VM3Z57sCWBlurodfOg7WER6BrzVr/XRRz4jFmy/mAcqf4GGK+GxuZKuSCXfRW
bZlEDqqesJFtjTDt5bpSCuyuPh8UnfcZsjAID6QIW9P8xz5526zvjs2JtN9Q3j7K
6EYx4lpVZMWhCY2y8tFX6b70dZwNAqe6RsE8mHooESBY7qNmHsYZgpmmvTZlKjq5
GVjE9y7xaXLU0wEr4m8b5Zrj635dDZ/yHJzf+BAfRuvej6lU9vcXpO4j/UlWeyPN
8DxhnCFbf8buzUCBhmJyX8fABBqRWGr/NZf+2iwyspbe3Z2fdnrrcXwVqYIQvBmb
oMhoSY7+w7BP7vvTMerItWhLZU3pBCwAuVWRJ4nfVHLSFGoyssx1u13abQXz0x1k
kSTKeMVkvJxw7HgopQQdyVg/ZrnipVBSxcQEDAOZiRzHHFtPZDTn/n2gjducLhTF
W/VkbWt/dmjV7LyGSenTJAR5Pl2+TPtQpItC3ZVAseorzLbI+46RyF9tabi24xYs
55pWiiTU/q2nl37FgMPiRSHYOou2c/0cS4Iv5sbiza9ctEoqnPJKNADqQQm3yY+D
dX14JaLc9Iu3mZYw0ho7/+aVuvpkDiJYPqmf5aGs7brotPRsDxLVpD7raECP6fHm
6Fw2vFY609E0YUQW1N/7nmAf1AuMT/0MljxEjFx3O3rPnSJVm09zTOgZqUecmRrZ
GFFZKYgTWvO78hXKaZ7xUkcs4QVwUfR6w/4qi7TJr/3EZiqi2v6cNMQQtsLaDh3s
nShrApe8VTBTRswbGOlVP+9RHI1fkWmNJnZr0Ct7/t3GhTwRE3wHfQ96CSU6+i1P
jI57y2Rj0E5p46A2QLqv9kYvD6L2DAcX0vQwvRRTg5Of6E5iUhIY9U05Fl1DvdpF
DjdrwY6lTSqmNX/hDLD+Hp1AP/LKeGRGElg5O0EGTdm5JTd6PeB+l2NHYh7w1GwI
+hcflxFXaFaGU5TUhVKN1ODo3qnuzrXHKXC25RdoMH+Kfa0ZhqvleT6FDceiUeB5
m67e/blgFQinVsjrrRh/v8vCndSZeoC/yNkI6g8USs6aQjimX6/ZXDUO5Lh6TbUD
6LMmEr2cMCqY8YEmjU7dfx9IcsLVbNV++zi8Tu5WhQCWF/6yhxcEFhjzUG6XeZSI
NEAUMK0BYHjP+Ju+JhDcbIJ6lMYbeuDeNB6QRfhwEwpInB16Ltt7nORvIqKMsGDx
obNnDx+FwG2VMPGUVN9/qon6VFCodxpOyV6qVqWsGkOo3uYA5C3LNDCIyohW0x/a
rTExqaN7jL4qW1XFfXRid7ZY0WG8QFGjZvJYtdvzHqPBajcPkK1U0gPCSDdIcYVO
OuwAnwPBuFoaR96zBlSk+YQCfa1J6HyakHeebFOQ04aQTWoagZ5yMJxN1qycviBz
Pyf9tFpOxt9wD0QJr6XadWcfdIwj+2VnUECBuB8qtS5kzPyb2V7oa5WWw85sNTZY
fNPKG0fMAkCF/ZSXXovrh9soem6mKgB8JrKUwS1MqSDBfk2iDVRcTklOhnSorqKB
zssPuSI9f/WscBzWIbSyECCaB0k6r2lLaXFsyE6W92wTiMhDFAvt1po5Bl5l+Fgx
5kuQjaM2AP1HgQThmgKm6/3joEm7QL2XLWUgYfN2rRXjWZ4DoQZtfqLJ7lTDRPOn
e36z1xmyHAblOEeldp9uU4ybhZbLot+xfnBRnTg35IwLkwg4ddibBm9JAxEVT+as
vFbI6eu2yNzU+lCO2cvHRZ6SJR93sia4GORp5HdhhDdhCfzASt3hOqSMa13y/R4R
zFQZJeoajNAhLtHmMk4Zsc/kqdumLoC+K3ObabJyZ20dAjw3qt44iED0TSk8Q7ow
M0WnZEt9Db0ZP2W+hi/kmMR1/jbTBJBmnfJKuNZ1W6Hy32rw1M/gnrfbJSgaLODG
/TVq32i6U2y9Du3NMeWEBcB+1h9X63O6d2Njje3gLWHJZeWcM9afvZ3dBNu3rref
nuGMVn4/PAg4fog66Lohyq0pMu0X1VJbMsGk+pFuofRlxwDzXr2kBihGCNXHBAG6
dXSnvskw8jkynlfw19vXki/iL6i38UA4de80X+Gx2ezBFxFo7r4Qru0r3AEoH9sq
QdfjEz6PkFjVdYI0B1kDzRI+/hYuiSJQOSydWNFn3i7FVpqSVunn3iiSBT74hA7n
7F9gxxCU+flacW8xk+cW5kRxIcRJjY7c4UzfZDSgNaP6NhfK2/FlK8GtHFAXriR3
iu75qgEyBVuCZEobKFA2Wl4u1ocDRGHdjBeHt0p4gaJ1H+1SG1f9nfiIz4OJUgpC
Fbeh4j4gq3DrCSME8OjHZhZZziQ5oWDCrdwMyYFtRDXZErJ06I/T9WQUvpP0HQNT
0OiGRN7F9yxWLdcJjZrrXEvnpl4N0vZOo1oox2e0S4GtnSW1agBJbi2SaMhun9D/
v5RkH9rsQfZ1bgv3oiY40+YE02v4G+Aq4gpB+90XlgP6DsNEIg6rbrZbWrTQPzCh
2LDpvj7w/gBeCqQbZO5BnnE2rdaNK1BKISsrA4sNTbbIhMCoOPWIetd8VeDOaBsP
kN/w4yb1BwzSUkpypMsXKQ5vRYQU5byav5ZVFt4zGLqmikeUlIf6xFqdO2jhKKtl
XD7BSNY03U+eKpbQdIoqnOaCjXDCoN1jnr2hdOuXKIT3JZfJd74pMqHvGlcDBj7q
tXYDcBd6LjSY6sSCOnBbpZckQM2hC9lDJWre152Y3wDuGbILZ7rVAfB370uXvlNg
+nkxylL0D39gdXRtGIMdU/O8KtahyskzmC2qngSzv/GDw5mySVv/PXmBUnkk+dDV
HTCf0LpQTyrBBXUwUrtQYLKSiIJbdwQQd1OWQU1Ui8gjWl8tjts7cTaC6aDyedfz
vhHsdayIwcDYhlRDLU9l5D9EzSsDxaiwvaf6EXCarBMAzJ67tmN5bbvNtgPZVUTi
0wRdDrKJTcJd9bAO+9j8HJRD9NSi5fJBN29kzHUcafzzgukJOq462mkrHatD2eh1
41Dq5gtIbrSSRjOWMHJSjcfIFW4pXMeibfvyQj3h/xqK64VRSIb4M9MXcaHozsP1
T4EgEg7UmUc5mgLobpeOY8peIhnEmjkPkMvWX83h9le/pDighlLz4T4w+MoFHt9U
85GWGpMBJFeET7lIIDmKjo+v9YBSwsBatCul2gj2qOiTUeyx5bJx+X4DZzvol1lg
F77O6IRBqU+BKq6TNDyvuGx4lrmz1QC/iP72ZHyohq5sia4Iw2e6LHCf8WDlP/Om
SwYyrbGtj3zVIAN2oWfc9WSXoSumGJH58VMA8lY6AU+cvy1Mxoa6IQStT0cFsSUy
ublEoKnwXGudluDD5vm+7eMeX9NwhA/vk0HQinehe3ci0oEBknAnBAUtZitC7S+5
GSsX9dZQVwYM1E3wWPt/XaKcltSrDdwNQ4CnPoVy2CJjnhCpYAniGehoa+QHelNa
mRFNcJTuj1yhUNG9AifbyWpNj7+wWw9L5J6kTdYHOutTVpl2LX0itUTeMFofgSXj
tXIsLigz0on/oSl5l61f98nB1/zHi+RvYigU8/oW6pfPSPW+iISTNAJ3OD2y9FlZ
2qwp1cbSH2Rab7AnWQwlq9kD7NTJDZVDb8FyfD0rQxBXbOqvdWWWqiSMYMTfpaOw
goMMUB56p0qTJqh/v2LKPauovmIDM0pURecMuEdzAFYthL3DzIBP5oYQ8PvtlrFc
o/FOutnKjhgKwP7GsSraRiXO5wxnrmLABmSifmKc8/FdlGx41RnOtBW8bGf9vmJw
9x2a9bQLK10L8X6lA+3w3OpKnBIApYJYJxPJTaRiiX1HlM7ReK05jk5Npt04LQJW
PCMhv9h4yR3kdM3nN9TglQE2oSeWhFDrdktQ7e95RdWy6GUkCLrmj1hhH2kEANW8
OysW9+GecuDktA/rCkpNvMuJH+rq7jISUfXCZAlwUtMcCgI0K9KzAukjULyo0Tdq
e8TsjuV8MjgMqw61Rrft0kb8mRurXQ0Y9krEgTft07WqHuU98QdyoN3acmP0kZBs
T2QtA4Hw+r4KGTC5M2T7GvRXWuCyr5TbG25zGb/TyHiyktqXHmSKV1PqLmzDLDUJ
s0DYHvjN6OXLDDQ/2TyjLyXfWBxqH1X4jbw9Ys8DsO5Ya0+UFU8FpX9Qm7Vwex8Q
M+kvv878j2A421GCl+Pvsz8jH0jJkVM2Y6tQUN8FAIg9O5JoRgtdCymyJ/gY5Q8v
yZiIAoSLRla8+486SgXhTu8X1AY9tq97NcjHeZ0lmi4RqkXIYkrhj9QkIQoMk/gs
CQbexWlmm9xVzHVFwYkZyiuMI2K+L3nVIXaY/FKZDzGVy92kJCV9ouzdSVo2UhdD
uHKJAifU23lhzqM2EIFiM4Kvf+EREEBRkRpdERZ7vBIlWK5ZByoT6gPyzUnyQ0zF
LqaLk0h5jU7lI3ns7EicRwl3cRYZJoecSt7jQRK0OIbBVqQoXldDm5vbEKOiooYi
cieFbGyqUnxBgZ2z6XRsGGAI1dwmNZmI7squX2+wr4c6DvodU/dyklxWTUqA9/5e
/hiyiuq29uIr67H+Ra2sPr35xsDHn9qlpyxyspnBgZxuT4T7EL7iWdo4npc/BOwW
o1FNr3erYsvqpHFcTtj3Y3jyV4cCp56rZuVKsgR+ZUrKpe9SB/leOxZwX4QiDdAD
EG/up2ss7P4g+qRDDm811agZ5mpxAQghYPwQYvuwFFuzq3byUVSIDKd18E0LmdWV
X7j3UmVKajA4cnQl6m6OfcTaFwoBxnmOG0GoURW2aTQuwK4cTJ2mWbceFSRSiTnn
tLs8VbRUdsz6sItcs7INEM/eaIGh3YDdZsxOVP/nZ4iC42JNfOQAmGTccYWhifY+
/nXY7Jf5KdDsR7eE36N+Up7+DOMZuWtJr5ChOZ4JxBwN7BP4y+k7hAnNYU88fEhJ
cwMVMXWTaaoeJNElIAX8ILNrjBS+PkdvTrLaQsYspO/pVMC+0zNjbeeSLp42KKD2
T9fGu6G0PKUXMsF9XfEeiS13Fyiah2QjySxHEszhkJIOHCFiRgRJMkmGio2jrB1g
EKGF4dx0Zyw3WO7Efrnqq0n3IYUzaYELkWbw+RYimgY9d5lYA3oYtxOpqrC2fZz1
S0qkMRphY+2sJQgMDGy3jhRlvXafgaIgX6aXUpYNnDWa9CxzzAbej6vxk6P0ZG5D
ppB7aR+5ef/NpOeQ/jgMJ4BsIADEfwM63Uu2mil0Cd2mBg6hJnVUw1US9NJvJS/G
gtJaAAHEpU+Ge2C5Oq6kOmfjuW3a6h7gW2USn/XfykT4JqXe5Khz9WPtPcclZzpN
Qp8tq+yD2YjDuNP0rXo/gr3UB5/9O2A0I15C4zAuAuDLeWCrVkTsQQNzatWd9kpu
vAQveK0+BDHc+zbUl3zWsq7Aq/y27tWhVcRNebRlP4I07+DXTt9TuEm+5kk1m+iv
4yeRILC21Ohrert4Z1gBfsFk5FxoayrFtcxpkl5MpDa7mJQBoaZ+faTnhxfJ/5UK
YlNExrmeXKiyHWoSVnNhZsFGGTSzvvGF/qm+kJkMCz6KRZdvu7tJCujzzCXQoD/V
jRyy+deg4r3LCOuegiTv6/C56/p5zeFgvc+9F8tX4yAJoINgJQhN9pBZLGgCbhOG
kTXUim8wjNMrft5R9ExloIzR1bg/+pI7ODeP/BU1k+scc1PAwwGsvAkltp8SQbEq
E5Gfz8Jdp770f7iTgJsUZMhLlnBApS+79Zdgh+mHlAHlfNmhiXZLTeSZszqMmUay
wUORyc1hKHawyIwXxJtvSNkGqp3Zsr9St0waHtiFKlo3SiYOE4TGRb/OlC4mbLfU
3sU0pTohp7hANbisEzqbo+oj1eUI3T+uTn9h/9cZgnMD0QSKo6QaahV9CXkjc2Lm
+IaP+0zkcoCVSVTvJBX6LobclluCdLCyjDcJQjPEe2GD6U/omAh4BV119U/6wGFf
5PCjloeFKYsqp52DjJpdZEiEOnQ8n6VMAVsX1JNMnRfPzm4Yh5jh2LtJorM3UV15
S+gb5Njq7UosYX9/agsvITwUB3UynU5YPwLgn3tWpF2+hv2HiyNJi8LOjLxyv3a+
B+0Je5MgzGtCQJx487bUjtAimuhxHBXj3eKoP8tW749Mtdfl3ERcqMWnHR5udu42
+L4bhZSl6TUeibzUPUF6NrYT9vzJnTXmg9CicwQDvX9GnzaknjmxNHo8pPR7/Ach
CO7yR5YFrkmqmr9Kr63D+ZH04r51NMT53QfiQAlhxS6FQXFkhl9garNoCvgR+Dbx
WpHKvp/UbBEUcaN6Gh5MRyrBeg4Vcj+xwkQ8i7TaMyX4fefuQD2TiRozCbOkcJgu
wmLcxTs2Rss5TQI2g89RBAWWZ7SpIbrr3aR/UYCJWhviZtRuu8CZDSzyfeN69Mle
UJq+u8iacpKJHXGYMg8Oj6q+yJxhTukNEaAmfch9KJ/XGlF7e1OHnRSdczK+/FIK
ccHYgfR2GdLGXZ0Hf4zC0xh2iZugBEgL7SmhvNBfi8yJNy44thgrABeZGlBRptBV
QFaOsoguEGFmFXgMmsWHGw8D7X9rZ+MPk0Q3qUiyLU7mK4etvm6bvTUUWmJb6rAc
T2X0BESsHIFIMyy0h+PjSTQpDtW5EYGKxbYWnfTScWbwHvMXRTxHyCH4Ff6yNP5p
o+WLx7XgUu42cquznGN2rAc6g+EnraDSEUPwxa3jrTc+TkR71sJoQxwHvBDjKntc
eTQPhreKN4Mulzq7eKJsmuKv1of2VRrkXxsINJia4jpVDv1QYtPykB6fIovwCytS
3sE2/WwNZY5Ah/LnKe9EGOKHS0FuPYgDWejH0UR3C/vvPnr2w6gwGN4t1659D3Xw
8b+bBDKQ2MPt1glUcePfQFnHuL7kdlrp0U+T26kXICrgtaGmMbwPqBSX8WwX0NjR
xXrfoc1aPIZx8JKb8ZKvOc68trJDknXNjvsDpmRgOOU1Gt0B8YYHbexR15Ae8Y5s
G7mkAwipvY4qoL2vVYs+hgmbwSSHWqX6whBIwSUbCvLdXbEBn4dFfPJQ+S+YQI5I
3Ajmjxgx44QPQwFWSJ8v09db9AO03N3ChX5kIUwcO3smRVWMHjN/vvwu/8rw9xoF
wSGbrKWNAykVtZxiRL3zZFnhM511PhuTWQGpFS7SWqc9u2C9s2noukTEbRB+UN+O
2DkjyQgvrnDJwvjDjvrdpN7NZ86S0HMY66SL3T+Rv/ldh2W9PpCRcqKbMFLJedkC
hMutU1xKENYGhSy+ryTftj2onjOVz8I0NPjL+EP43+pjb9tyXog0ou15rFwOOX6Q
kUWeeaZffQSEOhB4bhNYBRbvL5YaDlw8HPBWJWi2PIy1NVPCVQ/TnomjFF1Vq0En
0fvcEKHqUd0AXUnWEtARNbjocddteABL3g3NtGsf+MvmfMjE5EJdk8668IpkqZ5g
GnhSZCJNi2lJDeyEzENcfdGz+rkP0HTyJaMvhJ4/JwWtWyFu918BV4Qexod9skbn
UHvHIL5Krlmb9SnyasGCjl6yY9VZtTSTkaB8vLYPXEL6ePzXBRXpD5S5okoysmtO
vNjJK2uYFhpETaa+ccLi99tq6PuAN2RQm1vTr1lXtK9MRkJx9KPBsk95NJVFyAfs
X5VPxIwoMIrGyF5xj1QxJkUOosQngDzXpDpCrGpV5JSUXkGCvDG7HpxZQQWq9Gci
BEC+1rDOVHdwyAl7DRzdyNVNiBnb7YVbE62LS8Di+vmlOwNogtRnc0e8huYUZQJF
nq4zn/BKQOKRxC8hpcAZH0gGdi5StfQ4LlONNXhrnxuA5yz++/ieST2S/c5rvy1c
Q0/6IeeHjObL7n5xIYe8JFpkMFqPcI2BPQ7ifKU4iC8kjU7VuzOsl6Y34oSXWV9w
MenzVzdOJJcnp47q55Egi6qxmA1V4LTMcMuctMTv/Ahiz7QcVNgMdR9pMt9SgvIQ
xSDQdFMgdguDJVVhy55Hxfdpz/tuaCM3F0Ltm+NVIHp4yo/0kyXm6sSMorW1fIOD
S87mXzsBI5sSqIUUJsdBIWRk2NLi327Uku36N3NPsx22LjxvwMGcp3Cyoxs2nH76
lTVxtn1Wfk9hiWm+peXXB24plb1Y5mUqA21rYJM8b7Cu5WLQvEPvhsO3CStqNHVi
bSLH5LCjyumcKrkfHO4yy3SrptFRs4LkWfDC09tThpwkG0I4x1jkxhjjDtiGp0Kr
cugSWcKJZuE+LBe/xm7r9sq125l1F2J9Pvjn7xX7nwBRN/rdGSAQ90mWOsAthclu
BrQaRiR9KQCqGraa1kgm2sskEmLzk52LrHsmCDkFi6UcFT1gX1F9nf3/y8NjXk4g
FRUXT5MqNo4qKaRmZoFD0S05+IGXZdkZmexujAXeF8ZweKKk9hhdc1cqQ6Dx2QHJ
HCBTjMyceAQqYFn0gTqxdBRytiNXGOligYBm1pPUQtRKJTRIwNFU+i+88DX9XqAP
h4b/flIHQu5zhq0W+ayzyy+w2yCl1Hwpv1FKB2f6Zk/npeREpE1D+oHv7S5lspBV
H/AaABS8sndQkFD65E4VZjHvNeJY1KbUFgP91IW8A5NmpduIbRCrIWo9yEr3Mwfg
bbZa0/7Gv0uEb3CkiYp2iZDYQKZmhXcTdgT8Sw/SanhqgSa7S+l5HhoLNixcfgdN
MrO8kdNuRximIF04fV+h58bX6v6tSv6vHhsS0cp6tbaVODtKv7gXWRV/NxmQPsqt
exFbfU5WBmpno+ivHwGX+bgqpDxXh0ZEdPQb+CRBhCTUC5ateq2TtGDnUTBZ8g7l
QmiBPW3nB89j1Ka9XeGnXEK3GUpSu3UJNcIWr05lwYZKzUeCE4EHULf1EVOpCTeJ
58QEg9XJFraV40IoilvH1xLXpRrJCy/D8bLvAymjCkLk4T12rEGHN2LlSPiMUfgZ
nYNt64UHvFI1cBYSrFxxGXmF60nLUeDlPGRokyeuPbJkRdm7LB/LTdgd58llnHVq
ze3RDaXSvZLjbC0cGkJTkb8Jr0X5C4Zmsah7g/ErIwQ2rQEx/WJXlRDjMGfs6PtV
HhRRn8Sq/9OTYWTrZrSI1N6NKCpjtndUEVMIf8M/EQtZ0eeSWh67GCkkEvXhEagM
bkas0vNM9SV71lt5Iu35sN5kChnNd8FN3ts1hQG+8EaUbR/42Pji3XMSykdqE7fU
oD4PJcRwsRVE4EaEb0oSgzCRfVrcFrP6hfeW2OMrEEvpvCDpTINl0ry5KqVgeTCN
wsXfVnmFmTc4RNW+/+qAUV9+5rUkuAgJnSTWrmEUjAvoZvoJ5SHJuiYTtJDF36o2
5DIHvAMjRjKg1fbnlIVod03aSK5ZpvD7+L12dT1kROEfENtHXF6kMAc8VnDL5r3v
j1id5/X3qIG8iJb9oBNLJcgRdlJluGNv3eRlh5x+FIkSehJoC+h3CNuwy4BCSJ3O
MUcSoaztrdDRcib9N0quXEgtHmosxwOLk6qXMHeDLf2rlNdpWA2yplZWp8frBCpe
pOQpOLiKkyotpfSTUK7ilJIM4+TuPMpFKUb4Q13APh308ARhAEZrtcU4vc3yVW7Y
HfEJjmQNY/w3nJqnce8w3BC80WAmN8xx52VwRyXCtXh+pIUtsqKR87I09L9uxgZl
JhevZYYyhlyxmwgJQ/oqpcCC2Frox8q3EoLJo4OW9EGjS2DadNSlUfzH2TrOIdCM
sJ+E+UNWaeZ11WbFi1Z6kxXUPdmDhCIG2R2mUqOZRJwrqCc2eHixoclpTolIE64Y
XOb7/UKw/HV1S7OCpdzMpwFlkntd/1I7MImhpSNgAa4PpU8YdhW5Mrq/Jhrx6zPn
tFd1UhoVrNrt2ZB/FEXvsrQXyC9wJTA9UixdkapCbNenY6hhUY1YP9034kIoeAfO
boPAxrec0dVHpP3258ZL7FLr3o3Ly2R9dwXx+gm5ZmX/CGpvBpPqa9cIuC1NjQs+
sRLZNJH5ZbDn4XLcahFs3JZ/4EmgRnUdbLvHSw1fcQMholVHRYr1sWVf9QyqRyEE
opgYFrvbgsyMe5j+iNHOYucxJgHpLOGxd1acUrPwPcKe8L5/rXt7dLhOdjo9eND6
1ZwAWnHgl8CsdzPrKmZfIuMg/hL+1qE7hipSwE7YfQjfpzj2X3bstjc/5HtoI6br
62IcNCO8WMCUlbdjMjAUo93/lGCIebRkFxO+ZvGMmEb8yM0/ddzASl/qsSWmPZeW
PMi6IbetCJXSWJBCfABc6NIEcmZ5doZ3IL6n06NrudRh6g485k+BlpVbsMPkS5qM
dJEHeppc23WzV0SrwbiUYOEJcYKZKJ6gn1Hhmyk986xgguFN0sLKdstEPmn1n5dA
/Qdd0uN+z9Emf9tvfXRY5yvqZPeZfuxvDIQezjOAf6pEB9nbdMNHRMEPtbjLKlTi
15BDCU4FWocnZRPnvyg+og82aLJ+g+n05ioXscf66BZCf7tVBv2Dg7LK9wrzuLki
RvinbYRT+C2uehWx45MMllpZuhCClolH8FjXnU5gP9n+O6BLMj9GwmvlJmcP9bqv
dHlnJH1Liym/X7C/kQEcZLfnOMaAfZ3bUNSj3jaV3OnqRbMtRjlR5+kwXd+FOFJB
PqsDPuwjdK4DF8WfiqJKjFSL/uLa9tdNrLVGdBwj8TfrA91GzMzIa0wWFR+1OpgL
ZQxvW7g2l2NvsCM/lEalOHFxywVVqadZh4scYW1Z42YmFJaWBnWqGSd7zySAkYr0
wSZ8Cuev6qSUTc8Ua0adSJ+4WMlR8WlbJEKjshaj0NTu1TEDYSFuVpryIxG/fyya
aRXt7aYlLjTdSkUsM8bWcPGtM65c4MhyJPihTHuRJVbOPA/ZXA8pDJuvH70cS6td
WP6nWJR0QX7eUJp7wohwQWtKII6isfcis5KVnHxWMOFYZ3BEUabtx5P6UcXh7KRL
8HIJX28f7QsZp7BXw7q1G+aQKVk2r6/BpL1sBYKTgohN8PwfDtka2UP0o/wof/kc
RUuma9MZ+3mA6Ue6TNzPGWVtXItEP+CwdR5reLMKDycnY6oJBcRkuk5KvQoAa/g6
IE33AjT1J4oAQodLeP+hb80oWSiK/vC3klqm1YGaFuo3D4eBlcxCnM8EC7pEQM7A
0NXfudilW0rRfa1w6jfOc8N0i8XUZO+BmutT41Mq59AVG0e8NbzX6+dyNJvZ8s0O
XMU8XpxaEkNRjC2K15x1FCtBBXy5c8sc3VzvhTbewLV/n34nafcaHknY0cWSiFub
6UNoNwoN9CmB2900NA9Sl4p83fTcX0BwhDqPBxBuJNlUOnDmkjcxYzfXVF33VVNh
7PG89BXeKu5iNZGG2beaCj2sgtCSk1TBQJ7DrtKL5nY3gOCH4QebSm0K8sb9Ik39
jo1BedGC+F1i3niw/PYswFNPYVEWd2qza6rfC67DbJ43/ag7J0is7P1MUIyEYtq7
jiYLOx+FA5FYqpRJIel8OmkJYONw6s1EnbO0HWqRvU2en5/tfM/wUQLteoL9Wrmn
WdHmWR9ets38pERCJRMhlW5rV7Jk+QVQxXuFFWFhYS3u5ui1QDJxL1v2Gr0JHKkx
gKA3l35kTmAOyWOkNtd1XLVngiu7mQp3ceLhNidZ3LMFK5/iwXB3azCAPmNRGlG0
/t5nVJwktktV5lKkkdcPwEIeDlqCoVG45nSoVqdk95kzVYs1tWeFcgUzRdrUGK/7
DjYPRqma5MnPo1eAFb6iCTaQXbQVQQCarD/9vhnTrP7A4E0gRgbNm3NM8F78IZWP
MrRbxWP0jFqfVTpzogSDBXUg6PFvo1pc8PwZA2VYSFXDLDHJiRpAUaxtvjWc//yH
ZujNZiYbx3TCndC+Nk693wpZ8+vAUJNCCp8yieWQUyCreGSpW5W24KUFcMlB/TnY
YLCfTBGwUmXDyazCOzAqWaAYsHy4se8abFWgbZBKK3ENM1bYc3jj8fFYPNGAU9Ll
P7WDZDRnym726/Fp/dKts4McgK2Z2sc/UlqybyDF+xlyWHTN6u9+w0krGt+9TsYE
+6hFP9mP1/UNAOPkO3Q1SqhhFBCHSNK6FoyN9AjsiLm9P+y+znAvS8cR55y8+yLK
Fyb1i1LZyc5vSTpglSF43R+mMOxNf/cxmdv5bqYVJ4CXgJ3BG8sKo92C18RFGxTk
VCnyYHNwkmuwxyArTC1/6w15XI8FslQ6mZk1/K0TORv2duRylUnoO65GXQbMFjNW
aWYVPS3P87CFCTwjGsQwVqGdzyWmTxF6bT1I//sfRzXmhwAfdiRAhgeOqRi8R2BZ
cLgkr+FWF/fPH8Gf7YMGjNFlp7fTskiI8iEgkAsFfv3KDcxbm/Ot/p8hN8/WbRKJ
lccbvOO/1/z6u2jd6hxqec9gBbOc4vkX9VBuEJHXp5E4niPZFCrnp1uPVVW8ewTO
qs75jx8lq7wGhqkQ83gDDdjSfLPQ3qtMusDT2M9ZIg5y+y7FZRylW5LcjFNwIplw
bSnvucAik6/RHBpeBTOj52hTedbszfhKLzXFQs0FQcWp1sUFw+fhSyJgGa6jghgw
0JGnrzIYGXfW2kOC+I51p3OICMRgaKl/0McuQGZZ/9XILeDYK4OGm1inaK5nKNWi
1QSkUFWa+Xk/dnptArvHQM1nPnjJg0Ye2/TcnCn6YKY6NTDPfDZM6YwLbpW1BJUm
BTDXokMZfSNudxGC1g/4LVBOjsVimBD4SwXEtd/9RaA6i+lnkN5jpnMrCjk4SzOg
WchSCh0GKl0IRdLKOcIyypDa2GqgMMK1pGgczp0jqMfJ47k21mMSV8fTdsRIyWjK
2+Xp4LmUBUd4dQRfG8wVt0Jhwf/Q7Kl/s19/UjvWq+Fw+xHXdKVyao9gBWPnq22J
WGxmyoD5DpB6MDqJo44vUMCWZRFxkgQD+4lmThruAJNN52/U56HBPedNzVuMhmUW
G61LLJhtbGJ2VYiMGUW78KaBMH961Y3DS5w7vQgxP6ojjRbndSlwijdvU4sj8PWj
GBON8/b401O0vnedc9d9he8vZNos+LtBQysf4343K9Uy2/Sw7/pre0WsgmUP4zFi
WmEAH5MSLUMv6cypsHnDgj7Kkecs0kIna1z3I5pPz3McpU4sFB1OjjEj0NATvDri
ULInbPexAEylPLGT7mDYYQQjxTWGS783rKB175ptBHW8YTUTYEv54Ye/0V5j2gjd
wfvcNuE5QktRl4ogL4Bp3edmLIwwtMkEAbn/xJe7zLsIKghfZ0XmBkJLABbc6jkQ
uoXY5JqTIZByPU9p+U3KAlTY85Y5Kqdc8pQ7YpD0XSnoHcD17qby9CFTVwngqLHr
8XLRH/lnIlN6jpK8r7ntOv0QBEWahBS+45UHr2sCR23pJKE6bILocCpiPNsz/42o
YN0+6Xcck4PjTne2nQrfqaj0vLbzLFZFt8BRJrpcjdw1dk/0zb43RcTDXaXqQSqP
4GmaaRkJ67LnOy4wRugmd1JZ9aAuPKwEQ37P4faCSSlOziFUjO5LYHc4bmm1tvdl
9M6Qr/Jv2DKQC311LvFc6W/RPB9PfU4WW9jAYJHyRSWjr0SbZQDUKGUrQvDR9oEG
XfStT0wkGpp8/V836ONsZvEov8TuLC42XN8EuEe/b7BspUAequUdDiSQtME8AIli
QObqjmGAj0ctq/prwjbXJslOoU/smlfqMJbE+N4TWi5XzdJFk947k/o7VMjm4OZ4
EpjbLvLUIXXAHDLoEfbOE2a+y2LK1dAHuC6iK2pYmMF1ZqaW5PUWcUpWpfSresuw
ekitHVQcXqjq7ZBXLoGWEjQb1px2g1VAjuNlrTucLkJESDkhMfWTYPaKBXaQx/kz
W0A1IMO2dAXHgpQsVUJRbSXw/fa8olUlad6UBBeXnO0Zc5P8sQVPNkQzo++0fe+Z
yoLyVL3S2gYKvcKwIItEUPzAfNRQ/tMmHE4iZtScUg6rcLc7q+XHHPg0dbbTMIao
jqRY8YwnFlrDtY0MNi6PTLB7Cm55Us5VNnwAegAvMTdpl0pdoWhBQWZ0Y6xOabt+
wmmaq7pzH1g7b2n8NJZ4xYz2Tnuw88D+o9hECYkrhYXqaLS9+CHCFNZtzcpBOPfJ
gqykGCz1/peqdQruNiIcLKezdaEaDNFzT8CvJSI9x0WXQ5ibLj68KLvSfE/lBnOA
CFHHrvROLA+6aNQMPw70KkGEfW8MdKED05L0vxo9pvxnPC83bIb+g4nxH4Zf+gMC
z9IWCxMzt+3TlYz49AuXXrpAOgxzZGcCV8BXEIxJrC/1WvQVUxz63TjJXun8QOxS
izQfp19cO+QiAi5NnrjQiNq6EiBhN0DZwq6F5jTbPEPYipHyC5mBr1K/oIEg6KsC
Ieg2FGsLyFm7n2dnMyN/w0xBZDAtj3ikyGCOMQCs5OYF44FLepFSJjz43+znzO9v
7iDun6i3SfeNZRMCr0B0cVFqQn3FQuZRkp3N8KMATamWhSigDPIC/XrjA5rhzd2O
yhJDml8WeFm39KpCW0waxwf/ZuDBR2ILUUeHWkYsuzTgwQrcrdpKurZ0gx1RwjeT
qCiFGu6X0lriffQ/Vc4co70TeI87HrIn3soZrV4KRzTQqTVGCDgcvL6nIY+6DprT
CRKmTSgQfKprVXTIeMgC0sprwdIQcbQFoaUlCdL3QBwBEoE14cCLYamf1JZvOSeW
U3KgKy61XORdevJr9eE5O1nSoOp+7J5l8R5PNgnk83/178mpd5kL6hD/rBfHBMOd
PE0mgr/LWxZreqX4VmDrUeHW5WbrfUiQGv8f7MqxAGOZNcmXErNc/mDjH5kMAP3z
b5gyK2KedV/6IStP1MOgGkYjgN+3duCwnc1f3KoSnMhnB0qWuTvFwAL/MiSHaMgP
jfJh2MP47dq4PooyHSDuYPcsPpvcPewbJI+tR33XXiJ6oUYMHFIBabKEmLYyJEpH
sGvRmPyFBFe/AFHUyLk86PsLHz4zszu7/KDoFMhjeD0vZcnaZzQthcO9WFnN3wII
tsqodc+vZNbSwqoMptfn2MQTHOdSLBHYBLSa5/++gtaeeb/RT+uV9O2h0+0j1Dxn
J5v4I0SmQUdaSx55XmxslD5NQKeV+QNvYhwYtbBJAmNZqutoFtMQ2bhsrBPshCwQ
wPCOkAf3cZbFH/wh7NgEyL1oF5hqt2bbW2uy8hkZzfFg+x/SC2z722ctC1evJrsF
WXTgG4C8MbViuQMFx+mvyTFptlo4ys4qaHoqYLUviG5gnkF21vKbtjZyRneH9NWE
sixXcNMOfRfMtXKS2xmBSxNZEtckutH3UBH+Miu/OtgScx1xYB5IEyquyeLc1SZg
RW04j37suoOffMEv9J7qnDs5EfMEXh3lpqh+wNmzhG53dNzYx6aMgFSFnsXiE5wa
uVJ0bZFD+JLIBNIMoc1Owxc+T86PAigz9cgKV0XX8AhzdZSHbfol5p0Tri3734G6
4dOK6L+2qbDukbg9fTPFcGL4kN7AMqf/PgMqCAo4Pu6RTc+LdSCjzc6PYo2dPvR8
r0AnMFipaxiQi0Piz93/ZEv3CqENNVTq/FjXZGKAoocJe8qhICqhFhuGjRZ7o3cB
A0J8BMh6Az19dw3t4j4Q60man6tnNEDRH3pWL5s4EsKA+QmRBeZMeIySg58REZ+p
ovpoxU4AgS95wfPsxNlns6uur4y/VXltBB9va5ZHeIpVBTH/5JorUaYoYms19FZl
P/TNK9D+5Zff1zb4k7X+yN0MfHx/Gi6T9lZKtU3HK3dd1WQKtUBe8rJCeHKkxk+V
1uBYn+3PPQbs7EjUfRYub/wpJqM3JBXbGdErfMIJfdaxKPG7nmK1kBS7kJ3HXdfy
NMmr9B1eZXPy572zEAqZTE6O+fkMH2icKX8lrEIMRX637CrXgOwFqgAosNTc9brQ
rxmRWmfXf76utPhQv8Z+XZsabA3CLsJa/BEv1zpE1gky7ZVuih9f7/N4KKsQ/EWG
hGU/YMq1KrrftMjB7Xsouom4/qa8cFvY4wvE/DyAaelRA699iRMSZfrhw9ynJpiD
COqRATYO567QX7HI4OYMAV/n9TkgCRiuBwlZOBNw5megqnv2nYCksyXYwKhZ77lr
vDEPqS6l1IVzSoE2LxPSWbAt+3qxXxzWf8UDwm36BjfEUHheMupnmlfNQ3q6pLuo
fQX9M66iKhUTEnFzvXsNU73m2+GTL07+9ZkwbM0eWawDP9W67cwSXdzykldSrZ/2
sBkP4obgSeFoVoe3jS/tqruSVM8+mOuzbYzV80jWSA9vu8IGAVLH5SnZF6zk9i5o
CyGwzhAMo/f+XkU7yEKjJSEBweqn/CB1I5OJYnmD8gVoYt+THQZFO2gj4nuNsnpX
aqeGyIyIBhLJX9wNqJXNUdFvjSg0Yv/JEC0hq1yYi3vgIpfu6cgXaEr73p6Ee2CT
6p7ea00m+JCqrXPHdhZnHC1d2MLv8FPkmYuM022XHoBat9KIWN/NtVL6xoFQXMxY
sJkTZTwUNiT2TjKcy3CqtCJL8shSsL9H2wOYcvKcVRe1jHwvIrqGGkFiKBQ/c6Wf
mZpwCUFCOzTHvAB33payYMECSxZBmD0FYjB2clfOJExAeS6u9cyhW3GgvJuXMrar
TYmRC5fiMmF0GOn4HSnsnjSGn+khZe0x1L6qAkfRXGG+EmqaKIyeF56HWDoPkfLN
v3q0R9nIq7VQCg/hqsmYCW3SS4VohvKRAy1QJXanXZPuH8vsf0dFzzqDN/ADMjTa
4oU7MELAU03wOPWCJ5Ll+mKaNx/4UwFWE9uWDo8ngsAXCwSdLjKi6aogpPlqfzoG
E3+9XSde+NEnOVHlonculrOFosyXK7RmJ8c6A8HTM3P2eRTOjKhGKPTZtSd+h0pH
488fT6Zna+U1/Z83vXyqBCE84iWMuvc83lr6/3xShDkJXUuMn60IWs0c2AcPAuWw
Zd+lB0PGXjdhm/4RF0hPOj8rtK3fr/JODUNsDdLU6UAfJll6+n/knOmUC2/XL+d1
rKdUUfCw2z14L0z2CAsA7NamvrLcJtdu9VjQ19C5L88Ge/NBouNecl851Id6vQbk
BUbq3kz4knEZ/MMpPGF00UuiaqupRrQ0v3hg0SQ7tvrao3S6HK8KvYgcaYUWaS5g
jv014xhGswv+im/FyUeLxrHfsmwpDvr0Y22TGVV/t8bsrpTmxCR5DYGvaFHiwhjr
i9W8juLY5hqewa/YQrjaP+4EN4vlDcIGGuUGiTrtJhxTv5MAX4ccR+LSNUH+SRfr
72oFRExFecZLROngys14vcTURGuQ4eQgdPP9X6SCT+diOQLVLSOj+yhUYolEBWf7
Il4P67CxA6IhwlkQH2a+t0uZE5ThEoL1NXpZu5b49TGTTr6uLImW+00Ndbw5b/z9
4Yd/qgdhPe8+HuT6WvIoXXTUoH6f0uIS+7w74jcYr9M349yfKakDQw3djN8HVWip
nJI72LOP+XOpPmH+6LfUMKSCOQ7OMf1OBgTW4ug1IabTbAdi4DIOzKpXQZv5Fkko
DaPzJBNuwgeKlJAITWmQ6XptSUAOtKGdMBcgzdIrQpbcwIIdk0x0eEs1pu88qjmZ
dGSRxmU85OipjybtYbLYxhXxl1QBmf2OWHnAOyWWJeW+L+vDE8dk7qULy7oWWP+V
i7UOvFYFJmDS87Dj/wKBZooh5GVG/vGJl11ZBcWApIyn5JYe7OTyuK6X8v2+bmcj
Nfe31dDx/lvFQhG0X2yDfsJMVaKbo2TG5OLeGRKi7NsnreVOWqf+sKw8ZSJIekER
EqL+V4jjlPwJKkyTPt+eBCqiTIYGriV0qZP0j68KB0JuRKxJ4WuuuupZ1Z2lIRsO
jGENPZMV9OevsbEnI1/TSPe1NiMPuouThS2FtlhS6/tSd92OdDEz0EPGdoJ0arhp
Q0Tmj39CieUN0sb7sN2qff2btiVw9fBbL+izhRwur19z21ZpN8vs9aUrZljnTXXB
oYYxwi92GhDxWuTYLypzVlUQBThAvXlnFrmE1wwKFtX9ZoRCkmhcquRSt5/5g8U/
sEfpuB/rEIhVmqHrdXpGaH2vElco02WqvewgrASgjn6eONiHD2mzEuKSIhFPhB1h
uvTDHLQwxnRxcK8snl12+X/2LEaBwF3oxg72DcAphNai6velMY85zBgRdLpnzLy4
CghnmXO4SdZ+28ofZ6fTKEkKfDkbbtTNHmteRGRGfynsurfETkg9VdM2ptV3FM64
LVOsggXPXP7t5V6X77vc49ZRIf6NJMWVJlVk0CXFmaeau6MbmXs8aLyL9JvvneGk
Gvol6L0D5toXjnM9YrVGM4WtJgiuGiPtfuanWGJ4Vc9it7VPcSIwvQ7o3x2Ful6S
YR1EUDX4lyoCiqF5r9fDcdGiVPz7MyTm1qcfkhAg0eroEe4HI/6VJCzSlkiXqzGe
HkDUg4Hf85TbPLEdjoy3KEe2bkD5Vv1xARmUfVwh8+8vnQi2f1EutA+zBGTaHzHz
yFdPu7GrsjCdaWyvIIKzIJswRurly9r6Q0HPyodehsusHrVA7+DpTnKVPf1A2Sjn
CQNFXEIcQYzbrtUpCFVssdpTHQyhfvVhSS8gwohPd5/cIr1MsgVtTeSQMNw2Eqzw
KONNx3vg4EZ2FG+aJhiAwnuMaVFacfSv2R1cTnpFSl/1Dda7yYD8NavwHrir3WRD
9lX8g2R3vV9E1fftTwerp9QABgh7cOhq3PXi7oRD35UvwFQbrCvB7x+jZ2rkZ8x9
caHkGtg+KJ+/kH1eZMm0+sqHDBxqZOE/71oNqHywh7lPHnq3ucLTnlJNnlGNXe2S
5EL+mDhkP7CiniuHVyvqTRHxiYMmJC/on7xQ63U/2UEvkewu1gUmS7Xj+rCDRJkO
0fsiVZiXcSBJw2V1kEZIEfJ+uVGKfGFF2c1Sb1+X1OE/UEtcGuvFojJFoU2OQi7q
C5djNj2sMjhX9NMmGPJ5/Oy4tgNzkmHEox1vI/brgcgHEZYZsGWq/8sJtnyFOKLm
7BApEstBtOHbZRnvH7TMCBU+doDRwb6X9F1+h36JED4qf0y0me35mhnB7FxCpXZP
3qbrGMo0fVnfmlyrYHjFtnvtDkWLhZA6lpsqKwiYIq+8pqfVsmojt25BkoS/Nlmt
qQlsN0MQMRHxJGXJEySk6RfM2rcvrtvoBDKzG9WHtw1NdzEVRYag0A6dMZJwZsEh
uArkgN5nsRV7VVSFaupWj3Uz/SCI8zFROH1+VbDfnwJH3spQ1RuN+hg6ke6X+u6p
6HboLk1NoJSLLPBU3L60XYg+9EtURLUN8KAyr2s/fBoXNKLWVmrlmESsWXDdk9UO
n2gXYxsYd5eD4FsJvXzmSR3Mxcw/jrWlXSZy9JxaILVt3fiMr82BEOrlyiZtf3ev
/JbeR48FQDC8ASDqaHMF8ZbUh8lUUivY/wVSHw4eRdf3Y3GbsS6BMMLvk6Qdsg5q
85KgvwHZTYZfrWCFrJLgxipIUt1jx4RT3IJfVB+Woxp3IbtSIxbhKO4SWcC/luIW
nB5niiFtAaUyEZWbMqmM4mbT0NKdz29YYJtaWN4hwlUcfEr4IcHPKeQ7txlLOjlR
pZq+AObVUdmgs9uP9y3XMFSfwqY5Io93zj7FePkOb+b7TfcVk2FV4rFVn5oJ4rCw
TtZsAggojI6I+PsfqmN86U++wT8EytpYy38wnKquC+eyN4G4YCDT+ez4r3d0CF+0
kGGm4FZaOLdcGpQNENTKHkTQRM2HTTrE9scjIlbdfyACbF9CCkYGRjYPCR5Td9hz
bGlWBdDSgB6RVlRKVGPocvwTITWFCrLTQLVq8tY+RvfRmug9W6FqoMazSk/qAPxX
PHJFI3I+FVXToXAC7tC6MYZXWNqrBwVPhAXbOYefHlDdnwAsIJcnjxeBnHuXHsZd
KX1DPzWjHFMZMYUmnsGjjmnort8mls3dzlPCl7yXxUerHwuqjsS7sGD69jXI2X+Q
GNN248SBirnf7caJ7nq1grmAu0hnwqUA3APz9Xyq/O8JdhexgwpuJLEiyvwALgRc
T/0veNkn0i3YXMBZOSzyL3NyTOfdFWM8k1zHtmw7Y1lCqO1lXY4c5PeZhF8CjYlQ
9FpTTXRpmnE30bHzAuQGetabaDUByTM4Lqmgx8E2RhbGlYxMFRG60pPSVg96qwFE
xJa9WAKoMO5fpw2zeU8567+q9JplatZxoRFoeJWSq2el0+u5eqK6VZDLC7Axi2Zs
UMNhyrtRkBsOWN5uo8H/CMcdReTNeSR740htMp2EUjkAwG1Ok1tStsjPQsNbJbPr
6WKLqeoj7BLetdhRg5CXaTXPg7KC25uthSKOUGSTeqQ79JE5/KbW+VadUm166ca8
/vA9FlgONE3TMlUaF7CgEZ7bwL2g3HduXdLo8HspzR+3UXkxkC9Cfwu5okXOAPE6
zjGmAzdJTr3kitawqFNzDjIAxFKdLovgeQS7mPA+a7Ap0JfdqDGNrcMSgEsOsqVq
58f+54I0K8CLf57onNGfC6H1dZD1OVJebe2gA5y0392z2IZ2c9rW7E/xIoaA+irp
q93LzBKbVf74SSWBv5QFK+zSmT84l1ZF8r5qQ+qTIVHRQmROr9ORwGC2rR2fnxgR
IteaJH3HY6K/iP5M21tUqu5DFIU+mECuim+I5Ky2IeO422B3M03iOA91nkv+0A1I
wLxFmK2JLBbWzrtr8GVT1KCXuj1nDp1JMOEeUTdKaxcL9XHOdfaykiozvZcdwlzh
kNnmqR8Kt6xlRPxgoEThcUs45Mau6h22mjgNPgw1KoJV2dYGs65aSxnLJjjRLhZg
LsurakHKPh9/R3n4gJ1PlERLIMYLElB0LOLofJfkFDJ3JO1vWixwQ9jNX1QghUxO
R3QNWLXfhycbtCFjQqDIEv9iX7NTdvtzW/LhDowVC8zFJsvLY+Q6krGgLxMVXBfv
taVKr1KZc8KX/Qq3gttG3pSMjpCl1v4UD4s7mKKXL6HTTy/DwW3tyQe22eEny4uR
06xUrpIxSf5Uu2H2qKzhIJ/n7WdYJSrkS1ApDMu8EXYLx96q2klCSAT0RSmP8my2
7RD7sv58iTjvbKS2uRsLJYn3UocFeC7GBiFg39BfpYg96yGa0Aoz6tSwFcCROR1x
kLVMp+ic3MMNJ2JElkm+A35cu+J5CKmRhBMIaWdgqdrMdqRljgHss3/GPuKHADm8
/S39922rDB4ELLIO3N1Ggvn8Me4nddACMh5NXYYyLOIj8L3/QM4u9QgCar1S7DEv
8QDsWyosE6EOIjOAiI/Xd5uYtddr+s4OjJjQ39Z/OQaMm1Zi7n62F42c5ObUjdXR
nPUp7kGE3uKD+hPeJ9pXYB4KaCgOvfZbgaXZw2dj/L5aMP9w5MsTx2uaexWoGiIq
a4Xtvb/34nzMqCymgc3R/okEN04p2uLqAyEM8QnN/4sGUgbUy+V27Q5CDo0m3cyA
5sxmudvOLLQvQdCXSfzxi1TFnKksN7gKNca9MbaexZm5y+NqFZVF/reWLY57Wldn
53rxX5akWokWgWRU1yj/jOJC9Y1fVXFoJiSu5rZddl3c4L0K+n/F5RFrgrcJmBCj
WRhxE78WjI/1QSnNqfVpnSspEAh0MQ6tUsxVtJkZyhp3zWi+KpvU7rKWwy07AIyN
smvst9H8af5w1dppD8EgBUZB7d+aMfpT41IeCTtVTLFJK+EiLExZSgxZtA4Sagv4
Iyk3e5TgQUGgy2etJblo5MKvFE1AQV/oMbZC1QMcFHjNi2kR2xxKD9XrG//VSjVj
tdex7rURQ2F1vASrcaVsK1kg9c1pQPmeXEan2trlnxbDut3FidK6J89c/FOXtVAJ
MvQNbcF8VRTFKRdF4hmQrIZv22l5WWdmovfh7U/V9RsCxOUpKRjRWKSM+RRn5xiM
5wGgLf4WkNXysDAftvXJBgm1Q4GJn4BgMwV1bdykKEDtNzFCK8Q/B3s5zpBvXltl
DUXVaRLMo5lRVSJf26fV4UhIFac8FAKUvGtlr0gmnms8zb1thzXIjdG4ccKgGEu6
1dU3FxebCWS+G+6us/UOAC28nySBRnEO11DjFvG4IUZkCDkC0pMjbj5kl8q3XnJY
3qBxWOt22/AJFfZ9QJb804Yn1gCXSYOyvPTIRWUVGmEYMSBDGpXL15gSXyF7uQcL
annmC0mTkbOe679ikTLBYQQ4Q5/fdiG12cmI4D0m7DmiApbfQoHM27uXnSxjXPJ0
M0pawaAhGoobEBLHoQ0S1tCxEBxk7Y6SyhidLFz9HKV6XBaZ1WjW9QLl076Ki9Hk
nd3KOFP7I5R5Z1MkHycp2plNIKLPiG3UCXhIF00ZbIyoE9HAwirAZnOAaRLchIC9
JAfxHDwrK6dherz0U0iNYs5Euu6VMNtHyp9xKYS1HaA2s6D4Ip/21gwrzyph6css
jfDbUckgJZQSsOOc8bwjr0kcddlXK7QWtZFs/ektX/Tae4JFX9o5w5MxGBrSwIMg
ADDBuxB5Obml6CcUQ6QoBllrUsb8iTUg73rmkcxfCpgJiBEO81/7pR5Aj9QLOvPS
/ZaL1hmxmEn+CigOUf48jlm+MKYcKIzM0JoKhVGLW6I+G4sH6amfhXjP6tER8nbX
3mQeF/08YspBQ5o6/lokRLXqWHJFFg/Ru8DIZa35+8ETC+agDqJrOKNgFw7z6zIn
4DSL425nMeBcWDcVbIjif9OjJDmtBkTZ9XXCTQUYi4AGVgN1vwzUQrzE4XNyaPXz
AR3meppQ+5Jf7DMGeyBs7JmDo/ZOg7NKwgyHfNeDU7maQ30TwrXxXrAqKjHw88hn
JIQOWt9HtcEPYc0gqPsNxQdXf8GAW7S9F3h0hUHaAstTyl0nzeGCttgFgulQiT3s
ubkwmzf3WQIIlxpvtzclodDIryFPaQx+kn43z9LdHXpacdCdrBGZFZ18BPNam3VB
RiU/M9GCxhTA9harKPdh8YaW44pVC92unnuEmGj7sD9R/MCZxGrIxhT+bf4cNcpn
dwHG0XX5SWAM94P8jnvOMlX/VPnGxEoC1qMg9BO+lsykUozIuxCQaz7FTONry/dt
ncYJNS1q90ldI+uAZaxGZkRFNTlfDYOb3HBCkpsvyQMFBXeZlpjTES1YSfLpEIo1
CjuQX9AMaZJFpkHkIs1Ly1cOhRyq1cmUcN7YxED+ewD1j0LYEn5MrmucE9xeDX8d
x1XoXRrScyiAZajhRva8S0e6EbTvCRasdtd6VLgqJpzE70/v9PAG3uf5HyzwicvZ
cYtV5NgcmWhQTWBQINIWm7mi7lBsnaAng52+a5ffCCqRDQZBb67mrWwwv2D2+snB
PvIqI9Url40hXAqVKtci99EU47tUuv89aK7FkZ0pZVnjkL6jcypm/lWFbsXzwB2E
6F28cyM50WMCxEId7c3sDSYve9SsV4YUuy6KzRWG7DNaMMp1uXn6L4UUXIeYJuew
7K3fxQVI5LReLi31+X9qN/8hBKHT6qdourLh7AoNR6LEyzL5N53fwto7E6rhQlfb
dGdGErWtFx3nelN73QLrnaR+IRqT/vF/gC3c+lzcONFUTd1Nywhl8QbZtBrd6HyJ
GpVyy2WxD+EWjiDcSX4r+XccTHJadaPSymCkTpjRpZHgUq5HVwqanLIc5iZykw95
6hZxJXpFxjfQnlW4QxVPTJ5PUMVZaFAqhUJK0vXhxzB46n7TnTU+3mYh+4Ns0YUH
r5v79Ry/An3c6gY87IRWF+dKagrqZWUABecNLbCJte6AdWu7HmqjeWG/P0bbjxs8
amsjaDwlSEDdKqByNeJKibsgh3YHgdneWhmYSWFvieHb6oAs9wDPk9sTAdbCP6Ad
EizlrcEvQ5CjKAkUx+2ANkVGoT9IqBgHW3hU3OXxewOzhEthHtsEOVJNyHmZWCS9
wqFQSd6j2Yf32BKx1ddHT3I3N5EhyqzpYBzlytpin/tn78k+wUKT4R1nrOAac4TM
rkfnWNdxLNCOiF3R9yeXySMixWsczM+KqSTkc1mAEvuaTDDLZu62m9v8SptriKOC
NYdYY1V3nhHaMaaTuQLN2FP6WyOMeQfZizKRpAb9KcNaPRy4qkRBprlnO7CB9Wxl
Dbga715OPhutBtOJRc2MEHwV9JUIUfBqllPg3zVEDQno0Bdp6h+6xSdDJuqP1hZ1
BoK6SIadtwCy35GjzWcEGS3lb4iO+NqM09LSAEqEt7jz0BRgD2CjYemWMcV16RTn
REsS/C6WkNJ29+r/vabr9hzPpWNaXQrWXqQ1bdnhQn/K2MuG1+0xbb4Jdcb18+1Q
TLvlzftL7u1ina2fxAD7rnD6vvsFVC8MYg/NcCK5DqqgOfUPpZUWp1G8c0M48ShT
mTJKEgWbVQWTsTDsQTAS4l16GPfshT0RuEXjq3/qVM2yqLRhBkPMtxzTZFPrhuBt
GcV6Wp85fEIKGi6Lo8d97z/Fc06AJr2JbL+XPnXlsxnvVJ69VZQFQQuG+DH4czaB
zakAC718FJ5X0tOws0NU8BHRphXPeiLHJH511Ucw27WvtQ9/O65yba1kom2Rstot
VVECk8gjUstegzBVtvdzebkX6CBO2veiowlQ1s1XxuhwwqeKwlxE+wF5X5z9s305
d96O6voNPdZaGpDyQYQ6hfnwzWzD6idkqMQn1G9xw2sCrmJfGi094a4f1ayTGZwh
fiJW2+15D0h92Ealdi6g68aRNnfTKEJ4NpxqSxV6VFVajUSxv2F34svOBwrhym3j
9wyD/GgcEwh1o9AyuxDAh9u8VKOZouQcbtcJT+/YDlDgUjIwJr1vh1e1tLylR4pd
eyJWpSm72qssypJi2Krk1mycABCjoD6jFjGs/Mjk/1I1WbVY6XmJ659RShaqWDko
o+1IcSWke+GD9BPxGDBrEyJCz/SNUuK3Rvwz0I6QaOweAxI9iFYnzY4MBbRJItKS
RpQK3hBEf1mt3vW3GI+TRahaRqUThoTq0kgjEYAVvCSorQZBN0kpL9ewZGUEEeZM
2UFao3t5AmjcgLHHTUi0GHB/pXRHDBaugEK2g2519N4iDAStL9rdJdnYS+jBOSn7
xr0U435P1wW0fcvp+cL6ThDsaeVilmmrTKC20CAZJ3Y6FnOVh4cT+sy649dSsHYS
1EsnvU3oCimMjLlScjBSCu8fhCrrkjzOmDU/OG5cQ2SwuBRqLPuu18hKrkz+PVH1
7mdtOxwY2Z5QZv6ChRXHcij+MIVvdU2AhGgFje0r3vdVVtzS9ATJ3DFLpTT7+7q7
bYHNEALFQr9rAxgZJFZqd+iKkuyPGVjSC6UAfGVwDlqOh0bi6hAeJgil1s4Gi866
bjsqaFjv4txx0fmYTTRXstW5sgRKHohlumlanwvvLp3gRBNkTw2KhOb+Nl/StPRC
Z5zCvRrppm7VOc8ZGA83r2m4V5jMY8XVgLNGk4mUGRakFGZFnCzOqoatE83Sm6Za
RnPFV46pIzfcuJvOkY0AjFCwdWmtx65b7xMuuGCMtOW96Nzrdg0JV6v0s1RbT5pK
vk1pN0dtnxKK7svtAtTPNvgfgeuwh1IcZnxZ9F1Mfdai5nDri3oLwM4ZTXvR9ZHO
ATZM+GCyuz8K1zo+t61OG4O5/AXuDuBqZmr6Y195eSJn+qquybJTlFXC5KxE1bSS
0SfIrCNgYDOPdCq6YqNfWzDxOrNRZFrkuouVltqaE7n5oYWSOrPM2EDaxKt4wxJ5
dRxt9PVLWfMV0KZwdnJU7t6O26SqRR3SBrG4zzBj2PrUaZc/1QMfykmTwR/6SyUk
H085XN37A5VBDnNJv4x7AYQx96XGBbqMlw2f3AYTSuZ3xZCwfN4bKu4bhvDPohwz
yR4EltALMNgLk85/ZG5ax/N/MUbRVAaBserO/CEtQ+McJm7wGM1DxylmKmZmMOVl
L4AAFQ1NahkhVA+iJPFdDQlyiwXnimfLPaSEl5Tfu8fod9TFvaSkSFPi++vwajgN
lPV9ONqAJOxES98xDQ/YUnc5g0oMAnn1/EbHp8XjNHApD+AErQ0rW3lqMOBpsiHx
jZUJSOW9Dkxmd7rz8ECjF1iBw0+fySvIn1QxJw3BRiY9XrlSjhNK8dKNyCd4whsE
zHgHY4AWHyUOK5NyS3maWeasfO2HDwIWIX9XK2IaMHFrX/r5cU08nexR5Jm1ZUs5
oZm8XxtfAh0TwvoO3jkAsxcHvwtvsOq46cHn94RUsocwRVrYjT0XSQTrXQfqRvqI
xRrU0E8ObXXKyg414GYsD2nlMcYmx2eDuTJYTp4Qad8kyVCDKVEfPc0YQn5aw/Kj
6ZADG6HpgesDO2VHNyxBiFOoMLkvcOGl96g8ICGjDG0rXePjjQidZ6fURicMKEAB
hBePRtcMDwyioc750Gp6o9FU+voBbh0crf+lrTywtbiMXJTZZM5we/eyvP0CulRh
4j3vrDxvOrTv94en3j7TC4ANKNBEIHiLZc2ymzfIVAgMaNQSOAkmZM/sc+I15gHI
xMTb2RkGxCUcELMMM3dR63bQJjSPgnEdDHYyHOhOCrpitLOx4J5zbaXTx7UAJbU9
MejgdCPDkYMNK5TxR5PqT4XtLQk3WtBv6dGLzdk5CKHcwxyg8KogtlK7dfzaeMt2
iBPX5ele4xHuFcl9DSsMxt5NpsSpz16SIk+CAu94ZnB92+mB4m20RzSUSnggmOlY
AKtEBnWImqNA/J/ckKSJycTIrk3APbJdvldM7UlA9zLOdY1ORDE+Qk7Qp04FrtTY
AlkQyGStHMV50m0J5T0V76LqT5nL3tj0Hq5L6jZYg+YyE4O4oIq6I1Gwa9VcvLZm
ozxK4K3Ky5+80pcj7zCp6rnN107q3w8THee1UcURyQ9D9MenwUtJop3SALfoacW6
4LXJZEqcztr2b1m8XZp964g1P+h90wcT2UmRSsC0H8HLMrx78Il6RMQK/cqDHhqp
U9yUgGUL5rxzVZlMiyWJHixq1yi4grAPuwk3nT4Q45a3rLA5gbyhKzE7AgKA+68q
FL6L7GekVvtkhGVvmAFsELo6j7WtPXvii5WLxYRDXLS7ziB9FkiyWq0ikmJUhrAd
99l0bAh25pnp/t/S7tk10o8Ih5kYkCmh4XX7VDwZyWzBv+jP3QMFhfCo0duj/sL+
SOWKu83x25iwEeJ6T5fudYUt0rgQNTitPRkKQt1ZRZFrQxANhX8uovaZDUphRgGC
M1llcKDDC2tI89rbKkcc8MzBAPjlpb3e2JfQ2Cq81R2mHg48DJ8+bDVepdPVluIR
bIMdbYtJ3NNBw2s8PuSh66DlqSfTZjeQxqGYfsCwnMG1XZ7eJbzlWrexVvkH2sF3
rVMgt61ujO9GI9ZU1F3RH/WKFLspIVtoBP2INLfpxQkcBAzIfSFm1TyHjJNs/lP5
5t6NNN4bBoxikH6z1kedD0SbnHlmjkZ8FmEShPZXqjfp4bhwPg+GP1s3hP20wiya
s9R7ewMykO2UF93pTu3wHmeiPg/sI0hrZ0TUTFlPsPDKOMcehBWW+fSdp7tp+oMz
ZRQcw/kXHr3NyOXtQcPZ8zPtsExiaKXD+S5Xwq3JGUJnMI4lINgLRs4ETfqhwVyY
1pa1gQ/8SJzXs+yqU2IDZBvDNO0T/240B5wsfQEaBf+n9bYMsRI220A47GuWHyVs
mToCEp8cWjrNPNq5P4WR+tVPpGJt6BR7H0lKlI9eHZna0NFxqCsKzVnuNDGIz5g3
R8SqFsArW0EQhtycMhtRJleVAXnk2Qfmj7EHCMS8yLzu49KLa4jGecRCyAdQkrxZ
HkigtdoGbYnnbX2Z+i8xzSI+Gsw/IaT1X39pxO0LKsLCxMjAevn/KetQTeJhyec7
uKJ8Sf2HrJ9mdLlVHNTWY4sKQSetQQgXVHZomfkPbRqMk3+Nl6uZM4A1ltonJ+EN
Z5JH4qmZX+gkpuZTF0HFzyw4JtwiY6XX7O4y0T6fQqSFWu2iORZlo/E0unazgbuP
fDZhJ8TzFicIFIlEhlh9iGfmvPW93soUCVOvc8TdDeI/iOacTzEsYDlR2FqqK6WA
VcfHWye+dXpGhvF7FPtKXg==
`pragma protect end_protected
