// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C6QW3munwD6aSpvmBl2ivwpiqh0mgkHtz4w3nLEVbmJAvP7nRSwMHgua5GXPkala
19Se+CykjhbMz3sBErw4jvPhezqdkMYwOiIUePWY94MlnZI7Ds/4KdK9NRi1arEW
+myUlERLmsWZxjjva322Ox+xjiKYulFxfmMFNkDBABU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12272)
m40s47/Wgs1yYZ6hju1CMJstkLvgyPgJUKy4P6tcs8BtsC4xRu+8S52L2P51m9O2
7ASYtkmISYq9WeMOMAQ8MaL+PAv0dJFdOc+GRaEyZnmmoVgdwnZcnIzX96m2kCpq
K8Q/oAB9R9WUss4IXtuovJO2GOk1dPDpjND4BxH13MnwIj6bJVW5MGexXhLfoyip
Eo150jqdhPJIr8jF+cvupmC2OEcu/g2IkjSiPPUL7GNVMsAL3GzKeEn4mQjnbtc+
xLvtv8yamxbUzGWRYJKhbggsOPPIw2EsRgepLwFcVtf36mL7IUNO7SQpGl0Q737Y
vtc9mm5CtdhnBW+XO0kE0raVbWVJk0kjTawms1dpVXGH3nM3f9QY7nUGbjAE8FCK
vAALRGqGbqtFPvLR2/IR9ZwPzlY96z6uIpuslSbJLcWU1aDChQkBm8d03UtcXYme
EN6PZHbNjUFDxRAhU6++49OmLjRZCDh7OtZQFZ5Eeb7tJst8A4Mwm9OQ+XPcBBZV
xpG6h8xLzQFEkVH8Lwv+hcRvH7iNqphiKm7OQ4F0O68iN8S84prjyxOgTu7gdQh5
ywuts0HaIHU6kMChykwvrxkfHw+qDJouYHeViLOgfntujiyCX/mWyn7Vwgu1DcHW
ou2BCVeQa4XrSG64ut226lEEMuDzVJYPK0u48F88KrKaMyd1/w9ofVKiM9TJ1Izi
WRxIINipFo4j/K4wTMnyN8hjroLApJp1fR8mHck4YdulGbMsPReRhYhTxJyQpHcU
qPpS6czXwq7iJtRNmeS0yGhLI792c5Z+n9swrTYtYfuviJbJSl2yhJDOmCAS3i63
AS23jfFTDQaH+bBQzJJHXv76Kjw+j5aoNGnoC9pSxi68lE9Qb7cI+RYGHWFHx7Vs
9BLI6ZUW7CIr8OhYGL7lT85kAIbYfHBpuZgkXYDK2J2+o+Qjwz7431xxw0ODG43w
oQPBypQZBSheo5CBd2fD8izgsVX1pkogW+JW0aRZ8VrZtpb1OMJOGGtc03twQg5W
ZTUiNiUL8c8XgvDIAjyO/PNlA5+xTN9ftk41X6Uks6Ugj6wTTbNzGocR3OeyXDul
TVZmB4gAAmdM9J/P/IxI8n8rKIXOEiI2VTRF+tW94Rq3a4oZrVVeCAu27muxGGwF
4xB2jQtkOECt15PwtVtI3i/jewqHyPFRdBg0feudrWpHyUp7dHDMi2kshqz1b86/
yXfVooadirnHlghB8pm/wBdvkRpurJ9dFI6Dusv4YgVhT80CO/QJDTQ8imxhCCBm
RCO+7V18YTk3BxmMLSPsEShGwNOqKBWkbkOZdYFXUWjZ6YHravpazn/NXWdXPTkk
E0q4hQO45nSPB6hn7PM9MnW9uPmP4QHwQlef5Rynv66EDDsGryQTtxC8mGc0uimK
8zS0LMN8dacJ3tCGuKY5k7qohd7h//C5e1ANyXwdSkDgpTs7C5UpdDQbAapeYmbh
sndaZ+EcJVBBFvpPBU8iwNrrNtI59nzUWOngbDxQKJcjedfyx4/YIQQpqkMr6Fje
urSDwlJy3TVRfjf9lPTdBxbZc31EPMfus4fhbpjU2FE1ohUGnVVT9CQ37duqQNI4
iBUip8JqGZGuCRm+7GyDPPlU69Ewte0yC0yHc+yNVzROKP1v/uiVGLiF3CFr7235
a3C9aYt0Gti0mOGHMijcT20Eg5hCsnhNYSO0qtq0yU8a4SkiX5kfLLiz1u1IoSLh
D++4E7VIyDNyLk2juIjIm2IR84gzGgwY6K8Bt91jjMCoqbkTMO0o8Jc/8s2vzUX1
Eoa61bRv+K9R8DlVxEoQ88G3YJxGKUxd4UabZrhkTVBd1Rm+5RMFzGNOsjJJ6mQr
zofm3UcUzcS31Xgc4sEaYt8pG2BtJHFFsvuViG7Tgce3iIUs3x302dqVaZV+MqJB
8eNr0OPT+k90rNHAseLRPmvDJd6qz+WcbZaZwAKk9wxIkc0TArfswuZT6NwKAg1L
taRSBqy4XDov6zDFerworfysfoazfpJp5ulOQgr9TjRbmQhIsFwb8qmuj5ikCHGy
c4fisN/aPWiplqmSEsftWkdIn3PGrgqKE7dCOEhcyrxCQuQgEtJ4OmR0jcTssN9u
jLNuFbwg3Q3lSizTa/mK99USRNfDgtHpe57oowsTHgGWdxfFBZLzrABE1TnuXPzk
zMHfDhN5dmE3o8B6nnx63Qims6jPsYcBh/lV8wvH+ugCSquSI9nXkEoK9bbtRu8X
djyGUerjT+WgaHOhjhA6wE0q4Txhqe41ucHqoyGnnYDGc5K1caNdX/5q9/L1uEZ+
2HQA6FPYxGGb9Hh3fPcqNC1kT4U5dgpM1Ct/CowYiLiuR9hV8a99u4HTFyPX77mA
7WuUNq9BXR3ydhJgKlaFIjvNtxiTVX3fONBy1FnyUrqEeIIkVf8NV8Fq+VS+Jnn1
lZQ9oKjuFjx6IM2F1G1/APfj5lYDL9KSBOZMtFEULJbxuha/NImkMLMm4KqjCKX9
MB+A+VpDrzNh4Vix0K5nIW5wmwsJMsXcEqKUFKzE4fkpGNfGhVM/nMxv8CFbs0FK
Hj6unFJktZOq6n5j4cDpkdBWFrr+gpkLorU6bxRhyXYVujHsh1TyIeoE0BrQJ4DP
jcBcFBopTROXQD19H22DkNq6fu4/bgm5r9hSOdJ/IuDLEeN1y5i2Vf/YM7DXSg8D
u8IUaGmtZhixAeKtaLi3a6rjfspIeG4GhiXH7H/bN53zNjEMiWGEFf3u/qO38L8A
dnlBXsj3GVdkLFJH2YaE8MglphIDOySIUfxJbkmfiti/QrF8Uhs+rC54fhToTpbv
+uSUr07U0EBXrnpuzvpAkGzr/PER2SpknYW6pdIxgMgrI43vtH7MAuoNpmTwnumi
bAT4SY+vAnTxynnU0VgQuLjGeNKyt3LG2rqkX0sc2Wi9hsrtf6EAkcIyFLSxPTRN
fhvPxAXm2FF09ClIzdfybNcfsnbxgdFAYwghRwbbt4L6zEWRw68tKSoRCN9tfEXR
t0Xw8OBd9v7kmMn7+clfROYfa7JsJxv4Mhnj51yKlba0/BO/iaBRdtAh8V+IEqms
KwuQPsW4wFBml7sk+11utE1GrHxY/bc6ZW1Utm87BgGxhbpU0Sn/OvjS6+t8Kgvk
glyDo8sg3SRNdEFFbnerJoU9v2WjID8YFzxiUfbOlumwnZ+PvTqyTaqJaWbJnsqb
kMF6thKoJ5iQCbE938PfvpaTSWVNqrHGbFkcg7hCtAQvVMqeAeaezK7TwCMVDYAH
i1PwDEEAdwKJ7J5qKa1r4L0MW+BfkT7qNNPUr8ouqKqIFPphJlHcXoUZoyOWl19D
j/l3hpa7u8Vo2c/inyXOoEMgvGIVtN/7pA1ssMaYPnYGp+1Hrzk5yXaGiXPhUPBW
1urI3NXyVrjCY+q/6wZKFvuggofOEqmsrIPtbZZStrHBJR/fr8AjbiUXA+FWMddu
3XKgvsJOiPZqNzGV9NiNOQCoddAb3ZErbTO5j5+BTeK4PsyOS9dYH2Q7JXWR1w9+
iVQeDwKNPhn5OoTVlYIcfKKjsculZJhEGoLzOGQ2gdfW3Pj3nl5fQttRNCFqAFhs
vtKpKE/cDVdTfxkTEmQe4qv2M7CQojzgKtXpYoUDfRf4JugxnT7Jj/4M9xRvVwXP
67rlvizGR5HqUl7FEY3UyRPCfn7pSwsBsNHgFR729CAJRxaw241gZ1Tek7Csn1Lf
I1iXvc45qdJlAXgfIPxdBd+HFCW1kyW/Uo+oHeEuA6VZphMZcN5yv4PB/0iPHY4j
I77SSWysANy6qXexx1Ljn8NPIIkQrgbi+foBcW6OK1Y+1ZWGAIfOk0bsbibRW/Rb
TNXTSA9pHV1xLwI/3H/DGtmFvhqR5x68ooqh13g8CQLIRoYm3ZUk8AS4IYQjKndb
kL6IQ5yJtXBvRFa2ydcY2LEeIT97z/VAha8xX2fYh1dIacG3zxpKEP//hK8rhnGl
TokEtExMlff5401zOshd3XWxlVPkmMtE2tPvFMhRz86nY7KPdz5D+pnB6qzR4xXx
vezIfxAEhPCBaFvHZW5Iu9topSJ65KA42+A38/aF18CONjGHwKDkJF4NLGemA+P6
UyI52vfk6oNKOWlLv9kz2Qbs8FLx4snr55dy/dg+KJIiDKuZlbZr4yUT4TTFn/MH
psh7+mxJKLnNCidsRnKVH0y9uChk5b2DyNhqIiMWALP/Z6eMwcCAirdKFiB2fwkH
KZ4ss/MxiO6qOrSiZMSwFpVmJSHjuZjH6QNtpDmEJoSgV3PdWnxm4DpYLVvSX0PL
VzyNW8l8POQRpizvcFw5HWi7JlYc+RtkUcJI2aUKCykQJKMuHhtT5T/e7Q7T3kYy
8wmT3juxgN+k4LeR/r/zDZ/KS+hgiD1JE33Qot9OmedWDc3wV3oLIixnrKEn10ks
3tkX6tCdruaKUYt+xacR+De7/KE5JW1RTxolieodM9zeo8eAZ1X4zRCnqvR+vx+u
rdmZxb6wCGxe6EnYe4RCPRVIFtlkSlUMcmQNPm+QM+BSPdBqesgxfmkmSkqY0Uab
YX8rYfQCucXY7DamJpIW/CyXdQRqRTA9p3Ocdc2UeZO17Wmn5B/R9b/+3nkVP/gE
5eQF2e6QJsMiEzzo8dydcVD+P/9dJllMHYw0zKTuI8DeG3CPg/LtOpRxN2cfJNP2
l6zKvzv+7FwuKsqDLqiY7auO/IPZC/mmKgmIMyB+ek8tkmV4yGODFs/bpYgulOwc
gl0mQ7pS9DG3RCwNKqpICTvZCSnGr4vDAEk99ttHEs2ljZdFsruwUcbi61X578Cb
vNpYcki0LzmlkBj6vJHYhdaUzHVoLOgmsoCt5xbZPaVHYUZ4v+z2hV6GwsWEtrWD
T7lyTqAfEoP+ovQOBO0wIfyfSKSZM433R9tpqJprUhfX9/RDOalRNA1rSNK6eB13
RnNZrfzug5JRqS8vhTaqYkxqYRjAEElJQABNb158oYRTJmVpgb1t84FH0cviNrGt
r5nJP7wzo4rPT8Kp4APoC8ivT7eJk+bmQa8kLUQ1jXj4uJcSb1y2UgKV4sTuQeie
DqKoopzhVbkqgUBdf8YilSkkg2Hrqikn1acmeNESAmbx8oiv3e+ZfgvCp0E/PLG4
fZF7exV3IW8o7noFplgG57u/scqN7k1boB3lxrbyjPLq76vguD839vtPRbkJEEpE
c3SMEZF1HnVRWY5eGVDX5Ur81zNva1RsDcLwAQBnK7KPH4z5rQhSmd5Y7lZoU+ar
wp+7uIRe8XPn//Zge5a8TM71o1Fsg1JFzBAvjwdvAHJ+STSUZZOuwMx4evUDZr6J
Z8OGZZmZggxg6P1oESNZc+ydwgeUeusXt1uel3HHPgcF8tkwk981U3ofKpX63FBy
3tiQQo4g0p+2ZxDM/uYHC3M36S7eodpdIOyZQXysT2Ap20KCNc3FqTVjGQZYy5+M
Ebz5f+RyqNQsOcZQ6mLroYIFcfCN8tlBmde5TisZb0NWvMjKTnRW7VnITaeM6plU
ukgBkr/iHxf/pOGUZx6GQbMqeKKLh2vKFk3kRgeAsua+OU83YafoM8p83aJH76RF
wmNhIMmq4cflkNww+wehCWK0W496CNxDJWUOHxavQ1SHS6tCzL6zMyLetVDBpvrj
4Z4MNLkDjnHG0Y3bq6b+lArPuwRpWJ+TfbEAgDoo3NxnCaQrT7jDvkb4SKelkGGg
juemO189vLfrP3jodQZ1A2+sOxCyCRMt0EKij/iLl9st89gl0i15nQVT3bWNfSQR
0OBA85EVcEVsy7tDGHvgQRyeiG4IHkTaQengT3iFIHy9VZOa2LmvG/bAosK2dR40
bntpihTWj6hkxcKoZrO4AjPvdU0P7ZaXKfm7eswtNoQfDwMCnJ1WIu2KXhmg5x7P
AHJ4DeKOejsAvNfNSMQT05vqpwNPAeQy6tx/3wkl7efbQbgu1OP4h2N/E/Bw+cPU
DDUbdz2sMdM1zSM3YmXP9eViSxK/q3BKi/5RB1uKrl18XRoujeAiqM1Exb54KXtB
siTR7jaETf4H/JXIzD0GSPK8RFVJGDcq2E16p5fAeVEtK5m045TON+dU7RUowX0D
Lz/0EClgS94xjxpjezCXMAiJkJNPvN+yLOQ7tN8swOM/x60nrXrGqdb8bKPQHjGx
bnJMqn+O3nUPCY/b/xOL7Kgyu4p/mK7GMylMW/Lgf/qXLh8MiWjf8NlyW5V0S5vj
ocq/EdORUAoWEyoexqkMs+yjNR5yW7rdH08qB//pOLqAjrlJRu6BhlD76W4BH2z2
nDS63qn6XFbx0ZdbDjXA6EXAyCuypeaTjd5S5vDqW7Jfh6IzCHyg1AX82e8owrTk
gOJNKzpobzn8pTVZrYMR9OaRrwKhfWZZeFS7Aheud3eMvMDeK2F+4H8HS1hlJrij
+YQ+ohQNvxmQXzNSwBYWYgJ1i7y6xT3yMGU/TJ5FyAjzkbLhyAZbENvWWXcwwXmp
YBPf2V/iHIsrMZyFNxUbnritvBcU5lxESlm5jsBAOdePibnJOtZ7etfiA79BoARd
WYukidWBNH2p+9Uz/Lr4M31boZ7bHFrwiQD9u4DGboCTfnCF0L8D9xppp5sLg2xv
yum9TUBuGW6VivsqxfHyxlv215u55z7aJSCJwNkxTdA4dgwAVsPMe8lqVHbml6pv
wu+Q/vO5wnBYr7COWHPbd3Ar/zUv9W+KTr7qQjeaf6UmivC8wxssluCmRPc/o80d
afiH/9vi7ykr86AOoxRlCFqxksE39J+dLDLE1kJ5LG1wSWBLZAQIvhz/GYgG/kbI
34fGUs1cJ/qoMTAVQJ4hUI2gPTn/P4tB4Uopb1PPxrnDMtipjiC0Z2gcMR1Ie9DU
wtZOi7GGZGuwM+EVC+p1nngRVAy+XFQMCxeTXahPBPKwhfENuwe+H7xC2+JWqs2u
qOo7fTb3rm6pQibIby1aEPM/mNv8LrEvwKkEeMmdb9pty8Rlmqa3vd1AHz/+yjHX
dsI7fbZ5oAto73gK5qiJyzva9sHueOQFebnZ5a5NBwBE+Z8py8/+yMiU0knuO/j2
Xw1eHzzFevG1BtgZPSJpuk9gaAMmrDK54KSmVeJFQ5bGPrc4MhiAzGz5/cAbS62B
XL8G3kJaPV6e2M5pG/1hCDZ/IBK/Vykvrc8mWWw7X3X5Ul/BftajJaWvVLSmcGK0
ZKXjkBKZRYfZl5goUlpH250BKhlS4CRY47n2exW1Zp4bCbrTEByvSqmEi95RQiTp
ElWUXz0Rlut/L7F6MvhddG92xEvflJmqtkhrX1FQk7JMILUXFlMCHy53oAoRxIkw
ruv0DoncziBXRpsIr8cZsZyz95Y0EHVaLsafjlg2yURB5+YQypCmA91kRMUDVitJ
GMRpnGNN5YQhdGUOlBgcp81g/qn7ETUWZAqJy9AtP/6232cEbrNCdurokTDegh/r
F7ek2jalBhNN+D2euiomIlgY8n1KCcwFvmKz0Y/vYkAzW9FzQ5+4tNuXY7AGr1bg
66AqHtPQMgWVSU7pX8J/QqQBO1KdrRUab82ceeruiW+ngf5Mm8hwhlspjrImUN9P
3CTixoxHrhnZiX7LCAWb0MXjST078ZQHWQ3vRxZU2I19DiohQijmW+SN7Y+fDIIc
LrphkBc92fW/ZbsdVmtCbHYkPKOaesu6u89zntznCpWur/tDC4roLHo25sMfwfpc
XbHYQpIDtMFbn7E29iTcArxHPcDsipG7dSk5TYpIApuQPi3GeofMMtTwImTjtOrX
VY+NVDm3NUwkoCYv7X/x2S5Hrx6Vwg3xjGy8SuR66pYJQzzPOrcvIvQKhnN34gGC
G1P+n2zAlrzUL8Urwn4KlyANpZIXovtHzYNGniDrdqdJHiiSIrbfTZ6fYFirrbUl
dfgWSUTwoqyaSym0oO60pulLs9lTk9JXq4AySVInLVUr4ayVKF50O9qdhXthGpvn
0liAek5BLaZuFO1aGpW73/hPb97TOcTLZCZZZVOVPO6PWk3YPmMTeeM1/qG1qNSz
8FolJgSw8kBV9j+xH1aS/iCZT85wOctGEA3ACGXkkjVZQDCVr3SDEO0PkLVUaYQn
fawiPAtcha9+SgY4aezWEM97FNCLpSIPBy5ayGgdPgWU8QQ7LwBRXiEnrmEobE9R
4cth27ACM/EV21qXekLaDZyO8WVhIilTR5e1myN0AIWTpTygZO9h1rOYo0Sadff8
PQpZ97BW1sb/PuWlYS15mtH/y+/cIeYnQS47hfTW8bxTFIg42LDgTO7AkOga06ex
0/Fa01lK3hisY479+3lBQieRnEJuy7H2py9CP5Vzkhus3ZQRTwFWREEz/fMPCf+x
11uCVBbTiqJEkUyuWO8omECg3iPT6lIrdcuB+OscJOGIGbdZJa0+EdEDLk6GBXdS
QB7a61AW0//W7OUPMxiXVbw3j3nxJ740lalhWn37szI/ciVF251CqYAoncxr6CqE
SED6ROehP6YPUSSeWal5AnqIY3qoAF6VGXFysYZqULmAcI1YXfRsR/61IbDuK070
RvMpS5ngKlzbjwgGsOwmXMmIdT1T7S+bF2oZo9EbQ+sN0ArdS5S6MA1MN3FbwLHm
H0RrvjTHatjQ3p03fXxR3/todS5QSQslmdioA/5gyJE+ytMx8lqd0B9NLsPPJksc
hxf8ly6zORu9/PlUXiXsbVukBC54Ubj1lGlq38hPNsVnRWF6uVocSw7z7fY7KNqp
xOXRPZ306u8/eIjgHdAWGwDzglolpdENq/1Dtz3bykww+49q6Izfd80nsyhPQXPD
JDhgCoSJE35oS6e4Zb0h6fXTDG+ItJfvPXhwC6tO/NiE1LRqsH/QUFAFd/Edv1v7
HKwAAyW6SbvLHnKTYRe2IOyqPd7ku/qHigMzrpCVmEjh5uHmx2W6cFYkgibN3pzx
5bJNXNJqdyL/5SQuwiGDSFY5CekbVdgYkIZONh4qWRp2U16Wlac/evJXM3xVceHu
cj5KaDBy+utRdTNvNd6qI/KA2wyvmkOK3vnJQnF5lfX+8GUxXWWAu9JfzSQxEOoU
LNSZVgvHdvZwYYv997S+wVzUTpPzTiuxvEZ/Ri6CzJnJavfQAqVTT9eheNsEWwXk
GaFy24QmbpUonzR8VDOzv/Vc4R97Uyfbu9TcD5Y1Ge5A/f7Fe7GqW3EspuRPW6ki
q8LO8f6/pf5o7BNXzHeYX+FzrKdLv0JOttrEs+v/gK8qkBGIJsP8LR1bTgKlAJOZ
v+3TRz5fILhBfrM8Q5dpbbBCNceKPGb3a5UzeWkqNnl3NGW240yB7IB/+S+6fyYM
ATpiLALIQYixEckm3BK+il7PqVo6oVSP2PkP+Tq2AsD6ZjO+g09ooBnU56Bn3bl+
GZvfWiy8xi7cwE7No0Odjht1EOc3SmemXmtoR0GHXfyxaYikr8remwV9xVAKs/m+
fKQ0juaXSFhRKpneaBGBBizGOmAaL03PNlurW8A2MPsFWdV/ruSLMIlAhPGkL35w
iNekcjEL1CyX1QfZfIf5DbCuoJ5iYUQvz7cgRSq3vMPbOJ5wsVgG8POu9qhRPIBo
JswJGxUfWuOFlEBDUX9+lu7CDxCL6TrfsoxrISHOQwxlF3wR0WiYnxhe3WPLOm+L
gEHPToussO2d5kK2P7J8JcTy2ABinO5qLtkRUkVNus4uFJZSeFiVRDOdAWouULsl
vxaoj+B9j21bdLgK/G7FlgXtUP4R4fL7/y4zRCfJAdME5yv178eEsUIF8ZZAg+Ad
62iGQxwHq6g1gL0Wr2yu/ZPoqiiaxhRc25ij/KVUR3xRrmGD4fbhpJ5ytQJSy7H+
SdT2BJX5ektHxtyGBi3/iIEqcbU+ptTD3AAsG0BCxvXVLyMbXmYb6whMDr+BNjgt
N6+EVGVHDnb4LlSNHbJfSEe+0BMLTXENgRtb7cYyxbJJ6kNyOv2iRxXLhVeNE5VB
5OPL9NBelB1kmv1Vn9fWOu90QJimJgmOKmfiY+NlMrklxB61Wtd9G7VbzWBVmRYb
w35sp15Ow1o8zsv9xyVLtIQA3PjKIjRcR6GJy2LSc4FfPs42apimpp3JTP1EUjZo
pZ/9noafJgT3zDq8r2wD3+cYdDex1AYRm85TpcrECjVIcNeFVdPxxvCaERSSZkW3
fI44aT5VuHAd5cGP/HkbOStefF8TRfUnpKNS0e8jjWKPfys2irQJzGxrOMkXCg6T
QTc0I3sYpm54ozQI3lXJQYdNgpvV8cx9cjogM8asi14/k9PTKkgx3UmlwIy/Z6cP
pzn108awp8eD62UK+akpGssb+a827E6fKo0y29vHG5/VrO6myPB6ydy8djJ5BrNH
yiNKB+T03KyF1H4y/0tsQM3gUftHOYMYiHoBumORqGgKEL39fTYp+iAidBU9NdnL
zIekJ8o4bFOgurfZoDVSxh7Q06p+Hi7tQo8C49rDTfLCoMsxdeSyZTTXdrYzZYzk
F8ph5JZH6kvossCpKFiYeTLSSYelxhLGGaPDdASNPqAdL9F/7ohawf78Jsv/BNtg
z4g7V1oTKwlsiiMTf43minYqstYXRtOoV+HwjfNwOq8QpMsZFqJ/36VusYeb4aQA
lJTK7hhQhz27kDNEBZy1m1hunLQwy+Xtkhuv2ZYnnFMVC+1Hd1aljBchrsDr5QWC
a+n184X8VwXnZeONgnl0SvQN5NXCqF/yP+DHuF0ACgKBkKCVFw7v3qTcdy5wKxhz
CKz4kpIF8UGVwoaBCX2XErIuKiexeI469xvaruqd6mOPGdxxRHsiFsiJ5Lcqh543
HTKaGkDGpiWyetyK3QTBTNG/yo5J4orBeCmnTnoLy4aPYIFXOjDOS3N5CHRQwB38
pVJSsqiF2ugguVR0PM0orspeHVBO4oczCGeiE6u963kw8TePgUM0oxUtxNMPwv9i
R9ct3foUFacrt1cZmB+LLoKzNuBZFqTo0FSev4lq20RDQeBjKlx4fUiD+XH+l71H
HLbcH1MpVIkHkNsEgVB2pXjmb5vWYJqnwR0oilpeSynXBmIICMrd6pD6oRarAd6U
zImDUOc5lc4eHkHnVDrH7EzI0l3Tw3VC28UF90CI+i0JBCaj4zZ229a0QhgHxljH
WYBbXRah88NKMHbZ1eszmNSv30U4JrQXI6yyXDzNy483BOTgrj1fm0WkIsG7iBw4
1iZO0a5kItDMcKsuB5dpado/4/tzqev6HE/UovKzy4OGKOjkt2vL19pLGBX7heNV
YGH5O9twOHQWf1vbyuKAn57I+dfD+wjaI5SHhgU9q23KjccfE9A8vQq2Err4RZ0p
jTQl4JwO2+fCwtyXWC6js+Z2zM50KWFgXpuKYv4Q1jAX2ig3nXc0/g5r9e8ge0Tq
wcS+lSsMoBK17mpU7O35kFFKBrFT4MTmxnB3zIx72Vw9Aco863CLjV9+7T1ten1C
EuAvuWCrK9N75HjWBNr1U10iLa6rK6bYZmiIIr8KlDoXagXAgVUEJC4vFD/vT4Fg
5C6e2eomS9kaJJAWhch1rU91IxTs5YJGD0xv3HNvuPwRIwqqeU4y2Rfs/ytmGRwQ
2HhFE0xgWCA/lVwGNAte/7m+tHXzsJnjZk6HgsHO2tfVm67gU7XMp3oDvZ4sW0d8
/awjDu99WB7DWLBSelzaE/pyzcykHI3YBgt5hHTOCnChg4Z25tp1OwSmgf8WKlKQ
Yji1zf8VxLKdRjlUiFK7JbNYnXKEn6kmBlZLadYG4Am/jKce/AKRU0CLL205IIL5
orD7dXGS/aIXSbtikCsXhVZxsexxx2xVddsIqm6wKjNaywbnFVsIriPPviJXX1HH
6olOyJCa7KffmS97H39MzDDl5gm+emU5uDiKCt2Muk2novN8OsgSLJsCOkp5FV4X
qslxVrCiiK0hCCwr42KhDYZvgQmluRjxq15oscKXCWmk0im1YmcsPACStTDFhYWD
ty9z1pjiC6szGSfcj6A4Tg88UL0Ljmy+TWFQe7sG5VQdvmnq4FxJCYqFrxWRmnLv
DIKD7AsOOj8MCC2lxqBMa9GtwOkUmy+xzH7QCAywYXWbmDs0lXgHHkV8spmsJ59U
IJd5YEF2yh38XCUYNorXoi41/3+VaObBW8UqFUHMZ+7qnIQZrEEV9Sa1WBb0ZqKf
x9IBxw+hD93zwI+Wi4PEhwMG9QpX7xyhXd2gKfmIZJUPaVEsilMivx02M0BPggN6
tLqoDtmdFH4RfTwfkb4abfj7tbHcbZ94gIsdE6Zg0OHqMI8cYAHGiZ9bYlmzHInM
X2ns8ojj+cPPlN1eqANRMp/RahBs2LtD9zQPTDywMvyZMRgQ3OReHuic0SY0NmiX
TTH1gx+lwiiGPtZ/vNEhpNuuyXnrRifvBwfnOoFlQuae0kvgsWF04c6LQda6MlFm
RKL5EQrfdUotONx835rlnP5MSfJKJvKVaMzAVTDwc87Onr2SarUmwRxj+3MGdOIE
duodaIRS7II8hhd2Fz5XHgjqHE3i9dQpfo12wgOQqZkJdtWGvXLlc3SdasCuqre3
H0KOOO/gve7WS2sxdvBkUaBPFqoExEiS8GLR4U7uOooMf93PpeWdDsODuyqrKSzi
HsLufgpc10N2hOP83ZI6BJVxJjZuinNkS5H4Ps0uiNai2zW3oNLKO6mIVAb0bR/1
wETpkSelEakuFgW9oMwPpDIEqx7eNMjyzZK379GPU/CaGTjjwulQ4mzPzmS1AEWX
ciuBKbK0JXWZqE4AXf4j+jNUrDpo/TS9X76cUW+dQulxl4+svDW1GKjjsZjAGSm5
stpW46CzO/DTbWTHmx47sZPUWWhnG1I+01UUryUfVi9UXrPzdoECvixpuvMdHv76
I+R2g1OsX8zdPGBSaITSSPcrOG1O3qFVn18aHFbXo/T+ktAAhGuk6yh/x2wbP4Jz
IXhPAbSpz49Lm1QZugXy7s2kzhio/YzSYB10eZjiXFTo0ajzbAl2QS/E+SrYi6Fc
vJ28NeYMMHMcopcu1LjMu57Tpcpp2Tc+mvC+j57EN1zeuMmvzJuEEvXC7m98OnP0
dSDMJ4uMcJtKhIIxtLVxDbq+YwNEZ0giyVQrpgF6rxVPMUZtbSNP6EX3hJwj1Xyo
/eGw13e4ApajYC1slnaVmA5EDOgmJmImOMNIqfp9m4NUzui1x1y7m8OV9FiIpCL2
6KrR7UBEFrHB4WZ93nJyyirpRkVxNp1GGsHbqsc+i2Opk1E+c2XfbaCq3j6NPvzC
qGAQ85XY1QGTfwDHTziJaP5dCRJ77BVsgS8Lz7NwmfnBVHhgHpi25efTEtD5U5Mp
0xaoI9FPL/oc2JNbFgIfTr1U4x13kX/2701oTy2IJiN6rT4hoyuHgmkrjoi2X11Z
fWhDmapB2KtrvNiNTt/gGAP3KKDYNdMqfvjYocC72GCFm8YA3Im/WYyCFS5Orvau
07zbw4JdSVIM7a1O8NZtMhSwpqSpimxYsZavbfr57TvVDRsGobMWKW6AS36NG9Vr
WptLmskHb8ZC85qBjvg++GN6WAQKpFN+mKb4RqtbzPmm+ZlS/dVdt7o/zP8tPG6z
9QoOs4okO70u1wRTwRN9bDFg0SyLiVi1/16CulqHS8vdBvNJx8KEXRu1I1YNDTRM
1jJFnpAgJEHOyraebhYAD/5w7t9jdTN6XQ3isKocfo8J/o6Vj+3mtjb81JJcEhJK
Aoohx5EAd87wjZ+Wni6gcpTQo2I3hqvFf3qMszkH6Zes6yBafRT2vMWQs2IR7eg/
qPgVJ86UmboIfK3hxpuC+qXRXx3SJNfT552jAp3ZvqZhyz+U72mpE+Z+XQFdg0Tn
a3R0ViZxoU23Ua8+ktvig4wvbRHIEEWe5GjSrJ6PXl9aV0huyMVxfhbSNJmC3IGA
Olvdg83lrb3lcwvZf9yNetE8ZCcN4RBnRDiOkQ7oWT8gws5r9H0uAq3HngJg3b6E
VI9n4pc57vS2iUxK2u+g6fwTSwOSQheigFNQJrAL30pm+ziAxfjFFvAIGZzZgT0/
hjKpx5/AOnYreYKp+jcdBosEG16yinkX8XCKFAQ/UeO1kqtmOB6+9kglDJKBEZgu
a0DQRBBTW1XKXhOy3iQcYJnoz4rbDtLoI8ldEdgIeaMLbIjg3QWo6B37Cwwfn/UR
X1Dm7tFRsNaZQtt+6DVTaon6Ncp3+OmZtlIwJ0w3ksPkWkial5bUx35EcbsFmLOy
WC6oplPBWQi2I9YAYKdFinru3kPG4naaKT4Fb2UuEBPDn0J5EqTvKI9RX9JFZEuT
YqUKnU1sDloF8W1oVxXaRFvxeyE7pebwq8UuwfYyNzHyDpYb2W4b9xoxzAfiysps
8YjLAV1BX3qsYIR46FL2MfcwChtSUyo93LmK2kCA2I7qdM6kV7T68p2sFHxI1An4
ffBfxlOwgjwAn83K1Bohbggf1l7nwaTihXCyFl89l/+juWFkIdLefpCS2fFL4Bia
7sEZ3iJwt/C2qEykMnMUyhoMdI5D4KnzKUnrDO8rDag5JbjfnfgX/hFYBnyc+7gf
yS0cBxT3wE98PxHfC0PHlXYC0sWGayYWR5EesNr0kH4WE2UBxdMgqrwV5U/ODVIN
D+FEjgt/MtlSOYl+kuPmtqd3aWaEnbvfmMTWfnNtzTmpr1UISJYW8lP3UCtQ+uhe
x6nWAMAeHjdelk0fLQYJlSAf8echGbkQXIK1QU1lsafq2Io3LeTUAd2OoIfTEJYE
DEDReLAXG45l06LM86t3nn9Gi1qCwiJIr9Aq5xQHmiJKdCTyMXTQtUIoV//GF+hZ
MuB+PAkhCWpk52afAEIZPp+93MnXfOr738IEDGMTUMLfOLnGAQ91cWaOg9gmNVdn
I4yHyWgB7u0PRCzXVwRFeWawMhJAMc8roira5eTCaI+PSBSRX3enZaeFHF5wP3Dx
9si8BwIpQ1kBx+Ota98nrWMV3bYIsHcbfPQe1lw6XBA8ImmYLvjM8uUVUQIIH7Ev
epQpSJlQH2JZnJAjH48RQTWx/YntG2mZuTy+bdsvxs5Btaknim0MdWf/U6/A6hax
ZOwZW3H6qjiFPKBJ2aOoe+kY/MKg1sPYj0nC333xaQc6cF0VvuFz2gjXC/AzDEOt
C0pJRpqrhBkXnkVxIDLa2ZwgJiD/0ySEkNVGXTfu4vWBOGQKFD36eeVCFz8TGf0l
U7+zAWIubhsyyA+j1pbVBIEB/oIkRiDeLfFVMLG4rBnoioTLyqjI0a6tiM+Wg7ml
dGaRb2DkrJbnF0GhvvS+X2qYgtLzle6oqV2qKDwatFIKcf1cpKBIrxEYEx2Qekvl
SSxWhTbRrdtVUVOcjl/WV9fq5iVSAMZKZOAfJvradrpiLUEDzSrXuuF1+GQHh/3c
Yzs7E6GNpkklOYJMGduxFah+JFNHeZ+k9o41b2FHqfdGKQ7I288/2WtjOfvqxi2K
qX+WMmhy16Pwb9qyJtyTY++YDeZ9X6r5sogWNYSgvS5+BFsUHrArRjRTcobWXrZo
g5xDXhCJvKfekqf2yEc494vns5efS6W6+/IHXxKmzYvM7iLvya7deiix8Hs6NAZw
DNs7lo7X/DwSDDhQah4yFLd9cHmh0xrmSZ1MLNvR022nUTuIVm3QgVQ8q3txUME8
9TtFaBjJVw1P3gURKJe7wbliNNDI2vBNr2DgxEw37n49Loot9+3Vi56kvpSyy3Rf
JoToSEQd2kwOuifGsXdPAhxcxSme7Y3m0RA9wPIKjU8+5MK23uc/viLEfUaNK1nA
W2hEYHGVRlQXqzV1ZofS7sNQCsed1XxvOrwPX+uX5LArP0Dxp94VBWhftmlrprap
32/AQxxLExym4DFa7EPz+qf8A1E+vvH/YeHdt5qK9xzNKXPxjtdN1mj3h5KgS1hs
j8Hb9YenSHdLRAp6RZU3OA10xakPXWh+XZFrkQbW99WWwvUAng0O5LraUU0xJzPj
4IL31AIuCexaKJBH5BeFILY3egD/8xrrZkW4XgW5A+TxNfbdy4blOYC+PZcUhMNI
zwtZjbRc5M7soJXpOrJnKXlgiD4b7Z9hubaFW4nd0C9e2u5Ks+lMOeuMbMPeTaAz
Guk5X/nH5q9etnEdkpz8PIkQWtvUAau9Z5JUi3ZSUiHxE2XgmIUNxscRKJcXNp2F
6W69lsp9zSr3BgDHoHlDuD3fYgHOe5rY18wZeRfLvUgk3Vw3fsphS/FSlCYZvEK9
zpokRdQLtYdXqpeTz8gAi/RvTKchZrcENnwKsYh2Gzi7vJK9m8Sr39+bJaCQCTLL
fYb2YBvY2gsVh9oIwqi06nT9PinRck9DTer8/s0QEtNa8TtCvkKpjfD/fPu1Azbf
ibzYLEYpxjH7eCBgtigGwTFJH1mgxyxP/c0KlLxYKJQIpHXVlpWw0PaZyn5r3uUN
d5z1mRCN+XdumOt9cnwotu1G+1uOa4GpUZbHQXEBdDs=
`pragma protect end_protected
