// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
haGoFlz8ZUZZMHxtpF32RrTuzF1pDEAfNuqDN2VD7uUhuGByQB6VtH+YpqgO78D0
CrGo9Mn+6hMhaPQR+Bfx3Lc1jZlYlQrkR7CTyFStFSeMpM2rHOqpTnVO1lbQ2zLD
DHRJwKU8EXLg+aB1ujCMRReV0HFZTbOH7huySkdCn7w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10480)
JmQtEjj7GviRJabqVDFnLvRS0xgPtGZo1rZiUEMxtgyj5wxoq6hcVhEX2uNGhPV5
M1KckmJAC8TZbIWNOqK7MbWRkTB8jiV+gnsnYl5NPkD67aHtkyiCU99/8zKn3LGI
TsTe1FmQbKqKwbBlJQDqHqNV3PewidJZ59RCCfyQAf0gB9sN0qhxK3mKxuBrCzWi
XiwqcwwLSbKkzWcIok4q7V5Oc8VJ6gjjQRZcZDnZGwnhiqp51+XQYNs4yZ9n9qMN
+0cmnl7HAsrvAK2tRWqVkq2iyV60oUi2esJvCX/yyftkx6M+qOgAfI/lvNVTMYfd
JdSjELvXW8ftUpeq8iH5+SYg45FWgzPpc9aUBA4FK86cG0GURArW9aPdAyXaqzBY
sLUmW+jE5CUMOlt08/XktGry5z8eeMx//jcEpK0b2kCCRXBBCUA78tANHjmbiVgV
wIl44QP4czc5gnfZMDM5TyWgvRxXQ44fBrJJk2GqdRh6ozPfHo3x5rUm7bztxgyf
3XOq+YIQVBeIW2iwk7b+8W+hT85TUenVV+bDmXEq3rmTA7lR9/4uwDaOJl5IqoDg
WANkMUUOQihL7ynFoNCLIF69zuUPmAIrP9i1tayMiaYXJEBXTK+jDEnGBxkT0XX3
J7CPpaOXpzQcqTGYKCWVN1kQr10KOVPKDN8vUBP0clmstf54M97xz73qZNZHYdJg
0UpLdyVc9zVIKntOQBJJj3/xUu2tbz7kX9ls6rNeFnbo4JfGYJMSPfAkQFqCYHfp
LuTGsyqMtpNQjccvANf6OsU2j9QQmCfqWzDpGH5TPQwwG8wUUUu/4HebDllpAIhJ
mjV9d/eXScVSmg8adEY/3OLZsyDtxjhvb/Ht7kb0LnCW9NT5af6DtvYNdL17JrLF
akRH0rruX7VJBSVAVoZr2tvlaxf9D2sQ0kpyjP3XjifA9giAqkrRJZzzhPLrhtSi
VxCqq89m42syIihqetGMbLBU/PtXGwpQr5P7o/cvWDsJ4PqkZTOykQkyGOzOs0C+
3Em4jMaFUqjqUm5EZDdOyLvoMTmusk+QsXEBLL2edSorWZK9TAJTZxykVG1Vd31e
d9p0hdk1zlFtyHCIPiljcYVANQ3/htWafq0y8Maj3u0poFHIhpLYVRPQgdabuhoN
IijKqhl1iXuNx0cBAwT3riObRXpxNmuIMe3V4Ja75AUM4N/PJsQ/oChGvdmGRk6R
YCKykM21F0O61WjW5SNpxEaH8foOjvak/U6PoJMWw5DrCf1f3qZQAIP2yvtYhcZ7
p8SvPA4wYttXwhuvBZkDljgO+u9cHrvKVxEQikH0Hw0d3KmlY1TCea7aecOcP0gs
76VjZiXBoDk8Pl1bCWdn7Wz//tc9nc04aQ3qJkR+sULOIkdqaL9X4Hbn4fXzr2gq
SfjEMx7c+olgQWeyEMowqVhMfM9Ml8rVIrS5JVUjA9E5P5Yq6l/9bb9GQqjpZ4hp
tfub290jtAK4K7EVpufv/eXE6kyFKpx031u7u6E2aMwA/NAjgoQD96y1nFZyHLa0
GRTSAybNuKvtQQeWxhiy6wD0kw34VCkgAV/cpRhI6VAyaEkKvEAOUwSiMNsbDIsZ
fHGy9Cd5fuJFhbNkCugm9UtiH+Kb0oXtStsU2H/vrnoowDalxvg/YS6yS+THdK3J
B9TGb0b4sA53zH4CO8QXHHpjYCpKRSI4Vp+9qpwTnLmYHUHVJeMhM/X/XtWxyKYY
LZ02yhkwoi45QjhIDJNBgQjfA1NddrYDJZXUtvgI564ugEGKpze2Oc7ZGvKiz+Lo
7muyoEUam2zyWtleYuqB16KwIj/LhXMBEwn1YWHswgd9ExSObHvXeiUFMWvQgVSs
d5zdG2Md/E7n3bOlnQA3p3fy46XhxyL/++zC4wNxxmYujHnkVL1L2nwTLeSAqN/m
hQuRpzrLtOynxoxmDxjN9zo1k4GwlyFnxPDpaV1XMm9EX+gVfUHV1SaRB/hEafAq
0A0irX6DpN6rYsCgjpvnpbBvLP4wq2P+m7LRHnNaH9vXVMKYayvdJuZv6HYS5kDm
dTFygNv6OFbFZQgE8n2Y7Ox7UqzYrMgHKC1vElZn/Il0owtcYX5b+V70G2lSIrlI
zaZYfNpamA0YHxCgLzJ/bq97mGuC8K6H5FcweQ5OJwJRbGNIW5ngUFDUhNMxjzPl
OWtd36TMN8PrJYRCgDZyTSI5XFyH4I8qHWsDHQsznszE+QkbdMgSNger/Q79LQsR
moGbgRe5p5e481oBj0ermouNphtKD/9IP2bgEs7RyNNJJaPcj5hv693jk3hrfNsa
bTw/SfFUU6lu+0W9GB0wG7OHcevvosIR2yc4mzYmy98GflNn8B0yqVxh0SjOH3YH
crlY+vupGCykdAZ9uUEHEBKtwHrz3C5/tQfdqO/4iUeAOOIO6kWzIRg7kbNiUcYH
8ZTZYWyuqLC7NqdQlG3mqEpBXzVxsGOaqEnwUi97ZFWi5gb38seGW0Tw8cYR7yed
mu924Blo8bICDt8sdHee1Yq+4ztvVCv6Ak0E7jMNap+KWYzSPLSgCM6osoVMaufs
hF40pqNlereNfBbOxReReVsfYuGV8xNmHP2htPdIaj3fhNG3nNwW12JsNqyUqNJo
p/oMBaS6LKmRAV9QPyS/VBF9TcsTZzB5EHmzbr1ZECawoq8RfI/OlVGTk/xpB/8/
DZKgG+ez5R/5YDErTHXRJgEON2wvI24rkT7UhR4WdJNVCsTAsQIp5NyvA57WrKmL
L1e45Kj4GzDA1nRs+KVHPIkXoTxf8MX/bOBENnTNnJtQSJt40JmzrIHBpurGsfnW
Kmpb69sCdPduR0UIOpMQcPVVsrRSYYXZbM38mBZzFufl22S7QCw9AP/uWa6DNPmJ
XT+JY1keONceSKA6jkIMjjy4Nfq1iAvNz32y8+keLXPE2O3SIWD/UvbJ8m2LrrTX
fbG4ok1DikQ1zAp1nydMYnGHITjzVjEzDyCHf5SnZlJEWK99kq920XHL53HGteWM
Jcjvb4ow7aVS/N9eOpDAVOnI6lepIbE5O5Oj5LIiuaA4RrLSNd4vqWA6q/4vCAVo
mxI3WaKHyep94mCKFxxLgGYQAf0tdYtSaAYtTJHCAwr0/rNQWiUASX9V4DsvbMrk
IqK3uGUb+AWwW8Ai4ET6C8b5K6b+LDr+jsV7FsRdRIhcPbQc4RNfoXBtQDyaOeXS
1m84Xl9hP1jCCWGKe0ybOvBPHUi90VpSo7QAS9IPynx5GT/XBXNmVYIoEGiQyDqK
COOK6aonj4wQItVb+/D+XZnsfDJAqfpCMDI9pom7taCjkc/nAPHcxDp8wdcPfhY3
rsBFfm2+Y/hQ+5U8IcxSpN7XRGLVJdOQPF2o+vPB4oOi0H5zcx/qAZYtLtUhCrUq
O8RXlf3Rawsv4EbfojL+h3CPfhtjYPze+bEbcGJMdyqOotIQLs/vGNQQSHjKqd1s
tOL5+xySHNNYQYvDmHpClSIVV9YyDC4mhhk0H3guQ2XCwGd9hyeU8V/tPdSrAUdT
EVi32BKrP7wetqAZn48Up+UiFojMjS47jowvtMx50c+95SRFr4qUs5xxtK8FdXoE
KAnxvEwFB/JdCJGxb+iPzhlDFizX+dOeWb67P3hM4QmS9PzVISPVPYJollbfEI9y
IaXC+8hKmH+WstVTgaVuas/RlN/tfCYfnCkSnMMSaIQ/KpJ20bNAFugk8Z1VLK9d
T/Y9ElqnhkTChykwdLNIqQ1PKlDlMwb040iEsU0JH2fHTQN61KxKr1wj5lDs0FQZ
LYHbs3sQqMBtB2pTI0gTYNrJzvkjOPYlP9Kz4bzbYmwYgJUV7CfwmZTdH2dgYjZn
rKj6uoUzCWi+dGJhdQusw+2eMs/G1uj9POuCOwrfUW0fDXvMZAoIXPB+/xW/n36M
fUAXGPmfxE3xupqGCh1ahIzYpFANAYEacFSw5FSAigVg+9oSmjKYi4cKkTKbzVw2
S1VImQUG8gTGhlU4ubR6ftBk54xqzUZvPdl5eLGvv9qJGxzuWjp7M8QG8RGT204S
cQ/RMuud6XGqm6hw0etv/bO+N8R9N5sSI24lRHApV3cW6F5j7zucTmlA33/yjX28
layf00OBonGcykHlz+owhqKDAYwtbl0yiRlCVldmXQQZPkrbEAUt7Hz/jTDJSvYl
c1FY5CK2hM0nnZ6XezV6ivQtLTBvVOKftNDMnFrKV7iskMmNvP2LBeU17oZZaGm5
ef7RJgDG27sPxcW9fwKCyqlc02yylWHtZbCk2TqOFDDPMeRu5JOaJO5xTbaoNX9a
1I98ocBl2KZdBCcl4CSACcd1pvddUOgKy4DEtiriNv1Ax2o928+qPLXiTWn7aWGn
FlKCIgs88o9yrnevwXwxfcPbY7LH3ziXUExoQVpsQ0G1CZssMDG9PnvRc2aZLtp1
+atoprSjl160CEhaRhcKTszqKof6egA4CRxUgWpqRXt1i1TA1jRPQH9EvtZ91qM5
6Z2WNWmQZ3Iud89os74IcaV6g1ElXS4vd7B7DZdfjsU4sv4GsFooMALXc/rK48Bj
ObNGClSs0mePpZ341V1bYWpVXFwl/ZFa0AukwKj7GETPbRzZgad/Hp7McvMACtcc
K7PbTN1BdtQWfJtr1kwoYIN3Rtn8Po+ndIDi3bjCzs8Q3CHcit+9OBsy7yI0WrJZ
D5jk12yM2/5Xx01ne/h/lLydI4R2y//c0UQlBYGsMOBBQnJARy4V6+squbI+Nhgt
HBP4G6eVu3t5CZODVefFDzc18MMEA2QZb+8pGfQ/zbBw8CLhvCH4mDPgD7nOt23M
tTBFPU1Z2tHgvZpjF6N59sZDDIuOm/cOO31bqM8La/DBIauO/OVd/HMsZytXfg+9
lv9gyvbsvMfYhIeB2JeCQNm4vnkFXfSU/uZjCfwG0g1y0zOggQ6y7+GtGEpJydUR
Uvyp8Bnht2YCS9TAJQycb7vXbr2CEW8sa5nD++99/pNrNJ3Fr4hM4RXxvEe5dWcu
XvnWItmsqhzLBT/ymDIThigwho09zToHxZjAovtHDVkC95X4Mqqqc19DRbcLTNGE
sRrc84zbZHtWlAbuB+bH8/dIuCbHrUbxevxGd3HTIDkEBZ/ur1z/i9IDE/Rd6TRF
eOcNcZzLGvp4CLVf6kJCmQetjcKlDhfJcPzPDszN2dCVyzzEYduxU3vH27esAAt1
Z9ItctvrWuBceboagP98BDRJw8vcTwxXiZXBmQxppuPB3xa6QMsH6ijYEcb80/+x
loRX4uyrC9h0lM32xAY+maEuO4NkcivxNWF7ytEc0/iIDye1bnw7joRPOmWri7hQ
R6J7IAaLN+YsW6pjAkji6kD5eZ0YKfL7JfS2bTI3z0x6c/4FIeegi8E41hG/eTmx
oqhSGY42sljSfWwqk2wQD8Vg06Q2mezjjRANtxaJ0r9LZ48RezG8Vud6YsalRafX
8qvJ5JDDlvC888xRIh1WburX1n2NfMs3Pu0Cii1zoMwSmTWb4/dvhnHS677RKPbp
aFlOJ8e7JaA7EOVUFbEfJRa2/mUWO24+cuO9f6yFg6dynAxi9UK4hcO3MLAz/M+T
fPz1dJA+XBvQFfS/yHg8PdJmV3oby5aZiOC/WsBUEhPPq9tswlPllLA6cz0m8h00
awOZqNhFT/W33An9u35/ZY1ccv/+Waay+Eam9ZVUi0OkydKGeaDeNgK69IbkCl1P
B0yhYoORpb91Id7UtKO20Q1KAJRoFJHkuKrCr/Lhjc5pNTU2PGUJgkvciFplcu9i
sAnjU+0AyzCjz0nGal492aR/pUO+EY7YmCm4fSvGSsFxHP1g3raH1snloN6efAya
6ELeNdyZ/EJ/hGMt7K7KHKnTmlfu5tLcDwM4UI7OjjmL1A4yabbNsh8F/1Cm24mG
U+nz8WqNHLMxhdqRKDDCe8wpYO5oBi/uJ5yOEBiqB33LpHSgrdQwUKytAY4fo377
Vkvqb3GXEcW1SOczQpuHs6viX3H8LXjph5H9sbRPjxWVnRTNrr66oYzHPjW0AY7m
Z5ob3nNyibK64P7OmK1ne5G4QQWliuoYTh+txc5ZiDuYot7LQHriWrr+ZtB7zCwU
XsX2MSDTz5TWeS65AVQNG7j0jS6WmEIFctwZ4D70We5e2TxNVXePzJhyESG4pvpJ
BfKNUFKizQBCpY1l5ziIetrFwF03rT03LmHUk5yt86cAYY46otpsfH/A1MNZ6XYO
L9WoQ3r8kZcgrAH6Cp9JWZTzIyc4raB0P+qmckWN+0+vHGYq8xjekiIbVbDKmJ8R
eVOHgx7u5Ms337/RagyF5XDEr88vIcHSjGAeCARwL2cGM2wBIHC1NJZuMk8QgnLX
chrRnSj/i9LXWM9s9zPjEpxUcJTt0pSVsKRgbLKfqdMsduLlb28I8QBi4SeC/JcP
QjlsD+XV7dMUIlcjcbNmhFTcSgfHlQXWdTuHtkOOafZPMD6B4lZEKf88pO07MrMS
fc9FFy50BgZhNOM21Ngyh4e2q+9AY3gAK+jRqrkCM3rtFFMOtDdvesQ32iMkCUXo
aISyCliM2VzB2Hi9OQmexdk5/SMVQxXW5G0MNGI85ebXaiWzV7aCAJKmCXRZhXbN
0Z5UJaz726tFP6adlo0aHa3L0Qs6exziQzhWlYyAQkwR3HF6XO6SDIZQ7yLGKMuD
bXebi4qX9nJMipQPKrWldzA4EX18HnZ6R3Js4hRXUNneoUY3kdxQejyIknNzaSn1
D068rnVXntEBlInWeca4OhUZ2nEHIqEj3AxjN9vKXLeGDI0I7W+wWok9+5JFsINn
2Cp+Q3gWMpUzsUJujpUv0kBxtNTBCjleXYszyELdBjxIErNJs/Io+T2XnTwrUm4/
8SriCCFIkqViSoOQ7E1rxpI7u3fAppKGeRc9hiuLAgii0//qm7W/qYwgevbk0+5i
tWFZRIrMiyDiod3+yXIDpuKnbcV49E3q4d6p2cV5drj8F1o/vbcdYgvQKcVhdinq
G4Xqaoug6vKYcPOlzIIEr1lTakhIgu1chwvToOv5fTt1iFGBj5JSmRGnRRQsVG8g
OiU0/39dGwL6yh9GiplUmqSMfyrqXusGoNI2grW8lVSJ+X8L+ZxtfdxYrGko+49d
2NDY+Z5aKRgcGpSqtQuybHPPCkIZQqxsrfuQ4xpNtZmCqN37F9s/gptGwsOchKo6
WY3oTWs7iEkngy6BjPGVE1ZyzOMJXeKKhmntE4kYr8OMqOMQhjzT6e3JiiC9l/vE
2YqHs8P2TNO5vzqVLV++RIr9+jA+iJD+72HJkQirTvCBr6Sza3NJvmGZstXgYjxX
CC0ZvwPxk6spSVlFucNu0UbbzFooeNgxUbOga0gPPq0PS+o+b6P8kCsdYQEk4BTV
TCpdurMtgIN6tmo59LPBrtFIRjRg2nrGoyLjv6VZ2VxS8DeLiZoLIwEPLxzy421a
BLfaLydI2kbsoaOarXyPQjctmwadBmQhnaA0s+yrqOyndBVSeeRsHJLWmco42UTs
TZsME0aNfReC2bP5GMZRFs5ylI1ygT3Nqd3wwcYls+vpPkovQ5juNdcJ9+Jjusp5
+0G1knyZnFvYeZ5Zyv+sG/G3JeyLGi12Y5Xywl9ltSGfMK8ieRZpHlti4+VymVPv
cYKJV9lE3Ue3toMA+ulbBFL/mX4vXIuHFvli/35NYVuW6RWLw5W1jASaAVk19B7h
+dAFgoFyr6fs1lB4UG1hGB6HSzUcf03O7G6FZd23R/wHHInanAjJ9zNex4Y8FXDe
OJ34TiHgsmi43exNGQGHt1bgHFMu6WVl6XxRAOXNTbkrn3+4dVgrPhHRfq/JtWc4
0qJCcUGLCW1TrmLyahpXu6ImrBhdzYxrddekkAXHVyCxnAzvEE595ebiAw93BKZj
4lQTJA1Vpt3RQZTZR96TBbwkkUxKkV1cB6TKlRCCPR/r8iLst5QnUeAQJhKvMRfK
Xil/GeReQvZ2hutXA0s4b4JClhH/UF0mzUbHmmevbr9Cw7zxGj1EESwZkJzxMS5+
j7xiBhRnFeCIihBeS+qvUYkQgR0pedohPxGBYlLaPxWqaFAb5muCOLifUZoo0RyZ
tq+h9KDoOCn+xgN+Eqk6SBbQIe5OzwXBrjzhL++9sO3CZTqcqhhYTGbeGXgz3TOe
iaItR2CfkBaw6/MqBgmCVmm5kDVAU9L+g01q2b7nQ3LRl6TM5xcSs6SlvPRget1r
fB2RT7wIzA9hpzBO8nWacHv2FsY1/3TmlglAf8RWTDBFltxMezJJfYYXbJ+Mmlm4
sAH/N0Ug5s6/MBiABN6nu2V67bEkkf1yocztY6vdJ9JuJwF6maIY/nYbTG1D5/o3
dkC/FlgMl5Bh1QOnghTHihfDS8L0gGi+cLRXFXuK4pQan+e2uanTy5HA9O+ng3j6
DwDx+yjNYR4LPiOByz5hIelAWcY+jmnSg3/isX4VE9Ao5jqR9CVlHf/yTE6CZQpl
nJvXj0SDoFAiL/bDckPCr9H6TZ3Idq/rq2C3lamYVbVkvBgELrV2Byfn9U04fJqR
8SbMa7X+OHJq77b77llXjHTZ4HK5fdkQfUSPrK9HE2Lpr+fotVYGl46NEDmeTf5b
JknKX/MBWPZr2/V/NVLle77UGeOBKHK1RPnWwV110Ahnn5v/ESwbGYF4AB09vTtV
8Jgfm0yd8PLtzap/jU8XPm8+1v/jpSb9Az7rIlDuOWQY5pjjokdAE9paBj754i+E
uAK2fpZTrVLAEOjhUWMGbzwA7auOBMRxUcbSCLFh+NJTMcgKOwfhATsikdroHMck
BhEMvL3olSiLCrvqfuMavGM/dgNvRev0YH4PK1NP42nyg8AFidtPSZc7lBrpgd0d
CYBdRRHTXykHINYni88c77FJxa24dNV0SiradiW58b5chlFZboqLpD4y4Gf8x/mO
QGyamucNUWdDPW8evxJio4sKmT5o2mXyIqu6ssFtP85oINymiXnCg/UeMhd8JGcf
ef0BC2tdSv5lmagArsjh16aYxEtDXubmBXmyC5Sv1QAGN1vgK85HhWYlaFKBhmpQ
VeyyOffto7BajLZ0SP3pY+TizZKDAXJ9gG/Chh5Lgr55+I8iKaXZVCnniTtOAkjQ
OulNhMcCERvvyMS9DXocMLhF3Qrwuh0ZOKL9u7v0zvHUYHtu+qukgaqGXKXx9r1z
+NmgfFRlVjjJtJmrwI5q9QVdR9Gsxv1Vgj8LbKWqwSaAc5J90GUuc2t3aPBOnHPe
JIT7US1ZSHwxV4pMO4T6DfU76RwGDdn64N+o/P5TV8QZkeLkVaWQOA2swqE+Gnsy
beR1VqGIG983Re6jgze30ogW9Ndzq9zW2pxDRtOJbEgNbW5uqGLZYlub7n6V4pgQ
wuPnqny1M3IultBKb4cICjTa/42Eq00ACj+1QVpONBxPvwkYqciXsgEW4diyE8B2
DvACu2D8Nf2XorjTnBky39O6Q9CY0HyhSvr+81sRbLrDt5ii4UgopJsLnp3/8fAd
AQA5DtcqQAtDuiJ6OuRs2B96fkmqDgYk9TibrjfCG2P88XJABDfeLnWnBu+ctZyy
ZRbAfEcZuiYiTx/S7Hpw/2/0ke7OXPv5Gm2kzP5WM024HAMQ/KdJ7aCZnTv6ZZLD
t1OqIw9rVjd01A6T6HWnq1bc8VjGWKL/JrWJo3vc28QHaXX4s7u+ksQrjAHdgKjm
85AFtubuU2ESv9gEW+rk3inZvp2mgeh/jHtc1vxoH0Xlgx5NiC0GjOu0Z7j2Bj1G
yRZhh+y33rPQnBCRZe3wYB+zTVoqfUdyFeypClRNalsGZwUgtLcT8Sz0o3/DP2vo
zN784RHpMhPmZN2XMoUOLVRFcIx5TvG5rL6vE2rtpPomMolTVtZ5TcqmmIYdF8aB
IHEv6jcTzpogpnLFoR2KJWK7r1qF3mOsvWAtnZEp0QxBzdZb86A4fyjJOP+6aams
T28nNV1s/O6uCcGgYptB/4s5yo4wbuTjP0q4JosuGFHDMDxoJHmPEJJQqfzCWd05
aZ4iZrfDfr6svK4xHygjKpBU+NL1+cZfVnAs1C/JXrfgNWp+YRMMUXVydOQLM3qM
ZZJj0/YTur3+srwtON2lDWnCOn0XZUozdw85FpAWU/0IhANk4DoITrwAdpTL60h1
nZYDRggv37CXbQrevGQqUXEkieDNWo97snBmgbL/BKlmVmBvinolmJJ5+54gBa8N
DE60jJQwK050l7S//r59j9YFvN38ZN97irgfYxUOw6uDrlnINCDcx+qMZY4idg8V
Js/x+8fkfEJgfpYI4fKV5HeaX6FuFnpxLqyIuD5rJ6rC4GJvlFXnAg7zejUSowIR
BI1/nsqpQymxJiZJ4KppfZFrYt/NdKV3yyBCuwjIF9Hikkbpur8TFpRb00QI/LQg
HsmsBpQ66oA3EDQcLlcFYMh8dVxP8UwimEiyi+pBH4Ke7VVdyyYJ2TvudHqcvZKU
VdoFntEx82OF0i0zDTGM21HG29ekwHjyF5dW/t1Bu2UqSke/ZjSl5uNridok32iu
dFjPA8/H5y0/v00AxvnnOkuVEzaqg36ftwkz0d+HZHQc8YkvXzreRmY7aOXZnagA
X3xjtAQ+vKjil/Llz8UlRPfHs6uCksKXUKeE78k+EXgGNMI8Tbaky4WdLoT0AKfk
B37cI0DMhrjdU4xCS2uttx4SkmOFe4m2nVCllB7WYZjmHfCz2OwIxK620gwv707G
r5WkEpTRrlq8xEPTqI3N/jQh/DSJbeos1/BkxvaRQg0GqV2XQX/jdRMnEIsZNDGE
20EcMSeLAAZ3/A2+QsU2J5+n+bmR5ArpBsf0izn5bT2dzVev0cnHcHWholwhQHRn
kgIQ2Yu6xVpwDc7LgvZlP0Ym9lnCPjyN3xZ/sxfSJcplJ3CWOvrGHSONZWQ6FuMf
LzFgp/AWZapUdDSynIFUbAY81Uk+ETrh7ydhcGqEkSeP/WTTgO0rAHLPceUtsEc5
5i3vrNvqjzwa5nCQ+U4G3FhW41jdskRWsA9w3AmXaGTNFLfR7LImUU1UlUCmfrGJ
qYtdF7U0G9HAM5t1yD7mg01XCPAh6kwYezHmn52MdO5uEDfoGQf1x9NToARLxIz1
AVfLxWip8XDs1EQg/P0aFPESGeA5gKuOsKPQeCuk3OuKo0JCHnmg2PvOMC0mS4m4
qvaoyMBGmyTlpRmzrYl93dYBIoF7tQPA9Mq9YDXtAUrwLzeMzVdvJV48XUWEX3MB
jTui5Ac9Jdage3HFhAUuVRjtsyKyauclXhkhlV99i95pyU9eJfWqn/SC2VBLpepX
wkYTHc8h9EuufS06gY+A52Ltewyw/eMx/lGcVDziUMlXt3pb/E46TK8s4+hlPXrr
tH7Bvw0DdhzpsRcK4HBMbQtGhcRxdO9uAEQrEVCXV7QD6zsvcvjH6cRVW9zXGmWf
aEUETGW0e3OGzVnZF1jDjt1f5Ns55HHJ9B81FLIl28RTvv98F3kXL/IVkk5TUyat
agssbk7NbzrN60+//JnxnLEelZG+6hPvN5o/mFEbSB63pGuw9HwA4o/21eWc2/pE
eCXP0mgk6UFfRXnXfCjvVZLq8/nVEyUbn2lGTCwVuWhnQYXrNDTW84YqneyzrS0V
LB2c6eGLdetY6wIkPD/KARe6NrBeABCZyTUnKKFrEs1GWPp4JRff5r6KfBceOeyH
znlydokKSpKURWEuAx0bKZCuYLZ4tHUldZ6P3U8LVy0agQ9Kcr8IBKZGPNRpe8zC
7UPwYhMnnJuVOyqNP+4ffdIGzHYbpd7RZ+lQMwf+nXPJiMXWzzcYoGaVW3CDw1+0
J/7x1njp5dx/IwdzTwNXSC2zl45Loa7N+KqWD6o6+kmv3oFFBBO6gJI3MuFOBSx+
9UCUC4vqrOLqNnbALCdCSO/XoXwwj1YjC1n8iq3+uGxYQcg7U+OvgbQDCMbYoSHM
P56aXFiWXjYbD3Rkc1tbq5ZNNMpCM8bd04HBQz0uzbKvuFzsWAcxyekA4q+12zUY
CFEf8G2wi+Mgww3/KropwnMor8KPq6tbo7ApeXYapfHiMwGBUKpmpor6cQeyJxe6
Q4yL/EPe2BfX5li8wcEpSuel5ikLKwqDAM6medah4tJFAGtz2ez8sl7vQ7nlral+
vW288dKTv2CM2EmEiVZ9pOsRd3jWr0p87Zn3DjHRM8dN/oXCtmVXpWUZKtN7xm2K
ZgpVmE3tz6qA5FxIxteVzOMMqVEhEZI9Amgg5NMS8Nbbhk0yWsbhbdFaRawqu90n
ygImslNLrZ0QuQ/S9D+aUUV3df4r2xxC+l1AoVvndicAeqG39NgNjOW6495HzOic
pHOGVBHecz+alEv0BpA393dMd0/A82oG/9CJaHJUMQ/VqeDwcyDxaRRxOAXh+Poo
iB25lJiueUYMCjfrdisBNCqwqsRHl+YpS6FIvqJaRr/XtdahHTkXeBlJl+S1J1UK
1hgF6gbGdwbmCeLH/s0Xi2K1hQhvGoOckTJwPyNhZ/Ev1SR3UV42VInK9Rkk+8HL
Rgoiq6FmUQUJiyv6y2VQbZNql2FMmv23fCA24zrn1RRp+otQaxXZv9VWztSCniQO
PQv5r3XpxhhVa99WgsrkQkzw9PGJYcQCe6TooAyHASeQsJA4rV40k7F+ORjCsyny
KByVfLKPheeVypQEFFYm/RiTPjZiywP8EcUG9QYg4Z8qe7I8i47qGRWPauwKn9bi
eoqjO5OdcqakxlMKocJyrScVS20rQpnE5lE66KYNJj+YDFJydJBmFoTQIu76ggtm
U/5lym5JrVmVQ4B9rw0o/r/Qylbue2dDBWb4G5OEoW81FEv84DefARVb+aOQt9ir
Z7n73KmqOvA3Jv+i37I3J0P3v13hXY/gL1Vvsq2IVww+z7PqYNZJiWm7IUXThOvV
61SeYpA1izFJywqzZuoBXPyr2v9yWr1MkE57JCTzEHK/XxJ8m16OdEXRV5RXWySt
VZEknivwyRnWjwb/67iFyr/Gyn84jTwm6eTP/whbVsRUKKBpxageP/vXCl4Ijw6Q
PW/6Vff3tfxOtYF4skaR6qk+gxmIGiSIyzJ2pA/SZnZ8ZXnToutWz25l5OLd/sAe
HC5E4g3UovfYhLQ8SJqC2MGV+6IU+cyfprWHZCKMED7dFrFJ+weNH9D0j5hVvDxS
6VQ8SjOHvqQlmY0PgvfEZ1UDCCYzLCKqYcbLJXR5Ngn44j1lJCOMDPR5wXMgfzSX
ZD1F6ctMUtG3zgk+zymZaejFZ5xb8fDPZDqUZcM76hk6NrTrcnD91JiE7sQgWYLH
hL6tAHNU0c9Barn29tu+r/rzITFAhha/38v1LHj/8AS5ZK1uAtN32YMF+nLGJYu1
P6wpkoa0mHQRyJfOMD4q2ISMR1//m339XCzB/qVF0JYLw1zZWM4b2YoC5ZAR7jVM
65PgnSLOge48A4uJDZSmSYDyU7vPI9ud0Ve5+K6gAtAKg7z3n1hOHc2QZi+GpY+D
dLQB/GJ0W0phbIRbNiEznplQe2BkrFkzDGKAfh+NrSIwghoWkEyMhO8SzoEB+mwo
01ixKQ8FU6AlC1XFXZNuYVCesbTGz/5Mf2GOe8veL7aTIPjYhSWlO7TOOPKRbT++
uoWI0TBf/oLriCnsnuO7XSSTep5SdfJJRkxG5VR+F7AUG/GXt5RHYKgzix+pGLLN
6NaHUGk3CrvFN06i0R4FvBbjwJvhVsnri0KBYqSQOrDy/S2YrhdBPkvLclIv6f4g
lCbXcV5B7r1EDeVdVlWWEeLTKSYDHwU/ER1XuGrFVdbPgAHcZ8Boxxcb9eOJeHwh
4IhYSg7QH1UlFLyVCbgCwYQ1zSaOUKo0ucCHag++c7mlrDpyR3os/FXR47upGcdn
2hVY0XXma3TXb0JWfArjz6nqgZauD7Y6Bb0G0mM0+qvBEdFZLBWODeRTJiulKi8r
DRk2k6WFTlp8rxiHpub/SpWjdqFPjT7C8Pn5JpSw8gVYdHtelP6hkLEDKCZcXipM
SaoZt4rsR+QpgWtlpIcRXw==
`pragma protect end_protected
