library ieee;
use ieee.std_logic_1164.all;

entity dac is
end dac;

-- DAC8532

architecture Behavioral of dac is

begin


end Behavioral;

