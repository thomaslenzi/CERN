// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:09 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OeNng7dYyu3IF/TeN0pZ7Nb3amOLkp7UJrXGT/JxcNQ+sM8SC/z2DaM1jwmT9vlO
If7CdceL82QZWAjsdmBHz0EMCC37l54nbuaq5GJWt3+99y8620N97q/fIEYpqnn4
Zte8VREkN+AG8wviVQCelPGIX697zLdIuQeNOoP5kuM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
WM2G3kEP3Pvsjc/IoJYXfFzg76DMOCxYrJbn1FrsaFlh3WWFtYSomwmMJ96uW0qT
6FrE9TBgvR5xbt3rUko7zPclscPx5zzsX4p7ErvZKcAPSlywrxe6r2avpUy0JyEp
n1l2t+YRih7FgZVHy63KQYLbK3xyIe57Pjr4wnleissbwSDRbKjtWMnxpA/CfW7a
kpULhQ0sATcssaBSDuK4HXJNcXCfup+eD7dXuSNi/dYe+YOe4rcrbuM2/67i+05Z
7GKbeav+AThFFOTkv/tuCTR9uMQcz9kb8FptehVIrG5zwXyf53wvakk/fA4+TKG8
bPUirU2b5OeFLWsmYHekTRjFIFotVOrthmZfNHv+Eiaw2xKiskJjgjPkUb1VRdK+
JECyj0G2jYddjvr4VBabKuMYR5IkmfCAzrd7pN5zVb/KPNVDOVNAAlujxZbFxiHx
XEOfGmSL4fpfF3yJbuErmH0FK2kJzaUBe4QzIxNzZBvb/StAzK1y9AMQH5AuLv2L
8P3NneOIdxMvYgNBxCzAhupOfXXWyBQpnmO0vAn+g32cMNxcmiG7mQ9nBazB1/ik
Aa4M6VUF0FS7wWFGQx+PpzHW/GjrZTPK7N8A94DfAikBOdUouOANZNiuUOXo/JAh
XOBxtlyA4+uPxdoqm6Nr1nCJfVbT+SOIDZm1pvN7C1/zP4aMZmnqCowWUshihdHL
c3hXZqc14HX6/cTlW7URBKi/9Tcf13hIKnI4bZCn1Fx/Gjix9Nf6+K14IDVypJMj
s/ruR4NDP7PY2TV6fLIWtxdKIEm1LPAW7eLogCECWq8xn9Q2B+c4m/BfNmiRB/yE
Uo0XNWVaMrSPMTr5nHhJcvR8BEjie76XzPXwDYVXa3uiwLLQPY6DupvSIQSI8oOo
y8OXjFtcPcsH08+3BBCWDxdsQrxcwyB5Ko2dKuGhwd53cAW/ZcqIdITiX/d2UnRh
oyVTeUMXJms9/qoGTfRG7ncW+IPi8/evB3vx8cml25Uvj1NwT5Bb3Z0Ey+ph+s13
+hQeCS4Vim/Mj02WtRzv/WFMFlzjqgBtMGmzhACmRiPg0bxdSQzwWX7l26pe8nsm
gtkMtcdo1POHDtB4N5QuBsLTZiIeQDaA02PuweOGyWzwS72qzILjSW+719a6337E
xPV6FuFdoWqROLfccstMs+TsFdEy4lIpDiz1VsZBmrXhdNgm2mIslpI93fraIhTX
zXj55jx0P/UjAmUjHVyLkIv0AgaoeoMcoFqHTI/DwTM/3Qj3WbZkRxiilGNSqyie
Lfc/nvXXHaktdFIzahxt+U7J758xRsVZEwCiUQ1hXOONIATiTNL1Z2fdyh0UIdTt
cvRCMJ6uNlnpjNuCaDdG8Phqvv92ZhU36lGkM7EF1txbobUWvTHhBSU0PE5Wsnu3
oj2RCynJqhNEOnkJIG9Aw4Qhbe+PchZoMzdCv5t/FZJsxwV6u1EnwLLqL6u01HWs
I4bzhhCEj7zA6uZ4re0oH1skFasmo/YtGxdI8XRJeCYzQQqcLLoNvGU+D/YZvZyP
OFtfIW9LekLw0ifsjuztQpUSMwIFWqQ9asGzt+Zn6m3TbnyaDUPAstWU9cizRnat
GdjsEV1wpOOPF3FfUyo92Mue0alvss7P3pLVDC2hf0C7B0qnULgG3TSnQI0yvApp
52E3DD/8GG8zZEv4K4+gljLvW9e6h4K/CnI6GvqsVWxZ7X9+CuS6dBEBcd6i5jcE
aA8LIgbXLprzxoPqav93W/fFcdICu6/YlBKfRbpxaSxi8+elAQNnfN9WKNocPhcr
Q1h3YMzP0EnSWddFa9dD+QGiF45nMHqju8pGaC/3iYYRGhTxUJDkLC4D43/L9o/q
B3otP4rwKQJ7ZybehnFYG/y1fNZX/fLgtgghZO7vfTGQc7+ULSpCTdNPydx2c0Le
yrOrIC0ELAvQIfOG4LPyBydPrqVKXIOju4wL89n8bjkAWoB2Pm6n/JuEOGxT4l0H
kb2K0MkPjQuX3Ayj0el+H1GoNODpoNlJsSdU0zGWPLnzr4G9maX9dnCfRihImqRC
EIDKq1Ch9KpB+ATr2MkNy+du5R6PkluZ9lv9PAJD5rOHRLJ3UIPfq7d7DFW6Y6nj
c4bX6qIPQcAA+kyJDm9opcQc7wXmVxDXF4QgFckoRaMZ5WG9v9QKWy9Z7Bx1/uWC
bjTt1LEB49AtG0+gHHJ765cx8Avos4Ua5ruVFYiL7z2NbGUYMHBE383j5ZJrKNuR
0J0XB1kso+ZnZNZPl5fSP1OcPoJ7m1SaSjvU9WJtIyqyhMWJBu9tDb1w41imGvAX
GLgpHWxEzYwbQZ1Cw7X4inm2pbs36CIKnxn2z8VCeFyCWFgzZ6CYVgi3BDtRGNq0
xSnNR5KJo5AC0yZ42s2Vpu+UR030RbUo/KLnoopLItxnreLuSZafpJh9dmYTVMCV
qqSx/xGOBEEjhzGRiPBwfU5HqKhJDX1vmEFqWeXBOc5Wlbf91RlWAlBrw3hUer37
ylOyGf7NJt51SnZOM+YfrLRQII+b5k/asoc0potmBypaM1KPWLrgSeXtA1RPGMyn
kzh+nYsxeSbFcXrTPpocAwqMZbzcwlnshmu1eL5m8g/fJbdo+Gt+Pi73reZx+SVd
nOMQqMj1RHo+pnV8d2KU3eLDLX8IIgv7b1QDkVUSeh/JuGeydPBPVwyGH9rK8RuN
DL7QNhQ7yGztFN9PQ4SGl3vhWIMKqIZR4CDkvrejfC6j1gHraTE74JOZo6l++2wD
x7NwBOuUNGta7SAW19kwy+wrsUcsykthS7NVmYyf+OyEDSzcGJvFOCMMZRJAZZ+c
qfe5pR+LyibDi8MWowlACElsjxsIO2iM12IS51VLWjhxhNHpdxlhDgXXxWW+bnrC
4/zpXvVWCFctWuixLM1cT+6YXVUm6/CV+WPhO5KtA6vObqRORVTsuiI7X2ULCHUl
UGo9E+gYdsj/7Cn55sGGxRMvHglIBFnXu3r05ylHBeoxT9Dtd18QrN3quynGu+pK
g6Gh4OwudIddHJ0Y5zv9ZsJ6f7gsvDBGNoceZI4dRBbFzcUVchgvswqkFDi3mvTt
SeuOpITlLgcwCLCRcYx1QSMPKbI3QuQ981moz01d71WPOAMjSpGIRbX7i/UH/96c
zy60XX/GHAMYwStMFFtLr1/7Ow8H55EIUfN5glujxPDJx7TcvVWhEHLZ4U5mm4gx
j0EBseG0x/0oWWM7AA3zcoa6mRFBeV30NJrAQkJl2mH3MSQwbPK+leL7CCQ5bdb5
MG3I5ReGe4dpAsw2hNVAjP0OYbagEodCOHzsodDRCwIErU6QCTGf+6/HOGbL6taa
zi0lBbg6BIpR6+WWOzct5zeGQSO2dwlgE5D8LgDZ4c04f3ono/ZfB02O9i58k8HM
gCUk50CtgZ8ecV87buNfP0ntQa2bXJPPxH7cJu9aL1tpupCbnDPMpoOS+SXf8RMp
icyBoC+di84P9m1tMycLnyUYONyBv1BQB/IlX9M4qii/CZrvIMMxysO2KfmZz3HU
HJ3zYCXXMJ6tF978UbQonjFpNGwOdCBdDM3cg68auz/GE4cy4cIzwFmjUlSdSuAR
Rie4ExmQyl+2H4XghQxjGBiU7tezr2WyhB4/TU3as4kMPZ1SkU40qiAQKSvPpRrV
0rB7FVNYq6OFXBdzd97LnubZKzimz8Pbi4xH68YVwyBcHeirtRXdX8pJwYPPMmP7
7iD7FBaL8M5Z9Nc5mip/HZi2rHgfVOyPcuIdmF5nXfMtHpsi0rd1vN+KbPbaoyb3
9XN9tqlOv1q53bpb2exJoCsNEgslIPsF09+IlErIOJ9E9qDWzP4ZE9C55HV4fVfB
QAa5fmp1lA7T5VHlIlbL5Rlf/e4PlTCgb9FH899LzVNiJEMuuJ1B+g0I5Q+ueQC3
6w6jE5efhRBjDQcOJexrtudD7FDnnId8xiFU9LYkVKpudLi7Xtra8sr8x3Z9E7Ej
f+wcMMTf28/2Pc9O0KW7Si4QUSxDYbqHruD6vdNRZNL6qG3ZavYKCPQRIecqtW1m
YE4AnP9kqB02bcgtQC2GArzlrlVzNtUePwAeVwt6O9krwWL1qt5CZnRRM1x+JKul
VzuUO3cBvf7c4YSwekgPBOt7VdZu8dXyfRVOG5szck4oocyvme0daee7AuFeXhXe
/YoW5ujYfCokuvDa7zrdVwOwYx0NEjhh2cETEW1TyBIlx+5R8PRf1g4mhzIKeAyO
tOzUDIsG8hQ5ap4X03F12TUrID2soFI+eVto4KU8px6IkprqBd1UKPRBEmjRtRv7
ukvlT2J1+GI4A5UEqxw3dhyXDZt7FfLu4illieCW5Np5Fs7fhDG+82UBvzgMkNPC
daYbIxW51UQ4siqAGRqBmBZidJabrFAXxe3sC7J7Mgu531Shxyd5vV5c9n/RFN0q
XR4nrDFENeXjepDY3Wl7vhqlgFepMB0i4YLBsjs6ujI14YXHZKshFf9OPNXkCpJR
0e/vRnqRZrQbML/gfhLsSeMx6B9qYuxgCeQYCqWC5H2ST7ofVN1fkkMoeiDsY+RC
xK2lX5r1dHJS/oq61HUvxyIppVdJr6cZqLH3dmzoLVC4hNZzB1Zvb2ybIvy34d4O
7ODbBu4Na6f6YkNXjl6M5UjUnMPHG6dCRPFNYiwjLbg+l3qcqnj7KRSPLc+eLseF
HEIhD4Fvgl530NzpNoCX8+o9nJ3AasqTAoV05UoCtZWb+AjFtJarnalGZdkYKzjM
id3upNm8ExxayWa+352Wr/TmD7v7alSK6O94TAxhYP/WQ4eUHd6N3jhGV/xAKlEj
MB8cqdMU4k3S7pz7qQFM21q/JFsSRo0jo+oJdeNqI5x8viRCWAyMRMLgMJn4b/JN
vmVT0ysihT3zo/UdfVUkfD0US6obqoSfH44B1mZNgdElcKUPEOI8v3GcwDKoJLXn
8psdDFEZWK6hOFugUkGARoLiIVQofAgVEFqDJUwiL+6lgs6GN94GM4m/Ol4MfXQ4
JY/J/ParwggOx5K5LhDim27eS53J1lfKBdWhxCWbN/K4PfPjvDK6agZgznjZYrE9
LINXMr1mtcz5sDAhusYGLvlnlfBqtJ5FeC3IYwdVbZWGPr0hxYYcjA+BTbkDbUm6
guzgLceFtM4AVvOBXd8QJMCrtKLDHWRa0m5V16KNmeVGzrEcHl0r7f9RBtGlzPza
dtEfpNOp7R5o9rN34Do2cAEokLPzz7ZbKkOM7OJpuyAU0P2sABnArVjVz+e0xKiR
3943cJGzS+YCKOE28+k9H0CRqR7o8+/E9roAcPIF8n5//CRDMwQr8T5ssbhuvoRJ
8t41cAQjxrWZ1puYFY9sn/avi56RIKEb7d/8rvS7lHB9quGwuj5elWduETE1/hIg
ibGM7jFtr91GTR5zVNeKnEbqKrYiQOUvCFAYg9K0iXbaamtFzGaspiZk2aoSuFvU
dCKRMugQZjq2p8ucDdpuvCOSCEe4xLEY5EE8YtN+yR+Zphcb27d/Z5L7HbR2MpWC
LjBFKj0pK8kBs/mI5l2v6Lg3IaVnvyAGvgk0QJxnFPL4GbA0JVewiM8bK9w7I4Rj
Y+vKB6r1dmEnl4aEdUazfNIjO2s9PRR185ms2fTCyqM0dKToJOx86mJtcWJrJy9V
+9srOPPbP+XRrqS+ngRnqXesh+Bct0dlQAUNJVhuR1PxuXzAOtvDXOM+rXUzpjFu
sPAFvYkUuy0VrRUAj+A/O5Czber3q+t+BYHCclbfxVC9F/VuWJhfFQOHFLBusLM8
r4bhVf8nMS78iQkkIODV8gLWdvUiqjiacgTq4dzSWckzABGURwvVJXAqaKdKzdJw
W4hVGUlV+B7JGADKvIKfm+EOo9BpFi6nRWDO6buJVzg2rebJ4bRGJMxUyqpdgjms
NAKq1dwzDGkQ71cknmOJIMLFKw+JvtlO4ACuC4Tw42ySTrPJteMDz9Jo1TCElSCc
9rykah0MkA1SGpjr58pGDRt3p/+12RyMMjgmvEFTPW62Pts41ZpAccqfhJwjC+YH
daHfN64QryRZ6Dtp/WJ02Zr+/klLwvzp3uS4va/3W/GJso98Q4gvz+Iqshulbpt+
r2Jdvy3ZqMGAHBzN+tGNeiTRGzJ5WKWYPXMUvLJgnw1cNELyhEluaV3eDy7/lc1n
gPwoyRgPO4WLPTFsFbU1jQyvk8muM88UiGZxBBp3L3uI9wCHDtCvOE/jAsSsvlx1
G/csIGvmJfZiXR6y7UWVY+ns6gsyb4jBjNKuRoJS1cGqJymFlJWeazDBK2a7AaXu
+fEOGiUlew347y7IfQkV6G5riOm5f3Z5aL6OrbXal1lQy525uwF96zF4rtrXh1QI
FLGKVTFyc8zAFXSkGaMVRUaGQKBAApxBQeIyhVCDy6m03+Qc6ec1sb+XG3fCqYZH
yv9elEawsVWSMahOsAO0lduGqrTw8sA4vH8wq1XY2e3PT94nWWdd4gPAWXlDV2nW
v2HxBHtHy5Lt6+oh0sboPQ97d+Obi5SrM+RZcxGblhtgjdbHgop6X0nYBB5ORn2W
CsHDy5Zc23PtHT0V5wgbtUXVkJdg4UYKmSCZpVK48qiA3Iq3BkkKt/snWHeX7Ft7
d+tP8IP6DNKV9Dlap20EXt2myv5lkgBMDWdTpdgKVMJB3Xhsg0/x5mtKunxbilYs
dOjryrA7NmAaptwUnXbFQ+PR4s4XaDeJkQvmQKC7uudqOQ7DILrUWrYT16WZ9Jd/
9f2BShTkYI/qNBII/yowWXYuyA1VO4TY8FJNL7SBYr3idmpMgIJtM/ih07qys8GF
0k0HHSNm0jwwsN6EYqp0kbYczfvLrNpI5BtmvOuF255qDQGopxnycdSv4+4K/XRs
OjunhyMbEFSMEQHX0YNE48trTVMgm9Yr3KJ+eV1TudrZ9bGQ/qITEvB1ciGt+eJ7
qSSOHRTrL1MjO4d5NdPlwqzMs+OBhLOO674jt5ltOF8jO1K1U3tVhJAC8x2UJfnI
PYPBqITC1YZcmzN040PRTI6JqSJ/++ZmYX6QT982leDc+UDXWHMybn4wzxQG9dXE
nLXi+6T+0EnR1MUd2HPXv5+HBN9qAGW0PPqme0CaOoEXzcoIbPioF0ALOs9Usy5/
qxPadhylBPZE+3bKl2SIRUERhWt0pSk7gjH0+ph0nvsmJB0W4XAVaFV1Ek/YhFGx
+Bv+mX+G/4Ri3Y4W96ls05Loo9WZ2jDZQT1B/WJ5QDPZyExS8ipXkQOQVXc47Dhi
f4WBzt2caniCM+0seJfJ8bc3iWgCyATNZYAgfSYzQQ/9j7p/ulgxHpsGfYNiDuF7
OMaCIvNdrCxBEzaXlv6SeDBTsoUzO9/OA6QLkm4un6U4RNau02ujszHSbxfIVxU2
c5DslCj5UH/9NyCHJ5eUqzhD6TdybQ1AF3COeS3cCphAH60GSCI+6yL9Maosm7yl
AHUTWF+GENeszsSsvYwF5tfZYwoRcrvYoRgMIV+k3CF+j2jpSPogh8bT6+MDA0lQ
9Bg/nlonjqs2F3VBXNG2Qv6ItQnrJnhrqVsFb69NzPD80+CdZcUEb2O1Ti8TOaMO
X6h27kJlX9JGQibCIVIMylRLJFN7pSKpQSnEgnHjUAGdigJr+C5okLfFaa9hvU/0
nXkCEaUDpp+QInHElm+qNkmoIhVqAMZR9ZOMNYtdeFTN6cTpZRzockCqU271bSKM
yXWiBzQxlaQkbNcnG4hJ7YRs4+/FZBZ+MQ3TVNuygZYTKBMmyyIwkSDigjn80yBJ
ggCstk1zmYrW+zAZLH8FT2xjEyF9mbmYvGWGRVFW6jg2OQOvcogiHuBVszrUsIk4
+0Mrp3mw+yA9xJOi1oAEW2lBH96Iuzf03qph08qpcVSWLb2LLFXZpX0YqEMg//2Q
4rl6wR7fdeV5pw1Usc5+iZ0WXVqCJR4h3d4MUPNK4tJLMkdSqJgu8Y6vaxw3kqCE
Tiw78uLbRoRpciyDz2YNuYCtT8ne7hLoyMClGdUmXE1wV53RUz3JDAb8n8uc/JkO
hlR7td472wzt++Fb6BlRfCm0ga5PmGEn537uiSsQUOr5uwP1iH1bsc9zFBRsS3pM
TS6eqG2x4aeaL8D2yIdqnXPEsNHkpupYQsbPfZLJ/+poIzKjVnqb0eAZ7JyUyNLY
xy+njJpTY1i1j1WhNdDmLu8sOt//BzQdD9RhZDo3eZjXKjnamjhg0OLweSkKbrM/
QQPLfvfChGotQucMd8JoRuI9q2HRXQdN1A4DSlABfvtvimZvHBSSn1+C2w+ul9Qf
hSoPDOVzqLEnXpRE5bz0OWOn9lW2bZVn5xegnd4trCY0JV3/kWewO1HKIdcz8lK+
17362xSq2hCmygpCHw6hwt85sTIg6mz5tCMCaT3DTShgeTRSKzSx1yUG4F9l88+2
aClK2ORwZzeYjnKbXHzl9ivlDVRflld94abwHAkm+AFHL4jJ6wYFCVYVGT0FhGA4
jar+XA+7/JXfaF32ScUnsFFDD+puVJ+XC+n967IINTh1LHrQqPoDeMFkHvg0FX9P
/1shZ3I2n+B0YfKAF+FobCRb0/rqsvTOdmdty51/2p42YSEqYpLLV6PKyBZAOh5A
nI5Mcky7CDgby85I+rPLgAqat5IzVCP8zqi7IvmlpsAluZdoW8TjJuLEubRo4s5f
3dElYjakQWfiMFdDMqAkh/nQImqoatb3TMDykk97wZK/xBogoIreYIpKLZG0a40O
/S3TiJQFAiOQEhm0q7HOEu/1CKP7LKmEJD9XWVZi6MRkiwZW0nD237M2oIubX3rx
T1cYe3WdH+v35ZQmL4j8PynMG2i5mTCRHhUX+atBJXHuTx/f8MS99fuFc7ILRCmE
IlSyE9Jg2lf/fhqO/1loVoFrN/XC0Hf5T0ymBfERFsc400ANCIIBkCwiJq8riGzE
jvyfEhLnSzR/PcHZj8pzDJKcieTbOSFpxn/4suuAUhm3RHZvgSD2aU4KdCi98UL6
frsNSSBTIHVZeRzaISL0vO5Zfg1k9pAAVmwJmzeDeZvmrMT5LBq6OZ0jzSWzAVSh
L92MnXDIpe3LNAOE6Oq7DJEgrO7gCbAtGw+8D9poBMyS2aj8kUKVa9V4kXTWlorr
obMtsUez7/VZtercKEUWzaaYyswCf1SCPfoR33f58B0JEuLGmDiPwIGvVnUHsYKp
2A6x1llN18k0sj9bP4MJwhM3f0gcwUBUxD26fk+ke1xWKbjYZ/jQ6VvhCRfcL2JX
5R/u8nSzRDf8CEvjejhu3w66x1Mtm9GnmK9YiFWBL8uvkgjp1L/c0ANHZ6KIdHEm
caKy+HEYeR6daNLVE5VQ+Xd+xX7t5MAanjj/3kBrejQLxIGFbzo1QMlIer+86QTK
qYhDBuuSw3anOJhvo5ksxRhyT23aRfyKl3D+nVDi9DxIL9C/6fw9JmlhqS62ti5y
S67HX6fnYstXSZTX4Ek9kA5PaHZ5yj5MU7WyKD/WiTyX0q1pdVubYES90vRLSy1G
szGpe4dKN+OhbIueO7FyboVaSaMOyD3cBF0xzNLDSXqmD7xqSFaeSRx/lfsyEQTQ
kwG9w4gD1SWtihcAhV7hgB4TztX+M9T49q2zvC66/WDDL01OFbOgaCm/J9Nve4c7
94xF83kUtmme3J1p7jGDB6fTBT9twXawMUWGZFhjxnZlN4QmjSPw/XBcywfaCi5j
RvMei0jhbFLx7TVuRMQWhCxauwfDeLRoXxc3V+CdjIuwBVHEOgZDOouZ9i+7IeGM
8avVtyUvZByKV6qdsOiKQQaxqhmOHsjGrJA6BLBkMcPg7BucbvuuspGcY/abhO7i
jrp9CgtZrQ+OyXWIRiy6isV33bG/lLOK1v/8c4oTy613UZjaXnWhyu5n4zz/JdPd
F0sKUxH6XlpgXbh+hiM5NVbBueyOoNEKU00dgLIaPUDhao2nYVKOHtH8CV8Hgbtt
lQKiUDOERsm56+jXrytAaWuGXHjD/ajVF/iyFZTNMWZR3D/D7YLf7DxQoNiMGluW
kovNbOwV8FQSs1Mavv3+E5Oomq1wMa+eB+a6FzPjGpsxLVjd4te3ODv0TrprW19x
PJojI2MvbwVNYfGx9ffgoPC6+Qij5D/fN6d4E2xQ3rLJGuXcSbsHchWlhjfgpMhm
T/KotKgUUhhLPxf/aUisNLWlERJX4Y+Q2UCJNODVkAdsJgDbwRHW7mw/ynLocO4X
y3L7RAq9BPkcgGjNP0rerTbj7VvsvuIkQ3Oj2Q2Ac69tYk+OYAwIv7NyRPdFumdm
4Z+YlWip1nYXUF7Gj5PJxmTjvkBKcdO5fO7O+nvR656BVghvU8D7tXaP6zbouMOy
47P6o3HKp3t/tRavYinWCVA/z8eMR/pe0Qp3f2JE9cf2ZuMCAzoM/keMifsvb/Q2
ZmtLXtqi1xlbSd0DAHPT09TjLiSuS4aGBZkFAKFEulk3BZ0BO9MVe/hY03Gb+0vb
64LZQ2qYw/bX1avbS6YreQgmkM+ycl7C68+MeIQDpsRMSFuYhuwYEvA0rciHGE7k
CKX/GS2p/+BRKEURV2UOGckl6UB9kHMa36TAdpuJCoPhKZfPuAgqTDoJVVSawPpw
sT9ATk2LQAQ2UBwnhORU8xpHa2/OoANf9jREm5CJuY9o4cb/DMm0QN5xgfSYrKN3
+4phd5UJDgfdod23NO0NDYndfrmkJL3p8sw/obhBole9HlRrSTOs42urCA9QETmp
aQ3vCAGxJ3ebpU/imD546geDYeS5QsAQ8gBJjYIBFd/B1d14GsTx/VP1g5/3i8mH
MQqu4t7iksoT9XCDzAtZ7Hjw1WQoP9K1L6Fe5X4ZUCjxoPVgW04wdmw6dnwWTj0l
6Hzsiah97jzsyHy9eUix+Z4ABD7KIiq8Cv75P3XPIpshZ5pTT//eYWn4GG7+wQHJ
hiEfG538RQm/GFPyadKReWaohji+mIn/wgNidkfMO7oAfVpst+aXUQg5x7Usd4o3
QnCcUNZ6pdze0fXkszjSnvuXcXOAxZh1nPWSA8SMSXwJANLqTxJjOQ7DSAjMWOR/
WZYISF9cAPHSRquak+mP8x98EA1OFrUVd0d8/UN7typPLV4iAiRVvjVJgn7qXusQ
mdsy2siNpnRh6HmapBe0+LLXxPBn+uC+pydPJA+n6ae2cH2VuiITuFTKLTDA7csa
kbR/d/z5TLS2q6Qj0mAM3R3RCf6HVVybTnSf+TQQCf/Yqr5fym2AyAl3wEp5+Beg
xiY8bo/7rpaXxCJtym+AB1UyhsnakICtHYDo726GRCHXNsl2E+GFaRFAlLL/dR7S
L6vrmr6x2eGty0raJqr2MY2ed97WX16veDP4TWZCF82Q3xFZ79tVjxq5LYKnAkfL
BCRZv9kV6vsRWgMD/BSI0VPzpQQO+1eGjsVTO26WwGWq1cKofDaOv3+Z21tgvewJ
GEXyuKJ+Fkr+mxCfFettW4ZMumYnn7YXcOC1lQCYyU1rLVr+NAwR9P93xs9wRZwo
BGvlbCrK2bmxIEcEDVWwyR2PXEqh1EA20C4JQmBpl9xXOSf5xlhmm5e2+aA7spcr
4Az5BzJ7prFOBL0qj52r1gr8KcPIEEJeRVmxM/IAA8JVRABdkP7Rjm/6vQ6xE1/f
27XLTxOtenUgjOByGJI3pqaV9G+7USIZvQNSnWpsJKmFuS9/veVdW8Y/j4FU2qCb
9DiiVKwBEbjIm7hKPnXy+vBklICPZW5kXaT9NUaLQZN6WjlQtxVdZFRrh1HF84uC
HL5uITNzCqZKHbenxg+pY24/09ubbQtefYSehg/4bQCDW66fMrm3uaF0tdh+B012
yoKL/rdcSMrVQyamBOe1h18RuWYKl8waTFok2/DJZDRFUQ6L4qV04Uk4+xulp729
NmCDP2VvAW9c8dpxyv2+fliQuZ+SZuWfJ+1ClTUn7LRVKyekA3PnPCSY3+IjGWOv
PAHa7LgV7zlu2/nYrKt2kndL0n+tqirpgY7jd12lmLNYFuT+iDc8v3qPYYh21TdL
Rka3IXtVeppAWpvTQdQJ2sp0kPtWLExD+KreZ1shAn7l57e5EujsIoIZWUCZfjXM
Q39+RpKJQO5270Y0skONkYxLE9VqkJnDI06s4AihcCDf3SNe4rJFZCKHBmHtIllS
2cVNl/pWZ91PfHnUyXkVHLqjfy/fm2tbQbYc7zTzP7JsagI1sCrdOVkesgFrx28s
P62iwGnPanvYIbXkTCKlzFK1bxVruhI85ao5im36GMj1V0vZyNcj689OVJrWPOeI
12mzCqGFxS4NtK1TD5FzPoUqiXfJMUXanDHGltv/HxZiOkncb+FG2Kn9bLeXFAmW
hhR92p2gWGqjZ4TYd6y15z3k5KZuigIL0ZwbDjx3CD/y5l0uvVcyRSF6IV/dPUOZ
cN2ckujuAc5qGi+lbE3Y9eHC30dZVUqDguq6k+k+U9TvGtzHEYerDLJSwan4mMbf
/stNcE03bXbGqPnEgXcgVM+DEQUcTfR5xCP39hDNNn4AYTybdyYeSgT8gYo9WzoW
6X0uC+8+rbuQUCOgTPbfh9TeUCC8l3iVRALReciy+KqESJCiCBH1TUwNMOv3k0tO
I0XOPDXj8vOVr6N4AdAh+VbI4fmlwasOfHTj/VOu9GZXQgmLIgkM9kZyihZpuzc3
GN5BSqZTm/iuwUP53/uwBHpxg5CJ+nDypqC6eQIFMiUpGZFZs8kmRaAFqoUg74Yy
8E2U8Su+aFlBa2UXu6S8EDdFDMtnKL42K0R8Sb0Fu5MSm25mY8R9dgy5QI7YFi0O
ry59Dwscj9B17lYdJsS14O0664yaNALcsZvXKjPdmS7FeBk14izb1yTPkiyntguK
HfRkhVVpr2VSzNMwFwpdu+zRyB6ESOQ4LxJ/QSJtHGEPArjGvDHJ416xJmYlSHaA
aENHj6XgXLiQ1+lSBTNVi08gwAdmy0pp+dIj7SAgpfnZhVoyrQYrBvLzQkrn0JOv
s5eTUE9nqRkY6uRm0OpEDNr0Kt1YBvK7zKdXB2Jkv4oqSRoPMv6rb6ukDRgtmmBA
7g4SDU2tQg92DhW5cmEs6kj3RdCSWFGVNZ8te7/2JPnt5VXa2oxP4mU4o2TVLgra
166090lcNccJ4NXYrkZx6eBu9IPnGbBmt6CNjrbf1H/mUn8wtaITjUaoDQO3qAtI
lF/eG2eqBA/4L/Nnv6EixJgIyif/FTIFY7kHTVuGrRwuRObhBjPCHGHltsQhMaqc
c1bqVfZt8LW7txYmrzRyeuW7hzljQhOfPfGTMWeMzKv4lg7aQPJcBd8apVrdDhX8
DcsiW7KiMrw1Fy5gtlCzGnnTD92zlbpUZm0DxRVcY2nX3nrTutSytlB09N+jzwwt
w5Iexw+/W69mqyUjpq5eP8+h0mBuTyDjWIGo2Xoz+tV7Z4WMeKrnIvpgAM+Ok0j4
BHIQWNgokI+7uaV59tWLHRFMnD8srUt8Rgqemzucz7gMoGVTw3qysbkGVizQPTzc
plfvIl3iqrHpSddGpH/LMchJnIDIzn4x+9ZAfaYilQywmN+YK75zUoQbrNluUqm1
sXh6PvSfyA0BRR5FoNuJ0lgTErYtLRFxi/GNteG3SvH9G2hYoLyzM5H3yckUgg0R
bP0yg8YsO533nnSeglLCPNPEEcVm4wOoB3qsN5F4J7IJiezBO8LUk82zMeaPVAwq
JdPQMIjVAbnsh/cCfveohUlGQfLmb4Z1d0MCybaK1QzmBfiFJRQTHmzMhqMg8fiv
6/59k16XZE0+QlZ4DMQaqkU/mSH5jT7b0hWwYHKIlKHEHQLl0VDj2vByp4sIteW4
7iTaaXm8aC2rR1Wtj5PFhA+yJS2zqQ1ds9FGPoPqgY7M0VRJKx59aT2ffnqtLjZ1
HR6MVa1/nkJ4vvPj8VkcJPrmZ8Y1jD0pGElh9cdFqIEfuF20z0NEf4VLCNn2NXiM
OF8uApsGOG7iMZsJpHxub9miX5Tb1g5ELZBDBWmRmg4krHgA7KPbgwR38K5zbPsl
A7cdeej2anbRAlkbgXJyCnweIKLgDZScCQTJD1u8xVK8P7c0Zm3czANoVy5kPaQv
pfGmAk5slzwRaqsPhdgb2SNMhVHqplVH0/VEIKuF4vArC90eJILuK3AX4JPdhfH4
JxPdeoaEewnEgnCFCBMMmeqXZGaCEoDajZT5S1HS/K5UedYyOOzPJXFrfT4G/FDF
wQxqL4Yw/0a5FCI5l5M5ZsfE6XDvJFTBomO5BmPQt4oa1s9hGPCOmJNntPdcDJVU
zk7jta/tBZPKgYkRI9pg6W7bOR8RgTFUpTZKG/0a9yHzcehYCfQ61EXSKRrxVjBM
/Qy1zA8YiX+anwipxrMrFW5Fi7CcRgyB0ll7dfTiIjuMOq9ngQllgQ3Ew4vnf20f
5/Ka9QSVBuRLXYel74ePXB2NLGPE/iefrorHxvORNJy3aTcXsAoY3JF9x6SC4Adb
hPeDQHLpZrg17pd2vNkt6iSoYomD15qPAG0KRRXPbDahe2zeVJUN+tiUG3vYikjU
vnyhtAEUsGADxXOmKIPuXOx3KiAjCEls/jdj0bqz1MIfSsTnsGfo7fU6mu0hrYXM
KWNSC78BIGDUUKNv/X+lbgos0g820xbl2bc8RY299x3EJny8tJHhl5sK2E8jm7ec
fvfalxHfNyBjeK2a46zT7IWuEJVAijIemqF71unPxxVRjW8F0/G8laNXtX/zi33r
a05Qy8Sz4ijs1g8lP6QH7bWaZEBqvLVeLMuYsHjJVQuMrfyZ3d81TsdWWyzEeU8e
1e/BLJwsR52xhm0ZyV6EkTVYGTLv4Akkk+XiTo/SY6yMKFvLrqS4PW5Z4i0TGYkL
lByAWjQMhACLTaYT2MbfVBBOOKBPmm45cjeQjzBssXNoUqGxJd9bFV48GaDZ0QQo
pybEgIbHO5v/O9Teyk6AhavR4zYLcuKGfwpBHYPcSPoKf6K6z+iBUlbajkgbn1Py
bJProAJb6iG62Jv9ZUgBmF3br8Ibc6nAfSJrdcnDaUB8jKDny7D4rBHBxmA4xKzB
9p0jDZlGW0O2ydF7DQWruWp45ZW1hTzObSDgWibYV6fOxq9f87bjue6Y5jfxdmgw
1w+a/Fvzx5VuIzKAZZe8iYxgscKFSX37v9wCLWK+6/QAKotenxqMAzMd8aS2AjCb
AsUn2Lfj/l8UUg9jy65OhA/F/K8weV1jNXonm2eLUCmNK5vKGAhvCeXgv/sGfy8X
cUdHDAYMjAX88BOKfhyTJjI97HUq8Y+KdHIzLmbaRS87DUwJKasuz11oEtpbYLat
Arv9KNvbZeYXwUD7k2v6OmBe7laqXQJukjFjhCVhx4jCCSQ4r+NkRLQp5j/Z712L
lf9H7b/0PBNc9vPNYoaT+fDufwh/E7msT25B2K3v92u59ZlEXEq2YZ1K3Us58Qdp
9J9NNAAuU1fdYmH8Jn489bYaWI3VaoiVPEkl6YyKTiTHnYYKuN1fqUGpgg5PHXan
m8/X9pwacMTL2xzYBLo/yza0MczdWTngKATBbOlbHdQWuRGwIB83/n2GN1x0rSTI
I/bO1wqu9uUwNyn1mcSajNVuyXFR/rGDfmyuvOQ3wDZZOqJlRIlrLyQKLXrL8kfL
cyqVyGzINyembW8/0oJ/UTeQRbAXmu4+Lw4j2TukrGaF84v/f7gtnsVjR8XQ5WtR
Cs9LnRS95Uy9BVDcECMKEt6MS6Hxz03iigS5z4HtAAbhzcInHDdEy+GMWC6HUG7f
oskELrH9sJoyf8WA21e1AEHX660XyyC+VqN1sazGchFgIqhRpBojShC6bfFPGJ1Z
I0ZpeBo6jVOF9LpDR6W952l8HUoThm199H8uCMF+4TpSuJKhk9UqXC1qhi20kT+g
qrgLEcBCpjMXrG7luIjaiQiqFYYcVmXvZpbqKjkqyIN73nnQTmFr9ulnTioHZCgZ
tULSbeRkHZfd75jgtGedrHF6XiinukPPyUeDPspGkk+ZPgIBYy93WRbV1diFEDKk
tnjJMHAyhhtOzMKiVxbZcUIlqhfj6w370Ywsw7Ggm72uK50RQvAzNSJtUhLjf93q
rujJWhI3EqlXTHiS1Tq0J5EFAGj7hdONep9kRjclJH60jnJfe3bfslG5Gc6MlK3l
3twWXsBarF/9jaRS7z6F7jl6xDwdRBVOTq+dnnDBHNZ4KOF7QS2odxIt1+8EujkV
fcg3a++TQIVsILm3jykxfXstxc5ov3SIGlidzPi0KLJZMMViRjFOcWhEpX+gzvAo
9XAyOqPCI1GrHflZQF1bCO6TKuJgciQbAMu/f1stu5GGVDcVv0nJN+NLeYalXgmB
N0oiCtDtGLdrhGfpr5l1zvRGGXkfuANVZUgqWYsEyxtxeu4M20TahtfxDZZgRlvf
MIgZuuLr0bD/PMx5jCKAxL67s3lhhwrT/pfAY9QbfIPEZ/3cbWPVMUJZfgBrCitN
dZW+KYibadS3QuDj5jefDODre7iddI+6LssMEBiQrvZ7YKyxQshM/tP6wPyPDmjk
nA9BtTFh3Z/S72x57ZqJAS+pFUO5olg+fWpmYCJta4E+oc47aEnI9TlfQG1VDt/1
9Sr49GSlAhYzYXUoZtSXBzCNVfjEI9DACFlARr/ttcSpWWQej4oZcWpcQ1vTLFdw
UwrU7bGYrGw01HFNOaWN4rFQQ/wvz8BJvK7smEZlo4nnczlZ1WNftYh9cjLJqZbY
J/pwDdIdqParC9K8SZ3rBCNQSTY1uZh9XZw7WITYVfnLUOje+wU3Om4LNDD1/U0z
D9dDEwwcP/yIqQtfEqJklZbCyu1kBAUlU8bV5ZrKRYHcxrxY/yOvo7UZ5S8Bitro
q45bDihg7dg8qNfetjLQNCTpCglT3ZfCeHTinoeIcdmYc2uAhKLzUu+sIhfgs3TL
b+/hx2W6yVR9HtPBW/81iZzjJgo5J1+7ZFW4rUbDnpf47slf6csaMSjIHCfFnsAw
N0pAd5kJ45ruoPcbYePALdYdXrSLK7XUcYwYeNZhaurFGOcqXXYIDjV5nal11cfL
PTaXXEGXhBSVrED++7xFOoeJMKbfg1tPgZXLvmGwYNAJdLHu4Yz8j3IV+zQSYVTp
pMrRvE1EeQr7LAdVIekkRAsGINQxK7Z3w8rrvP9Ev31BPaEVn89Ot2NizjC34EPV
iQsGD7RSAgOCvshijyM4Q5VEZfSLH9i0r8F1JNJT4mMkxKDT+lJZ/rMSFLOcjbVZ
6Wfe0WOW4vTHFZ3fNJ8TLDnE630gNbD0Tvl+uvGsnjNkfU+Lgy7wPZ0SdlcePgNE
FFsTgiK4arjqIMBWOMV6d5MTcowwIvCd4dKPQkXMz7CgEixlj7NHhS6LCrpblsZB
3GUeDy1PU51OvsX4WO8cXQMNCFPw9nxN8iaoFGoukIriR43EEdph25+kYWxP1vdR
4f06jD8prHXRXXc3xbIIB9E6hTMmf/aJcUUQjhCJWWgVOT1aZF8eTCsUG/n6eGIt
zw3tjTIq+xZS9/WVrstcGh2GnuuS/ajzyjPex9WHQkHgyp6GgwJ7PoZ9eEHUV8s9
9KNQVAxf5bvU7tV1kc7VFK+OBtFDN7CDmyFC/5lzwlAumqDJm/jC2mV0vchLRzZa
zA0qpa+BBU4NMXn0FbsYJIquLt6VqssG5fPgzSyWKXK973Srdk2/2R+SaG/vpyQh
J3/5r/N5b0ObnzV3846ljM9EaltuGEINjbjM0xOgs+CeGHVoLvj6XX17K9BPojsB
s+LwdUt8W0lFfiMsvq3luIfvSNyF1+aVkHmXI3hCeHgkOO3ebdVQ8WTs9dRaJ2tD
HWiTjqmu7rHdbPhxLUm1TrqvsgDwHoIhzt0pFPwe3MRLEMt3CVF7SiMO5AnOvb9n
R6vtqvjhuSYFA2w8vb+WCSOKUJexhwzAIhVO9axIR8WlpFLobGKQvdLR/PrrwHF5
ubLKjTvHG6fugWhqT4ZhNZvTX2Epui2LA4H+oJmITJaMooXCtxlW4r3XEyJuXQrb
osVv6gev7ddi7SpT7mCDIm809L5y38x062kQQPf7AzDhhx8t41dGAJa7P3PDM/Ob
ChSAbMsqWM2w89EYLeXQoGvQAhF0UM1WLxX2DmQAC3enpwpCH/1t4ryiwmUD4QjZ
e3Hh1dbixjKOtu4N7CqNzHWPrAtRyEken5vZ3HJamkLMNKKudUlvdwciHEeJe54W
WVILoqJb5jiZuEX6D0QTnNUP5Cs2YuRgXij7zS/4FCGbrpZHTQS3zVCMgakg/BZ8
lkFGm3XYTKsYPG67sAi4iknhyEYtYt507QKYY9uAPFF8briZz094fpKN3Gmvcv2n
BYWWBnh8GLY5z9GWsXpCx94uLNNJUF9wVjdtrQHNz8z0ap1s63KybMTz10n+9y8T
b0tjnfhnywBgR/PVCjxbFR59S/DZal3UUCyfSKt+UXByfRB+Ku7PqB9BgVkoaLKv
i06JqVStPxku1TX9Ea06H51WQlpJal4P47AZqdh3AZXsQ65JyOVr/DriSDLKIkpq
O3ZUiBJHmsvvYAuT0x0wbyU1jURqRPMWHF+rWttPOwe9dxDV1HeGv4jgfm13iqVs
vezC5RAq2nFKd00cpmzwEkJXc/X7ls91xozXpTAq1WaI+1B8ohz8C3br6uz6vOPM
WdhX8c41mmg1X9DAJ6GO0Hz++ohD4gFcoltmoaOUL8kwLtEvhbovP218hlYcNhM5
7yJx+JnlZUlSvXwRT6bcWq+1wkpLewidKRuJC+tZEvJO+0PhC3h3lGr9n08DkPUp
XpNDWDyZemn2kxNv0/xg7NjPI9WZutnjlqmf/i02krflK4fR6oPg2isRg2jcnV1A
nBcQRReQJqaGAs+udegqzLUFXIM7GOjnW0v+9KBGOBIu6b8CHxCb/V9XKhLTo8k+
9thCaQF8D4pcR95xGzO+J/WQoXG9yMFQQb+34jyklu52FCg5sci3X+RJf7yjaFNy
ssoXqrFOVD4W7UOU6DZAAPXBhwhcuDm0ceAFOpDfand3fuXpMz5Msx74QC7xl57X
y15T1YYvs2k1u/gwOX+ZZPKAtJ+No/mUIUpI9ZygFRcmEg+7xAeh4tZ2kwHH9fp1
wUO4AGQl0sIb2jTp6X5x3B4mOw9SqPWHrLEpOh6Ih7SOFg+f9up0eRLtTw2VZZY3
5HfstGLE64sXJIo0oEesbI0YD+NfqcspCuVH7OIenz+CvCBsnVrs4osFrCPU3UVq
zo+ALXxD1Otx7NMVZCaxYCwosoGk7HZR9b1arZWoCiME4+SfpOYfbq+gshB6EeG1
G2DEmXfOSuqQwykxyWUIjMod92nlyQSKiS70LzG9M2btI5hjSrv6Mocb78D8ZXdm
Q+/D9Y6KEDpsz8UJi9OP7oWYUpzCzo3zxsnQPOFkBS8qD3oqnEp4OprXjGNWBa+X
g6QOTDm+WYpcEJckvUzAmVxlOQrhbDLdrOQt+mlNoBFsdKOrgCM+lcx/LwgXJ+Bq
EGNrGtxrL2X3chJtOQVQDYNnm2onuLTpRqXmelH/1orwkzp/AOWDiLXdI1UStye4
Eh+AySOYpr26VNMYrcr3u7wByl0Ly8g4o+rKlHzIW8ySbKS4KN4mTsSfJhbg8l+2
Gr1T/omff7/6QESEhk7JyDmaDYDwFS/D5o+06W2fheNXrzv9Ug8okRQfxHSiuoqe
4mX6M06wcD/tG2MOdIpWyrM2Cd69vjD1zM1Q6ox7SRb3dfbR20kaUa9uw5BjzeHO
gYSXmbT4x79NAeaOSgHdVE1mP3kQrpu6KcDcqivhZMPd0UaSaOeJvYJTyLxnE5/o
h2JejF4STlK2PvIJcJWw74Lm1fZVtmPO/QDrtosCYyxrHjQLh6KEW4FEFUGAr0nB
IlUBhPbfy9WxqWh2h8y0EvcZqL+49Md7uhPyKTbKM5PxOaY/BsvshnMwCexZDxy8
dD3CFT4iZY2sIuLXEf4SAXrUwo5epF0CMsqN5nr7D62+1tuwzoJSxHEArN4hdxqg
4l1o+pMk9XP44zVe9+SO9X8QgY7md5bG/MGMJL6CJXDuucDxmqwf6MWv9kwQXNLA
72oeLI1FN9qoguEhQqTnAfmhOgK8p2wyP8N9vdZ0nkYeHSeHl7UqpAa5qnzQEJDa
1q8nueLHcYOmVWqQpNGQs09OOHCu7CKPGOhQIMXfLK4tFaZ+c2kPBupFTH1voIAM
7wJMEA+cg1ZInB6/D0SckGa49sF94elOiFkzU0wyA26FrceJ1y+Hli4fQVCXe/lq
3WCUdbtoIascF3zVYh2+yunMawWq8hm2YTSU/61D4sCUSXANa8r5ZOmu5dIxT9dL
C+EcYqJoeVyUzLEm05Kja4wECA/LMIrVBpADfndycxZWRiPIw5C7f87M4CoL2rlZ
ZH9ZGoj3kawkDLgIxHd1LHsltazjyapb2Jg9VarRFL+njCqjHCc/sa+NQEpMhXAl
LapwCYvj1YfKurm9cx2PDmjBezcQo5dcLI1YBQvViWKQig0+hmKCqCyUR+Ox5cyg
weQfKdI2YpBwinAidFfepe+SfqcsYx4twAX+BJxER7rfmCzZ5l58oVYnmz1r3hQW
SxEnB1gMaFrDNzeogfD9Ha8JlcuQfkolsmJ9VNxFnauBjlqQDGAEVkimHWQUKvCM
ZClX3WLUTobKksiZhDEecR9X+1/xAFFzSRfklcJkLNNc78tZSjnJsszpZeW4c984
bz1OFU0vCromHS2y+1AZR8sI8e66LXvVpf9fodCPjOyAb/BLv49oB82wg8V4S4VL
xk421fw3USgwGf3mnZYztqXMzSoITHrgkyUXE+P9K2mBT4HaQ648xBaEloPwFDyj
0aGfXBVycVmbezpKJtdqWfXRwvyOTle3fKi6NiEf2xoAPj97pEnj2u9yjTQV2M5H
qTaFHH0CjpJW2QFvouPbPcf3ocNMhNcHEZMtQEJqEAYliXx9GLy4uMMD4l+J/W3x
nBmhKf6wsC2jRsQNLGLY/J1lRU9qCF4nrjSzX35m8aQ6NHJbTAdtb74Xau0mtRUB
oBkiy/Z47psZ5M5pkWHpy7eu2oYpyn6aiobO2Vqu5/Ng4VEpxoxXpuJMZAgnrYCy
CtOl6sUNGZVjktAtbco1WIWHvsu8pp9wRYvorSkncfxRKwRU2kwvTeEF5dfDrrCe
qvPt+n44mOnMmjH0BxD30HEddtxwrbvUYoqsgMnR+F1pNenCKICLFu0SSTB+yEjo
PZuNLE2lEgV02jvE9PhoFpkfKoo+R+TPSDiyFoEIEiiIQ0dY9P9KgpHkQzpVDygC
/MW4S+WVkBjRalDMRjELPnGz7RT5N+pMSJ6AsuqfYIU83ZgMyTFGesJT7xvVtin9
j/Es5LOcCF9YGpWY3LtCiIOZpJTCxWNTwsV8ubEXQTFks0ngM0aSOD2RzM/8AYBj
uDfYEdSsl2ARdxn3swQLMXQRtgHQqmIxdgpKU9Y8kJ7+WWpq5aig+RBTxmeKZJsm
ulxwkV9Q/ZuLugMUwTwYhrt3SNahd59QuSHXXySA2y5/nIkZMvDHvqEPIzHhyo1P
C3iNLyPaqGxbPJSlTvFWL3OjbxYMnfhwNJQ91ySArM2Buszk72w8MfpYBwU7SsAd
ufS0P/MUGlgDDc2Dx5YBmm4AEBCNJr989auC4zPtj6ldWRI/tpmUlJjq+18rXIDP
F/dJFSJEo4JHIPCObf2IwLkbMygtSVXynr/4ImC7mMWvMRRBcXjG1fw2b1VAFFMU
1nzEnY7zEodGgsUq0F26P/bAHhQ2xoUxb9N2QnaYWsqx5Hf4Ov1yRVPMbForMoVV
QhXCIBEmCrEJhb0f6N3+t1BcUhqr+cWKTG14G/JUHBqTHOPic/NnFHw1ZHRdyR1+
9Tl138XnXF54wVtu+HiDd3zUO9ObfhgE/gJuW1xAyFxrxP80zf0hyugwVw0NJoRc
rrM85qPq48DLUz4QL8/tiHGJ2W4tClahLEqALU+FEUR7THMzCc29oEgLvjBE40HK
uixl7DdzG2mdMDtJ70fGgG6h4Q/rkSsq4Dk8ZimGOI3unoEUlC4yz5uvxe3k1CBf
bxgiqt7DWrrXkj7ofVGgzeBNgcFPo/CTyAkXKPpOR8d3Hup0GpVuSFco50mT8f6u
O4LCEZPuaZMvhUMrEuJ/Q8sLq7Gp3SbQfZgWwS7KgSZ/m7sTSpQKBy75o2sH1rwv
HJoQL8TgTmFs3wTPTO/s2l3DCo9F7MUWSj7Y2KS8LjjUMEaTHMyywjW7DEwxU7//
FKc1dFdcZTSePIp4yU9srm/O0ZpY243oNc0whTPv2g5qQkPk6jUCZeUQqgQ+LKnh
mMpt5yzdoSos89PjKu464L/RlnMtW4Y2lZBmKHAGQrGHOs1qOdizY7ficyHXhPbk
/g5W7xxdyU9QMhziLd72QSXYXjdHX+f+fbQxf8jQ2o4yPwwDeDYO+AMJ8weUcLYQ
7HMgJmkysIpVUZCNE1VIUp3r+9IzHJtdBo92spVkuYDBpDl+H86K2ypI1lUoCRl7
IlO6zkgfETVUIXPCZam2xmMHMEp8Uqvvo5LUtjkKOe4h4G2qNfF+RGSO6/ThlGSz
2yP0MnYEwwpS+z3yfWnty5rCko6OA6YTXVtuuYJpaBVRLsuYFgq5XqUONApQYkxW
aW9ilizaP1IA37EBq11uIMottTo/8prH3w/8+qzqJbH1RsniYckUp/1zWo5vdUS4
fP5QCe3DA2UKrfQb6ae5xq16mYk6MIXmbdA5KbhvaxPWISOtws0HJgh7suRmMTLr
Qn0o4O4qyAB6uK/1HUtReFCoMSjb1nNIiS1C5jlXCGGOD71zVGeVuRQ0FIxrztzS
cXpCS2mEK+Do26/qjweh9HxQPQgzdE9Rd3YnORSDC5A9t8PMuchla+FFR9m7d8pW
NThkyugWtin1y5ubiFvw4TLU2qbF9CbCWgfuUHoCjByiHeE+Dz0Hq0hriFWctalG
mLgFPgQBXC56D8Ik303Isv5KRN1k9Aoeiy9t5M2UeMG+lzIEbZ4mebvdzFAncupb
UhB5NfiF/WOZ9TPfBDtdJ9fRA0iJlvlNmHH28K7Dz/1KaoZ7tCwzJbDxn5Babgpe
lTu/wI8fRBMxqOAZg2J2lT5RzhUwx3Fa20rL1cT2q2Ey7ZYq2G4X8lBUZi8/eUbI
l7Dout7qQm2rxX+SEdqlT53hl9bRYL5uFaT8hcymfoq64PRttHfcFBodBslLgQIJ
75QAYR8BrmxpUQYvMDTKjqHr+U8Ub3A9jwnCZimZeZS46jeSlp/8IUuo9wAzYKQW
vARUIFeQ9oWA7EfscHHYqP0D2We6XB3zP5LXqfOPkaNwhQ1PhWJn3BpOhxCIol4+
2b4HWcG51iCPRUpIufOTEIVhSRJwZ1Rh6n/gW8ZyyllR3i6i1++STSs1NlvhjxwZ
2gBS5KzOUcffz5yDcNMGZQ4noRm7K7zGQkyh3tIJAz3PRkc7WuE0eGmGvrbMqZBA
jReOOmC6aeQRPj58XjMzJDwwVlH8qtXCVR49gsGVWIH5aTk+rrIkJhWIvHpeH+SC
Zm/HdUvWKVy51NPV5z9/Eu1xlg2TyD93nSCt7vUWhvoShfQDxZtPTyvZ9ek6rsfO
pJkqGNyeH60FXZxddEsbLHnluKcGlNyYkvV4MdYy0kmvCD36FeXIkY5XcOE071+T
Au/0gQRzdqKc/dv9koiNPXlIp/BzD+xmAFBPYw9NfMqiTMrakCq/i7pjf/2fKKSV
rggKiUtg1K019CbaYbeRSZBStrmYUmkQfvtr7zsyR54dYJ47SKmlYj5snFL9+OQK
h1rd+KdhiMQBuX3kpQFZGmbvW9q/PmN8qIsCxkXzAv1LCJBsLZowLQmkSV/JX66H
IFy3d2tJlIJOCEageZ2uZbwtFigvJsWltaum59RSknqtcLjEkt3bkLAEwarQqH2E
3/Sy/rTh+0PGnZzpWaAux5fmfsP5Hhf2VnX+1Si36n5xziDMxd9ZMG1vmQEKbfGP
3x7C0r1/4CLgc6gGeZ5n6yetVWz89VucVz/rNBxJO2NIJi0MFEmywM6qVBqBLBvu
Y2wgD6rP95qFD6FxL8cuYFjnECGoTfK/AFxe+wMtBglkJ1Q6ZKLaALukpNrmbzL+
qxYHn/xyHqEiba4eNCwSr/XxkdgD/xZCd37ucZ6pFjh2+3GYctDW4wFZR3d7RuQc
ZjoQ+f1F0Azp4JklNsi0pOITmHj4p/YyS15rmOHRt6e5ec4bUzOrZX4lDMSSS9FK
buSA71PK0ifkbGvusptUXzzsFaLMh7pfQHfL0NKR1VqLtXw3rNbZTt55xu2KEFCK
cqcKxOh7TxN2tqf9Mzf/+3mehv91PXI+AIFJEScpEPFnsnchxfIuKFCRA1tH0BXV
k8gGJtsmOmQ3FzG0g7iwrnpS63uWuerJVqh2LWc2Bmo8mNtdnT5gg0yji2b9IdGU
Kan5SHmNjfz/QU+f/M8gnN91Z9nDea2/Sw6cHyc1NWqSwiw3eiXQkvQeM3wLmEDH
Oh1R2IbbB6jP9kw2hheyV7uFQGt/5YtlXrAU+43kPTf6n9ddswkZlruCBCrB2xhx
aVIffviRhrGa7V6C6yBmQu+/eKmkGIoADUciJnxAy8IzZLyDowCK/d3/Q2RyW98+
uUEAGBZBn1MkeLkc6Y0sAAEYNqKH3eqsBAo9aWCyPP+gVhcWr+Lmp/i/BYtpzonR
SGL5RF1pHiCdifrI9sn6AhXy9zRbGbEYVip8DsOdBsk2Qsu87QEh/OIHMmWCf6HP
Ijh9oEViRKxrLOkEdeehBuH01ntlTGjVEzvzB3Mn6NkiIqx/rjB6xkmcYxarwVwK
ufIaVDNl2suW1YmCR/dZqLYI4w/3Wb5v3EqT5hPZlGxcTewGexs/Y70XjUIDvlXq
qFFqNG+hWwLYXNjtpp/n6DMx82PiPwz9q9YihUq8aJ6vYuUGCrzLgJARBwOQn/FI
r39u2yM1VoYZ2N/1chI7hZs0Us4peuvsew7LOs3+HqL6SoDSKmUMMJzxsCp4/WSH
rhfiN804Dh3TC8fMXU3gVrCuA28T2ETKAjAWDLo4abPETKlFsBC2UZ6c40n0hrVx
Qe2xZ/7bSO3rxuZohw30nnGx5kC3JmqH4cYipsOchzr+POGo4OlMuojvr/DuqrID
ELwoqT70kWBc6Gl7hFVNMku66UI7/ziJ7h9yu5hYexocRpxs9ScGg2XqZI+GaUjz
GZ0+nmf4jyiEBInAdrDd5rmPQ0k4RK8nb6v0/CRgRMwzsS1xReZOi2qeoFd82JCQ
z3cEnMJYMNRu9DQWefeybtK2xiO9wJbNI8Uuieaih5OwJD2qNd3PeW2rqxCGCh6a
79hzFVlMBWNRbH281Ks+le3GdrIp9l3YNxLRY5eAObXvJRH/BQ525JkmJTATI7Bd
76muTJ6bA7M9sM6OwNCUIQLF6cc+k/5ad8e84xqeC/kDcMOv25MXF7AFypTnIhIh
s0Ws4KKx6yVHPAxtlDzhbhvRfiImFRYU6wSZ7EbChU7Yx2g9k2kZtkDnIESLdiIG
vs73C5pIi+IH4SoETakvTrOtg0yktdIRFdaPuhfhpvzP0YpUea8TWzAsHix9qcDH
SknV3KDneqKM1WbkWx2+O349mNCQrPdgJCTLsndtNxy2yYrzRX5OC7OaZI/2lCal
ZwhzpRghcs5whMNsHYlemD1PTqnHZb1a3JmKE49SWbW3awNnltvqY8sNgNZ6V5gl
IgdEbOfz/H7R+F6hY9FJ/cBo9aFxgqiNXyAb84WJazZ+oOAzdAZ6c8J/OmnNSthh
xBZ2GUrCipCSp5E6/cLVRrI6r3ABUGsvqAv6TeMlSyYljnhRZ2nG4TNCbOHcxskg
2i2XuxfQH9YnC6J5HCbbSizrfpMwYu+9EF5oiu01EbfLfAOA79Jvi43zeDMn8oyp
eMCeRNqdY+CzWxeEv/BcEDDgBS4/tH6FFXswhibLNrEOwQvwq0iC3VNkYY0P41/w
e0/aQZBaTPnjMr23i1UglKBce2AVpf7Rkht+Y4uspmZRnXcE7CO7DBP1aRjROkf0
AHPdmratRQ13+3CS+rM5fUnGFUy2t3sjOOSHtw3Lhm3ZbYtx84NsxDgs7/NYllOV
08K+f7iVSeqvK03e9zcIGHQIwet9g8dnrSYakg3VYqjX9K6ammzKQw/u5zPsouVg
o9rbOFaQy4wBEAsv7FiqoGNBdlZXrb6HsG6nxipjNLga61K4ojPANkU3rQtVrqSn
dSiNvO9IJhYcyvknDo+zYx5ulvwjUB0hxq2WvUjtPyNPecrmfaRJIFFUx4hL3gbB
xC8hMnYrmtbwk4p2GrpC/t4GpwhhmnXgt4j9BqTspt4ejZCKiRDruEoCImHMmOg6
phLXoz4K/vjAEnSM0G10JC0MkXUPPqLsgsUG7eDympZgd6btWLm62cE0soniFo8P
7r1PGV78ZZ/+h7FoXYutaFYrjaV10P0zbrlFGa06JUrT0XVeJv19I4bOAVAUvVsl
1dQTKaJC9surLaffjo6sVOzuCSXtqSNEARAO8dU97xFnNjKYakavfTYp0Pvqog6c
qhtvNfbIvAa2gBclpiP+HtTpDdqUXaz9ZQZu4y+UTQEJ+zsJuuUqpR2ipe4yyWBI
mK5I8HXbHvPPo3fFLEaPOpLi3sB3m0aYQFEy0MS9akMuKnqWrJlROOZqXqJxumV1
XCVgcWGTa+AuO+VZF0WuuQ==
`pragma protect end_protected
