// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BEjA4zvX5KBOKZgi6K9jwbTIkOKamy+Rmlu4Z6fy+kyCjUiIAWSFIAcbQ72cVGpY
30VR02h9SDHsdEjAHjRahh8FDUplAc6JHzMVe0eLSQ50PSnKmWrUcAo/2T1XXkUI
zc7EraHJRaAtTY2FhlGJWrCEQCEmWHNO6cuwrQFwnTE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4208)
LxPihn3LY7oy6RgjmMnMR/H8COxUhNPRd6WholxYAIQVKjGY1c+3hcHRAP3wsGUG
LBs0rexQobAKPHlAEoOtR312++zA8oyWkDzw/0EFs+rFwo1qZBdmm3fVtzzG9ru3
rmnVsHlcDGXl/NjYZxhqaHsVw4bvzV+SbpIw31Ytmq2Y2SEHXS0Mxnsx029rd85h
y6i2Z6FhR+VvzOyQuES7/4P2p0QlbIFYx58CB3qhS7c7VWEwlRmryg0ufbwfapMg
xf1vaWvyaWHyUbATPzGybqvNLPBrRbXwnoFRhqpU6y1FrO0UFcwN4qA9+aTFuSf2
E+ccBfDt2a4F6/BmKVldlxHRiIsAmqePWDHXdbtPc90BDv7tbnva6/tS39C3DzZZ
bkqA+iSa/pPHhrErwUB/sSr9pccQOy404xeyMm2bIwGFFDYeMDvvGUQFDxpYgor7
SAPrIAbuKL/SKJlcoseJTdtaX56uuAKZW4c4q35/WUrYdBzs4RXLrXR/e0sOO8zj
xgh1d7KFeYEantwyKBKutyfkVKkSVB4w9wSsn97s8n5qeuSgF/zdcb9cG1AsVtjh
uQXUyIbg3iczIZSLuolLO+hDLSmLISGq7kpy32mK1nOZCqRtAcXZpYsFGBD0++js
N16Ud7qd05xjFCraEfVyfMcf838GNtOWfxsVjB3a7GgAnYOnjITj3VJl1LJ+1MD0
h1g6G6/4YvBGXjuQ8Z/cszqsKC2PuJD3sHEoGz16gY5gc6mzFghFLELQwEGS52dR
9ndxbotF/fWxiaVvaVk6byy1wR3WYTrQPiwpRhKpuYYChulubIu37hGDbTNo4ima
9PpUYoJrh7sq/SwvOlDg4uPZtO4fZnpGOyMg45f2zWYR3rYJV3Pb6ArUJjsqf0Nq
qaX2NqmlO8Qkx0ne+1MWleU1ObXvyXUzu8y6N6E0kfTpIPLn144NTaPsxRiD1OPO
Z0adpsO0WCbiLSfo5LrV9fOWB76mBC4V9H5DK5uRU9zYcXelAlMMdLhQzOIp6QY6
X/Blx8JspRjygY3o5P62aX01tPZohPSNW1zDzg4jrGvvOzFKO9YPDbkajh0wAIGw
AS3gpCLNfT57lFwwNcWx3JYeuEhlo0lj+NZF4S/DzFX79s0Juz7pDBAh2QSSLnO8
ljsdTuyDy5ywd96co9tvseTumaJ+QYwu00VxKqDDiJF7u2SAby8O4UR5sAaO+J2v
gTUngui3+RmdzkkHc0Od4H7h3+DDIsQDjdEJHetOwKMPALkh4xa+OD8RfDI+TxbS
uAUGGA2wsBFCyxYG2JsdQBsHpkggAiMmNo4CxesJWYtwBeX4UC0mn480EGdnBxKQ
We4cMkMJ09K+513+ads3ap6uOVvUrXyMoNm/YxRC0EJ4Sh7jBNpzrVXqshYssifb
Q4q6pfzyQCwMlPvwcdSEmkkwyzRC1rgTUViWRAZhb186CNhldBl7EPpyVhps6B/F
N6xJOoWVkYeJFsHrQASxPYmgJ667KuOPbYq2LyLNDw9g01a3J2zAHSFuyK4+T4fH
WxaauWtQuj3EkrI3npXWpuN98POEhM2iXWfL9/b4gkiLpQ3+Hw6f+l+PcrjA/k3N
uIArmbcB1mReVND6WsPtN1Yjmzd7xrA+EURFMWkpCOegm5ahk1cbV5M2xk1JpYET
Dj5LHp6i8btZBzDvKV2A18cb2v1ajndQWDki/+Cx/ZKO1xFfbwkRR2aAT3p7Tjz+
VAGqElcKmgKLr/MzBtSgwY5Q316iuVJ/kwl2O5jCm0XlnjSnzTZ0HhauT51BOuyx
uptzgvv6YVydwratkMUTfvVoXhqdpB8OT2NxWXcv46myJqV3iqQR9M5B1kp47/wY
GI5mopDdS1AiuFgpEeT3aHU5SYeFyQEaXnrmbndlH7QF88hIoXV/0l7rbATeZCjg
mIChOacXQXpQ3AedbX28BUxo8q+QspWxBw79ktfBoZAmw/ZkC1L2YW4A+d4AORat
HRWySsLGySOcRVOB4j3U5kj7aSS54KNyEZapSXjr4FzBF6iBGkqpfajjSRroYnMo
N/uGjx1GhSlBvhhc4/4KTr8dnZ7Gcg3u9dmrcdgHvUMtQD4XWud5peAzf0UMjyij
FZh+TLRXIA+kq36+BxgAP0+ZFb9zslaaDvqyYXuvVRibz+bjmlPKxt7+8Uwiy7kO
OaABQPbpVluHEIh/Sss4E8c/l96KeNmPr1JghJc0N+U+u3zpB9RWYUZM0Z8bGubT
SwtCcfHwqx/CWXcG/0/bv0ULNXLKqHozFwFJ/ZX9PNUO640Yro+KxGPrMMxHGUM9
d6LoC5UPUzrxpWsLnTiQQxWsAd6Cyozw7N7l+LCm2fA4d/EejCoO6Gdv30pte7Pf
WRfbxajBDGDocAKCejzYDGsCMkkBaNd9jtxiOg7Ji+7wgKZDb1Y+UMSBdtP8a8XU
HBz6CwgEEa6m2FS/9IWXoadq4qZGWa0rJ+6878yHUYm6JRoFBNcR6yqvISdKHMsb
WG7vBjpetFWtNShb4emK5PELjC+U/l6spsrGqQCNH/6ZHXPtqo6BeKpz3CloI5xk
qcPng+xuZ+JaIQxaKjVPfF9F2Od58cngE/AZidgSsFnIMAOkQZLqUgEmmfD/ni2G
2jUXeuqZRLuTIHrlfhsK/xcjxEWoNbnQXNRufo6UqvbA+9QcPTnm/Iyf+XZlBAV8
R2/9k/I5UlvUIFyv0YtpfqK+PthDx9jNch/mbIVegGoxy0KXBpfXov8375duq6ZR
nNb93is+VyxPryazeMfmwwUqh7dZtUKAvAPRcN9VOzIIJns7LKiCW7n+uetpYasd
XcruIcctY14vzWQzzP/MJRE09miDmRyvLAGZsZXzySm69FBWCucAEIeXHJ592Gl5
vhGKasrh/9GjO2CKQjG++kI3QhNIyp98k9YQqhQ6rAOK9aUwBUnuvCgEFwBa3Mvq
aqFmdl/TEgtDb08G5SyiJXGueH4ZZZieIb2AMJfALRatZ4AE8XIfTs3DwAsSGvt0
w760e4syHnza2iw2Ki1GDT5guSAqp7fRE1X7kBAuV9+qBzo2V4KK00HM/YRTFElv
P0hlBOhthcyp/OGe75mpF0uhCN2R1g7sA4PnatId4AOhxXPvIwl8dUTccfLcyHKp
7aB4+x5VWP4yPn5b3wxgTXLaFdnEgE82vUKdetcXMcfmjSYs7Oks8Tv6x8TtxlN+
s9Oe6eVpBpY0j8n58bD16kI0/JU/6V4fULhhNNyfFo1cCF7KzeUCKrMuVLXe+FxG
7vr8/JMTzD0tzab8ci+zoqQV7u0SAUbqFTRQwxOys5SD66oohUvGdRV3ALEW8THz
wuYYg0N/B30GP8t6M7njBZkHkPy2j9BL6Jmun0R5+qkg1P1pjVZ5BGm0wMdxgydv
PITCrj4RA73dOJ6tjRzryzR+ugAWtbAvjaQnQqFVTpR8EX5JSpGUD1i2SLB0GC97
UWD8XRJleYOLqCJK8BjbBhRWsqED0hhwcNSzJCCRB5xIuni7R0NkJuMJGn0WfmYS
sr4PIJ8fgVBApVJnqYrhw5ju4rxnE+XM3f0QNLQRpzDoooOJvld8ybgjOyzB1V3r
sCOH1AuKa6helxO6FXGcbUGkgpeE0sLJStQBEMPWrtlvpOhzP1TjxT2OIdJVzFyU
AuJpH66hO+CUjLZfCloIKicMd/cuILNg72rkSBnJIWPuzFdBd6OEQzM0YAFp/Jv6
oXdOGweChSC6bpff8rCaiRZ3WrDWocStDMV0vzpgju+sP3kvYoPxZ3Rdd8D4+69R
t9FXUgunBybA1KReOiii5ufqPhNWjQuEFsduLSLgwJ9bCKQNAEATw5EDO0N905bR
nZGmUJ00rxwPHbs2lJjQj0yQyc04N6cqjrXctlVgeo8KAvVJJlw6qwh+sTO96AZf
rhmGFhJZ1wcGkoN725QFAYCGWZmM9U9sVTQbMII8tQ904NVkPDPt3XkJusBsilSC
TGprxVNrF9HSjPdcE4nWTI2kgkAudq7cO9tN1C2KLTtPw/O+SIMhJ3HQQLyyD3o4
/idIv2iY0qmQFTSLDu65dxdlYoIajK2Lzxas0dPcM2gNkNxX163pbLpARu0gD+uT
1w1/M7oswkr+lC/wsi0cOhk/LUoh9yzDN8VdV7QRRx9DRKVm35MR4MRM3RCiGqvs
w8MNhicjsoOsFHxfzyL7xL1anKlJ18MWFc8SLVxENuKeLU/P+SQFaO9Sup/bR1ph
F5yeAcMjme0e52nzViuH+XkRd5xcbfxtnVWjtIF2KsbRtnVHiBf7iB48KHeCDbs3
ngIZDuny21QFDAusA/dl/bBdUhHDbJWnbT/vJUbg2sJV7k/r+viXvgClskiHblws
pSLn08KYz8U7Ao3hldqCFse1pGnUAJ7Rjq8uLXuXd3eg+3s40x6AWR1qFLN1Cvbv
qnDx5UCDGFu+3JxRsPI4UlpLiNcddPmfjARd7JEa6mXi6WKiRdPEVAkAqheOJi6u
m6a7+b9Y3mVW7ub9rmwVPVmfY6qK5O7r7Y9K02bLjveQXSPOWaoHycl5JgSwOuo6
VV0Xw/cYP40SwvqSS5gxRklLXl4SkFQEym5RQiakvFKRBrlm1CNJyrTyFfzoV4Cz
TsgE9+yU0JZjyT1D4lQgNIMyTTYzCBQpEu6cOfqPo/f0XDShnTSLTwVMdQikbZTk
a18wUxZFIXrBQYLAf1HjA06jimdJoA84AXqOGZvT0Dk9oBCnlxbV1/ePhoTM1VqB
kgGP27lvnEMRpJ8N0fQJJLtNAMvhbRyEhnzZh39jDHNhBb1/FbkPq/+GtSZ9WIc2
jA1fwXTYVLJps2N7x1e/pQ2vUSkCTPFwgOq9WbFktxX7f87VYhj+4ca906hkOWG6
grB0wE3wJXJAKMj8qIhPPAKwqre168E5XAepd6F6G6i35WMRJ/iY3q1cufEADNcx
dNzoGI85PN/uWdawDUDzwaAj2xAojAteJfhhqxHm6j6MNwNTU3dfo9l0tEkYW8tb
pCLzz6VlUpvTocYZHWrkl0XpYHbh2kvOazeGN/dWOSn9DosTbCF/fmFmlxjIdiEk
dkoCO5oVW1xLJKxhvwLdcIY/a24vLfboOgcHJXDG5AYhXlz53Cyl0/ip8a/tEys0
R/KAV7ij0sgyy/Oh4zYKoZPk9kGiUGufW79YQYIPM5k0V+VFBmiUGiYQ7/e1tDWh
6LPp0y7iDTHaRZVEF1k/zCjCNUl34bdjk4olXmqAmFEwBoaovZtS9/URTqw8c9mF
ZM+nMj8YRAczw7TsPUgzV3+b+XUwwvgR8ASH7q9FctvDinSa5/tasfEELSUdcH7l
2Lq3Zn0XhcN3C5BPOz9KIOQhkzVlZre+RCNJidq5auu3SfIvn/tLHYyDPdWOd68T
+SWxldF24Ty3uuKlxCbUaYnVbhPzWazFnfTPyzFhGb4HGPnNe3TJ6+/LhjgINIFS
v1kXXwAJpTQwvchjK0ZgcDgJPZVBTY7OQlgyTy4g2QxWQVpvFo6TyVdLmYI9P8TS
6XUqEQHoUUg53C7YfyVHEvCW+vGzO90x6PN3ZMMiR7m07dgvEguBE/h5GgTMAChz
BOVK1I03i9mFgVAE48QXoTOFjIu5o9aSNPbxQ1A7Kig=
`pragma protect end_protected
