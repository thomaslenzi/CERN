// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:07 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rkU2ynF2ckG6bs1SOSgh5h7ay8sbBbS7tH/gvcHhL9nKguw/dd3AdarNPCTQeOD8
iPOtqXkz9En3HAuwihJHGUvqQTI+3IpnxMgh5iIrDWYYfbGfYhpW1/FbXuQCBBgU
doSPvig4Ei+V2hDXQ7KogtPmJl66Dlf6QOy0GtyDVz0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 183712)
SChgPEhvKp4F9NJaoXv/2/kp4p8mt0opbMtdHvpmlIzUxubZ7HXwGFApfpUe+Njt
PbF2Y8kiDFFzTJOUvq4ETIFLL3jg6Us4FjN+3g6MMq3vkPh9WIq92r884d9HYoup
EODXl+zcQucs2otsYofHqpEuePU6moP55UVqR9IMYw++10btulfXZDDPpNEEvRrE
0oCgUZ2gtxDA1jIMfvBM/s2odxqshksGoxYhSgkgmdELhyHXOOpVnbMvZzjntU24
whzRPM+K0XsbagLMHIzFB21f9bR37PPNgSDUqogjR0cPheRzHO1Nf2360CpVB2hk
svBbUoDfEd4xVV5BbPeXJ3T1MPFp84fyhrdG4HYq9XPXN7xup1ODq5fYjdNZ1ta1
mgxsDxY1ZjWi0N3m+ZxrdxAgdmG/peGrGFgXa6Yh3MaE6wOKZ0NiStSLlTgDT9QR
NbN86705A3OuQA97wImqM3YDDR/XMdgsNjLcfIXi7cxqTQ+n9hMgdUy44hDGqG20
AZZf5EmX0OkTgPYsJzwVMpL+Z2+rqMpGD2J2XXHcunxEsEivOSGq4dm/s8BrUpPy
unH4A0lL0BZqKsEhpyd23YPrinni6veBaLfazg2Sojzbnt2Dw/CMNZrsoZ58kdnk
eVpRNODpfJ6HNVSsgqxfUvKjdjbZ2lC3BYQ6ftJ8psMXooStbrsz96D+eBvWStWZ
ECfRxVJLyPB6R9qFq5Amysm88mc8dW8xb09Rr+fFAOPDMgZ6W3+cd0w2UQ8pdIcV
5AO3Z0Z3zwZ2FynUlKe6BYhn/0EbAbNvh9rtNGh2ThQYHkvZ8/Ssq/AjaQQIm+9B
dae99WuRFOquA4dxRjnpz4Y3+qgPW/Ie7UOBv1IWfYgMc/CFFgUdMvS/paNHGZZe
kugIqLwVkp2AVbE+jOSoeg2Q1ImNBjbigF/5otwzi62zhPsPKxhMHaLUuxHccwB1
TKhYhPOtnNl/cz8f9c2AzxzuGtOKfBinxVitACHvHaN3AGefHveJKbXwsK1qTVfC
DwINz5/xxj7VKcyHEvlj95lRYEfiQZZt0ObZeUQhLjbKuMR+wlvyRd6FQON+U5DI
sVW+mXm0YnJczbqTOHBpfecO1lbQe5oe9dtI1JbpMupYO9q+rytBC/qzDOFLfaBH
iJitZN3BWNRPyqG9s5JXRwIoBjDw6FC4e2CtjTJE8OLpCSx5ckxHWmjEl4JwmkqM
GtK75NF6d384IZT10aYaw1UjlNmMNWQuO9UcH3rJBg24gKJMztQHQV8OtN6Grc3G
+1HY0E8Gkveqr4Gvxp1hXYZaJihybz3IDCFp+a1hRdvhA1fapIyL+mXykTjfDOV0
Tp4j8FwVTFe4U5zl14a9VoCuEbU/s5aw64xjSRZbTTtZVVunMpTG5cimdY1AgjZL
v2Vz7EPnRYCOhK8eCdRknEcsDQrQuoe+wi+2uAcPHkE4NXUrL9VKfQJH5nNvzwqK
oXA37qaCLnNlEl1+jC/DFeO2+8/LvV4brNxUurZLDy80MVqAnKNHrzmdPCRmhcMo
DCaIQV5RMoTkgUIB5SHv6l6xUQtQW1ZIpa2UYbr+S/RB1hMg1Qp6oipTZorqpqo5
0+bRcJrq03anoraZhYMffteeUuZZ2u5AGyOQirtgzlVtOl8z7YIuLg/h7biicfsL
ZbvbnLPlxLQD5pzgJVBJ4Ks/Frz0mqhUbb+VJZYHIe4GeKLGjcCQvvcx0qhndlkd
1GSdEiwcC3lMSeXCbiFamYIkaDABI9diLdIkRWC/W/x0McBP7VqXADo4wGEmVUEY
eeTT+KBxtbTASsoQTZIoTbYi15CnXfT2WH5Qgrl11Rux/WFpbUUxvjRYxUQ1gJwe
++naB1gxUZVMazg+DlqhjB10k8DY2dNN+3L5/5waTD8q7Hu854vCB6HJZUpj+D7o
jbRumWyAbUErS4dsx5zZWRsTHD91900hd31KPIbRN3q6lV0iEiMx7W43nnml0kNV
FA/gKhPCAiRQPvEdtOi7YNGAls5Ppg3zclVVzpoFxjstrdqc2Alsg2riY2qD056q
8p0/oiKRw1/KA+HQQU1Z82xNslqatLUfRG5KfIi1oMKo3RrhhhIAanvxj+p9aVyp
LV/lrNUomykUNxc2Iextw9MZG2gnis714c/A7P1o6dGM8HI0+T/rTnW5XwGb74Xc
GfRVAvbp7Mja4ubKlCMqaRg1v+EIwnH0ZO2RETlklCeFFBZBiBQqVKoMhN77+1VV
PT94eH1EB6qgPJeNjI3jDBMlIDmbTz2LHiWUmYZPNI81P+3gbqrGa9r1carVl12L
KpITiD2r79E3pdB8w9Qhx8oGnRc8Yk3N2g37mYRBhIH6AGKZmhILWNRei9cVsOgI
/H9Kxefm0G+Iz0cKyMsQJfP7jiKCoS1hmjk8mq0T2rVKpSmyZS6X8EmFaCHrHfVc
NnVYZlEeMwl9k5SDDQg7P7sMHFtWvCNe7H3kyLwIFrsiLMRnFA1F58NFgsADQ9HG
gs+jyE3catmJuDywfUvQxX6nHvmKl7TQK22KtW0aUV8pTEcS0bhYAcY73xdyc6R2
zU7l5qV2UtcPB4SWGAdTCEg39tsUrRl4KZmMybhSruQxXLktwlXkxny2QRmM4kKX
y58P5Ut6GLPwoh2KcI3djhjnZ8k+iXuugEkhAgY63zUnCEAjPlHUGJjJjZSsxtMS
oo4QHw0af+6kBdexeOMl5AoCKLkDvwGRpNMpnzLEKh5yvwJS/C9hiBGlkIrDr5Cd
bx1ZDhlv1laNCXokFDaeo1vPLiQOTqm8T54dSrnaY347xmdhOAJ62JbjdJJJrt05
b6G6GvEHVelL/jfLaRd+OeO3skGrcQZgGmyjpg/fp61IT9cz67NE8XakO57rsa9S
5TFTZDf/9hASgAHVe0JyRPvM1SXd8K4cSDH9Y6hBrbb5jRPBMIqj7gVrodhsMgUP
XMhdNYAaWKhZS0rxbEqCO24BgDmvSm8gFzTCtvmPD72q7U5TLvXNe/wQsqdARlbn
bK+GU/AfduztxIqUl9Kb6SHwKRHjyihhvFrCSdIPXJj3a3JNe7OT9ito112l548z
Z7wWe37IdeeUmRjlvUKfoOVPDGfv/3CFOHnY1zRlZZejpa3DmF2e+kmp/Gp+TwfV
De74CraCxLVAzGQ+jjQhj9SDd+O6PQz4wzWJ1aXa9GDNgiTeInw5XQa5mblMTDhi
/ZYZSiPOIciYksRvyjHDNbsem5HTD1fdT2teBA03gUSJwsr8441Xh1rvL6wHKBTS
4JQLUBpRFdIGVxGcil28bX+w+a65elxs4mcnvrpM56ry5V9FjRWQjwuWddmDCPuN
KdrKquyACrsz7khE5BL8Uppm6YVbI5E0XAFNB9VZn5YBv/nR8GFBZPXEkOAPL4dL
c+r8UaPr5iViImiNC9TiuN/5oAbopMzV/hQYQxPXx8aLjzecLvpiKjyttdRrJ9EN
4nN2Xd201QnhF1qqQHHxb1AL/Ppf1J38/71sc85qBeYuXwOm4D1IqWfwV9+RZF9l
tceKocmYQBPn+sU6rAf4wO7OnPwQvacOqKrti1Gh1+XNbxO9CS6sDtHgGFx5mt+m
AumbPP53NJqfJcDFitpn2oJSt/4rawCckuMewG0C8aF3gKL9YY08hHKGCJvN+tiS
ls7fjJ9/4fxyIn2WY1Lxv0Jqg4+tBVCqgsohw0DIDLq43nLn707cdNWZNF1zUgl6
AgDVbFmYQhtMejQOXeQnPTn00u2iuwe7w5ypwtIc2+wA/U6BGaIbhAGFxKocjLVq
PsmRmX+L1unQrdMuQXPhWUB1HGEHiHqUvGySj9qrMZi/JAIsQ22Mr/HwSRLq2JEr
vv9bfbaqz+9nIBTYpco4yT31YCivdehFBql7aN539IK/Ek8X3Fk+fzsFDPhcfsZb
EGv/VhqEbwgxlmwb6HlOmEFhIeaSKGj6QgoHKRsp13gjgzfesDC1ReaqeDcBLjVM
zSs6HGOYu3/4kwC82w7wbXqkZBNpSJa8nQk6KZVOaj4sQM1w/RwnJNUvjRSwjebf
lqzLYBOvVATQqbLoXDxmawYBZgiiqDKCBLJfotoJwbdvjKb7jKQ2KloW3xlfYwE2
7lvqSQnFCd/WTuI7kDis9hezfNy9vxlkH/IKvnP99fQBJFYdYeSAgBMDoiqNT/oJ
Xyy+7gnYH3OstDIYhvagQfgKIiCpBWD6owxDuDkEyHUUc0cgmTpK0LhM9Ls7MJ4u
PzbQwFYJK5Z20Ik2mxlxlHpnlEi7Xpd2Qkibm0tf5Z+xemM5aUJytN6LTcSthhuV
TkPB5jSi9eible2ljCtUEVnJAQw/JETpLEVk4CGUHHFUJnGa76j2bx5YOt5dIYfo
SD8HxNDuUdTEECrJKygqEMF751vSWfUF5vpfSPW6RFq/mmzssIrJYbAvyulPLehO
9U9YJTKPPatlhgkpxiP0gpmWzHlAhucE+nEQX9o09kDIu0fnoA3Y1euDdr0h+34J
jFoED0He/geu9xfdZVAR5CAC3NNXcR4pb+R3a5hIhb+qWvm+NtodBwUceLQSl4DT
2ampLaeHMkQV7N7eXrfSaJ4/jqJoEdexmTJhiaF52/6V99N49grSBO/jTfNKCOVZ
vDSs1mXqAExLTL0Fmer/bi5ggcqyvqpB/weX2uygSR+RzuJWTGr7ATa0c3wc1VOj
jVTjQ6IIxxUZVO9UUS2rQQmIFV9sfd4K4rc9amIyx0KHxOB+sxiDVKZV9RTnZsPH
Vp2LgKaHKXONSlNl1zZZp4IwuQUuLcCGesVE4d9DmMFZjsWQ6zkzRVBTfymmTGhA
PUoEzvgNHEHoHcUF7OPzLLmLbMmfdx/C6ShdVihQwcxXIsBjGmMquLlujAonWQJX
6J0IoXxffXCI0ryIsntlGV5Ts9ZA5PJSJR21PU4cdsut6Z27rJL4vH5rdov7CkNQ
D3aLKo/jI4qMfmOeETLk8eRXWOe+Zfigd2ja0p639P4o1k1Htf+Nq91Q69ljKnkV
FJS6hqV7ZkPS6UXqoO4PUNNZRKcTySDn5tCK2fOhcT4P0dnJLv3nDmV0pAxqXwOB
a0L9SkFZ2J8GsYDmBEca71nyuYGhyns7Vf6wIPkABfN4Rzpx69AJhVh1jpds09yS
suPYHeTAVeX03MBmIttpXJqgeNygDYGnJcns43apKLPyaQ06YEykkHip44Rkvkvu
pV9/qWUR8YCSt7OcZSOmJCaU/sT6wrR/5K02yQxAHJklS7qrqicfZaAUE7otugTW
FI6kwsO5yO9+VL+Uc7UXpNoQEDHh+b0xyb3egun2hoe4MtRUlSTyvc6zorD9MZFF
DwCWHEiqOlmHpOnmUF8N6adt97jC0q2X6aq8jjSg6DoEVAEKs51Quk6FoyWaGS+j
jgAjo9fNKLrbqgsvaQ/c2fBQE+987k21A9HMHunl5UKTDrvrwh05ZsOiY56rnAZP
jgNNpan7PGwHUZZWn4IZXm4Nz2LySfdsT9p0RhWrNSe1b/cNs8rQ32BKLmDPgSfm
YtH2VMr9u/Uc07ZCo7s87Z9mxw5hHes7hLNlAkcVUErOSQPgLem7VMxcGqUAeRbB
WuZ6fX+vNG/RtnWuhQf0gB28nm2wuus9THEXOagmIxRqtvtTYx5Ph4AMVHGRZ0b1
5YRmmEGcwFmxcH4lOJomZstiriHqqPn2NhuYzMKJATA1QHkQ4iRZ/7cxNiAjj4PH
AALDmXiIKX2phe3L21azkcoQXgaMXFtpQCJSJE7QhbpCfAhZAdHZDd04Qcs/yJXC
ATYV9meIxOFL5b4Enhc7nViwKvdnD0ru3CG/kn5pJHH1/eo4cH1o9JewYnhBbfnH
1W+7bU9cx47KZV+IoXa0xJBvfSzm7luy5eaa97uvhNh6RBuQ81C/mTlo2mQxt4Uj
4FkZFkesaiZMUJ4WFd6nRzSL6hHb/k/TOhtU5GXD4UpRO2rRCD6GJMbOQi4DuEPn
QLvHt+kBGya0yRy35hJNWuDHQRvfzNJ69UVksWNl1J2Egi4/cMmTAGbcRCBKtN0Y
EWL5Zd08UyXuacGeP/HMw++HK8BCOnPTFQVHy8toFjVx+6D+2/f7uVA51tUHe/uE
3N1kXGBvUnoLNdqKd9LBRkRa+Bel9EFDXgwlUJ8OJL65pmPhMFspmeKtS//LRgfZ
38+FdTaPl0xMMAe/h9oyHgKVUUebAt1TrCAww4JPrTL31RIxDNuvAeloS9m75iHE
ZM91i7PjhYwV8iLDeJ75t+R+LgGbbtZbacLgcKOAcKuRm1njCcmY1XIBbnOLwYHH
FWvmLTZJ5nXL0ZxYkEnVJuxSDXEsE0wX8RQDOCjTDVJTtlPCRGK4Gh0mai1PNhEA
OUy36N2wCT60HyaWW9BWTxEwSbtwiDgowwa18AN1ChbNlzSLVSNCuVHxMcJIgyZZ
jkIzO9XyiCjpJoVeOmbbqoh5qM9u2kcI9H5JU7ih1Bv1m1C1EXPUvMD8ZpA4oR7T
6GEXnAQmyob2XoOw0kX3fV6C85dGEI3ZvQe5/OkeHIHfA+TST21neUdY63JRNyJ1
k3ZmzDrMArEt5cFtDIYkfmgprfSRdfCNh+EkAUO+Du1HsSSLcWd3q2X21ynyHhT1
Uc0+3FTY0bQBGZ1YHfj618OqZPX1rPbTEoAnvt5aXeDSJt03Y2pwTuNjHF+SSN8y
hcApnHsooodXCFimK0sxr66FP6czqsO2gTf8ArqEmfJEgzZlDFLHrljrmr9sMjS3
LTZbe94Izym84EFZBvCNQD7DcMuDvNFhfHGrqOGZj1rSKf5r+PUmGLiAhV6+72Zu
8U/B7SOjr9LHx2i2FROUva7qnOLv6u/Irj5g+0267Z4UQzrJpCvMj2SLoYnNuEcg
SNluhyqpAVF9V80iIQU/+PS9LLl1AlE4g+R9GcEpG1Jk4Q7uBq89bKfggGPtyfmW
tNgeWnI3Fu4Wz0SO/TS4ii5rFzvWoboga7WxJ37hsEOtJ3naNDzb8Unw/NAgeIfa
18bsfBjpkU0kOZq+f3QDO5Eq01woDAMMATgpfEWRjzK+t5eri4kmhrmJ49yRIS9c
uebecV4USZb27osryoOC/urWGEvrppcu1t6qFqbZhY6LCGR5GbHgI5ctp2m96Gi2
wWVKvs6ma7YCJmGUzL5tbIuTgo7QmtjtckcQ5731LnhWtO8p//WbBLapv4j53i6R
krMhYaDneniqHLHRLIXqaPM0s7aSQEiSZfwWMdthS7rW2wzKzLQbr6aitS9JE/eu
UHKE6u7fvnlt/VkBCWAqXwFXam34WdelV7LqRNhJR5s/J5Zw1doEV5xQx2OUw5YV
351m9twBtHeAa7IXvceJzNW5AOkU54O11WCRL3dlnHVPwtmYrnDoDK1jo1vOxz+c
o5hif2IJoSTQhjKuDmqzcTAjylvOs14qFQT/YWDam2oEzBI6PiH7HJuuzQxPZHUp
HS9iXlxVxX1Zy8exClUm9Q7pVwgGV4PT8HXNlYEQt01CX+jmbdeA/pd265QZabzn
dY3wXXmzbFB3o/BXsK79ciV64iXWRPFMKjNE5/xl3C6guJTvrwjrKMETjySnj3Ss
8Ma8OTSRm1oAw1Umx4zPXBTfbrMq+boiEl+gkbKGzHJVYr1ijv4Jb5OTr4yQStiF
p265sGEH5A8jQeC4Uw4VlQrT2C94G/nvVLn1eMwFbR7rqf/XNnPE6YtLD4Q6E+xz
ByfUA+ESBTEdvvMu/3XvSLe2RZjGoHQpx7UyGyQqrYsU+V8TYT9JPOimyxMsueId
zhFvE/DZ9N5QAtAWjOrzIf0rQi8cKrqMxcRED7GK+BXcvJPPbzwv2YF/zu5sN/UM
dBHoPNwAwc0Uerm5wpScRJxzGuNPrypf1CuUfEWtYUsc5dv+/v4lx/i1/P/pc1oQ
ZWdULgrLcFlu017vRcsLxJNKOYhmeYtrwN0hhsAxIJRyE1fVPBS0LFCjRXQV6IiK
t9bI0ahwJ7NObqYK+mIG8RhEXkDEQuwYKl0ny8dCveMleFOilDp7+N7w3l3OYZMl
1WVc4hFKlXVtQJeq7XgJ+gZYEeJ41DUCIQS2S1KNV7oPH8/TIO/mLxl9kprm8EUZ
0u07emS3mm7pvN0x43iu5wKhi+hcY0Hzq7MZxAUTsKhHLQwq623EBLtrtZlQqAAc
YWE68P46jn3IXn2JHQqCfCTFsyJ9G1UumZ57jp+QxMYmvWrbEBOU/izQXc6XyRWH
54bhZUFqM0OHxcYkuhgIdE1etCQeV/ePy89KhCPSchHdd3rN7YiOqWSZ868QMbji
g1Pyk704RGrxMKy2iMRS9ZUB5jKxpW+RKxDXLK0MV84qr4AYV7zlDZtE/nNIR1Sb
/HKtom0dW9jhaXjHwKnGLt77zRJlzCVpucWoHMtVLulLadUKhWHwa3jRA7CjqIPi
WiZaNYLl7R2PtUEpu7atwEEsiuxKoek4n/lEP3qEyXCt4Xjm4RKYCC61dtZ1cRMJ
rQvUGNjgfigHejWfegnU+e1DXeypLWY1srN8gmFUBF0kzbTf1ng9sGfxhDDML2Sj
OZ/QWfXHQ/mrTqGiV+9HtGGaKK/JZbRFEAb34itSJ0686yUEZCdE5YgXKbp+R9L0
5ttdWGaFrio7ZriHbLp1c74wHuZcBwpmfYGw0CoJfNnvypbi7iPnxivM63QbC7RN
UvV9DfhSvEkxwbDW3Xxqs9x75Eo1Bxg7djLMra95IJdOBwoDvYoFODOIomErZJEY
oVI47nNeMgxM2A05B2zApXcSuOIxDr+2/MF3ykO95rZJ2/jbaB2o3TkjldupXSnW
sG06hkSkyjdk0A67MXQiIBZrjbsYbH2VNzW0phmHON4iXUH9BYMEYD4k5U1Bizhz
EaxTywDebsCmdlKAtDyFv5F4qgwgNDkZJtRQx0KSy2oMdLBwdToof0f1HYlL9Dab
yn6FcMh1rySmNBh3K+ZDuFrcHDf4T68Jt7YXne9kTqvjKZTT0fzd+qavSEeheCOK
yCCczLTF8bsi0pqxCu5E/12+NyFEWFU0ft26BohsYbNMirXy1GjDzJ6dWZPFgVDI
JTKDLO5ZxAk974k1WKcWfHpkRmkewIPgUGyR7BgdiKOwSyYj+Ik7rpFUMlkXthGt
XVDhL73/gB92tug2v0NVpIY/WZXgb8/wnaMcF3yMF89D6u96SazkmEfLyI3c06sm
5peJtDUW8fhrtl2F+R8QP8kzY+tFAMf1vG5j0bu/YdCpvTQyGw3fw27/hvqtZMVe
7uzvSioYtnNsmesfPlaZWY650J97GtLES4A4Fl0oYtyyC/yWYTgnayNCp5rPHyvr
dtWy0l6zwDV9oqh0ESnsRqpWMcKk1AN3RHQksmCpgwL357/+x2yoY6ukbHkzTUX8
UxtM94ExVOJVYIiuuyr+W94WkWImSuEq3ctyl6CCkekWm0AHq/HVRi5K7mHXcEX7
idyE5RAbUzzZmnoit1YcZT8B0EHUxQeNd3wvAI4UVy6DeDT77RxedARP6KXMazHV
5yDzyHN/rbHo+BIrVr3chIO6RwTyGna95I3y98RQZwmTg9eAiQKB0ftGtSAisZDp
+IyWgWp5WC8rh8kPN3s/W/hExPGsbLQJweM1meMuvekt5EK7rHpa9R0RZhjYn+Aq
qKMAfoCviQ8DJneDRtrr35DXkyw7gvNehgqWmXac6bPBeSz4duFn4l3yrwbHl6x2
rF6HCJzjGQ/ndjmHCj5l0dTWVYzIWbZ4WrEzBpXP+CkmzTVLYKQezJPA6lKT5+fb
Z5NXUwsTw8sPZ2Z02WprVghoGeb+HSygY1vGCGEk9zoGm47829rFKVj5fnLv2RNH
Q+GkqSqSqfq6hDL1X13sxgYVzHetsKqzEgVnxDGOp/6J0nGeL2se4M7eaoMTXgEH
GPo4WunuQVaTTKXOlOGoyPrl8BbjUDJAOFw9wjjLdnUD7HhDVc+zSWsM40VfOEKL
jG7K8hb33GtxF7bo+VaUtBIFjb+/PgQiyE662sRQW9wlHrfuP/CyHQZ5E7WPwCjg
w5Z8H02zgW39xD11QAee4pdTuhbDzUWB+pAm5L5+AYLqhAMSfOEIKDItl3giX8sw
OEWb7wFRW6eJO61PeBYJO/DJU32JoR9F8puTVI4/uwOb9TgOjxVMyVYyFwCk/hdi
5Z7GfvBtFM9NZql50NkXM87RG9y4vcHbniVWgbpI8IcgDXauczeuvLb2z//l8vZe
y1eN+U+IV9wraT5zLA0apm9lsdHkJXwmT8sS+HSba+AyQ3orwZ6ntZ6iPZ/Gy0IR
HWdUUoqgxeuC0+Z9NtvA88egGJlChLLs/Esw9IgkwgyYmlzXStZ0JWeTC1ke5Y1H
2nR9W7bObgpFHP20bcMZ1QsIfmwoowzNHifq01mzavpf+BAbwR5xoG6knarTHCq5
HGSlQ9ujhpllFCrY1ynlRuKnfoLacCfawQxm8LFYjM1X+pPW4nqPRVDOI3y3JdfK
RihkPrK45uKsNyQWYX0JBdz7mzbxFCMjCV2WQ0vC4NZgQqeZ5WDCZPOcYVo3clVP
83eveETG97us7n0i69TTDNEVZkMta5mNIK9guGfZoIMkoXRnJ7jtyYvXf0moFhSe
42rvE1DDDSDI9UWzKWZtigZoEdZcV5cR9B57IF+afr9J3GINBlWr2/AuEwEHBIKQ
GHZl2Hg5LlykS0P0sQVq5LbK6GUqlj21bqw1onEdL8vaTXj3ENUPOPghHvPFcZyJ
T1DSz+Q8BFDCYrLVR6Zmy0f6EE6cJC8xccfTvx16of59dWypLYgYv9WfsV0YOERW
V5tVgST3xmA5KaF0XSCcUsn51uVuRbQDSO2qH/IAH+GVZF4hdCYACgVNMvO03xIZ
OycjohSCVUuRACIgh9/b7MvyVO4D9I5RjbFHmGzuc92w218ScYMVN1WdbRLWSHFy
V6e8XMDtvSQuPbKfeYp4lIFtD20RSS+szwtQIu/59IjOqbdFor1bQ2hi2S2mCLPo
9nbVNr1h3ov7Lu0hnYRua3EqkCN6QLoC/ptJTJq4kWrZoEU/1cbhTlyvOEMGbdmA
bK9SbFhR2nqmwW70XYeXPMEDnVyuxlSYeMUZiluZY/cCxLHd50GR/D1dKRwPJMfK
vV2PdQAxSvb4UtASC8zatf+FKAC5zEaFinAIDldxNyaO9TxGSQSpnSelE7K/3g1v
ukeqmbFxVHg6adCcTd+R19DvgJnb98nAOGba6fc9z853RGKj5Un//+EnQKE64mbu
6XKEtKHdXm7qgCWXjMl8NZdDU9/rz5pIqlYc9NonDxgQRMJEg0apIlU0LZmhcXrg
eNTg+kCa8wEvwbAJcyGUZNps+oUA4DoVR38GEIaoDQsGXfKibF2yWQctqF7WSmms
/ryO2ztudAExTg4OdEbZ924BhtaCZ7TWfS8YnrhcTHNvkgwsRQWXn2YXOZsNrl7b
1TmVCBOl2lBZEzSbLJhwp6Kln9FzF7cT0TLKqS2JJO4DeXy5L5acv6ddPOyrR23Y
d0gk2D9ikqDSaQCUwooW76H+8pYlftjK9oo6N0UZZpetDTNcIWiBUM4ue8DeN6IX
bbCl3iwJYFgvOCCya4ZAsBfxAlfhvLKc07vWZLciYSVwZHIwYlG6sKbEJuU/wFPU
VFgsa2du8WRpoVnRTzLcmHKlcWRf91wMrUW1gDeEKpIR9+EOehfRY/3/2VTAOEYL
wuhm5jj27EfsobJta5V1znpF1n0+uyW+mimUShD7rQzKYr+EldT2R8ABBA4BX6Vn
QrPNrgKsld9bcarYso505Xrt/OUqZRir8/VhP5x8JkB7g1rqm/4aKsccbLocr2FW
dT9LZHALQippUL+V/KgihZXRKaocE8D/91oLT/77gkikVifER8jj8Si6Xn5b89UU
Y8j7tsqXGKDXX0vWktrYe1Dkq2K6dKx51Zi12HakcDUTTbkZK4kBwy/9jA8LHS6j
7J5fVYwlBv3rFBkDdQ7MxNjh9NttfG/Z3CvTGKcA+CFhKko3DM+Fy7vbhb7PGwg3
utN8QxosZR50Q2iSx+RfyI2wqsj6PwkjvqJt8fufY1BBGMPbzuFKfkN3tjoCag3Y
OVE3ZSOxHz1B75m4jcK99zw1OmK3pD82Xb4wEydcqYIahl4SraWGsATUfBwMPF5B
UdspSeBaITftr9CmTmYHAVZgvWiho7iioRKLF4PVn4/quWr/iUSFNgsb6lYVryCQ
FZCkedKu4sitmtW13Euv/HY+zaMSSurfdbNYXS6NvzrmLsZTssfTfySKZ8bVzqs2
l6WaRL0gTPryf8PqgED2VKquESIUNlLCTCTRj49Gt+JWEvF+pNrGcMkOy1PwCEI/
+niVnnuLxxIVrVorgZAkjQyuoFyCpEs2aAfUbQgjiLu4Sw6XUQM7nW7SS1IroBaD
R4yLTX3aZD4RkFsmr98M27vjJWTTveOo6MO9/vB85004iHjpP/bvCp1no1ez37B6
ULNks87LUObUVK4tXKoFIsC/lClws+a1sSIsd34XYu3HYuOCvwHitHsX0wDCCqxV
4y3RSk9Mw+CkohC+jQJEwV1NbWBfxsAuVFQtnI3pqEu7HyTQOQCqhUzntbRVW3k7
7xffJQTpHp/5pCG6NirpQDDULBdeVu+3U0uOaot9dvniv09cVN3eGbiSAMGlgFFi
Uty2owdh84HkRUWZrYE1Gw/uFsccGcLjf5OBdSZzKYlIg7uFJrYYDaml1tkEbrHq
tlW4dG1aMkM/auahC4UO7Q//LPismFjtxGuMPyT9frLyktThdUAiW0QhED51Ob3Q
HAcMc1Dg+D9eJNp9+SFJOa5/bWx9aNNDDX9pNVgYW0flmmKOlHCtuZvLspUoAUf4
jm1QBmBFXDjOFZEpcE1CSFggv8KB46C8lPEJCmPNd2JYwRzl6ml0IdrksTjjwZUz
p6V/vMdagu1MN9RAFssT8KFedEKpWAfnNOchMksUrrawTiVfi3lTDmiscAMivQIw
eBAyUO0inYuMjOUDkA0jtQaPXCAUwpxuzKAQ1AQtlz5hHWnTXAGPwh7wNI4aIA4r
axfbXEDZejAfzZqPwVziQOyXSdCSZsEWsqx0JvqrBZ4L//otBfczL6wLRisVhrwj
TdpBMP4zmfVJ0LbuxFYGWnaJoRqKw3slKz21qA5JbF+XrEmboDsSeO6NRYbp7wFm
3od9/etq5epn6l9s9VTOSL+jqcHkJAGAAvMmIHyCUwR/F8GOfJZiGXn5j7B4u2bX
YRd23Zpv02LOVwJL122b0QDkzHt3ENWI1yVrLCB9NfJ2cFa8g2/HM7QFZbBxnu3n
gJWO9si2459uC5YTr0/xp4IPvnv9DqDO1nfbZ33J913w7ECpsjQQFpuBeNQ76VYm
+fMGETgfrDU7sBSJrhxXVwHTOC9RFUlXlA5GZpcv+DM/MrwaWvhRIXUV6+Gb0wQb
Pw5I084MCnZTgYLehoOCk0CJWdjXeUAZPaua76CZabgBwV0CLIwWADhWJzCjDQBC
kCOnFHRoNHTh6vXOgcwl/3opbbnXokmTHT138ijWqqD7PmaZMMmMkTUZZY4nM+We
kmRccIzX/zotQTBYGXViXJRHXkASIPj1VG2o2sXQSL9ezWQ8REUvAaPU7+Carb8v
J6f2ckQy4DVnqrowTt0v38tFKU/RiKwCTPhbgOYrQIhn1grgVzv8LlI0Zh2oLwY6
bjIvIuizgRIVVNg9cqMJ2Mifc2HxHxeqdX1O3ZcjBt7t8cm52Iiz6f5vgSkTS4ZJ
C21vnva9Kx1gwyWq+7jiJYVQ0zVNUlmDtngQngEuUmUDv2YRR5oggsMCpOOk3jqj
Y7ThecM+QXZQX8SyMm066OgZpAffi+0Gt436MnveTb/a7+TeZ7ckKECUagCrIFyi
mxWYKZ7uud+uJIm0542tffOjRdm60zvVxyIZRQjZc0Vlj/ni+VPOZjtipF88Cfr2
hOne2qnW4/nHFIsbyahmcScAjg/+W3HSYOzl8B9UuoM5xCwmLCU++XEp/khJ1Sz5
0G7LRJJoX6pbDOO1I3u9hewCCihfdIWpo4KcUJWcEaoEtfkV7bnHqN39Kpdjc/mV
ZDhkySDaXlzH3GOK1ZzZOAhjlRGJj/ZJppGHN/py6JMcch2/mcCac/pNcelp8sGB
Bt61hUawTeEamJqBnfkrv/TWANBAYzhKvMNfSZtuQPHkZYImTSRWYe8pGeQcF3rA
1DtJOWm1jU+d7yQHKMZAd77UoP3zi+H8jXXhmRSDuDFCC4OVpKr0SDRVuJroMLwV
7Ql/oYhtBbRwg4Q/QO9o7wYGP9RTqZWpkkYy/aihvdJLv9iwV1QWZ6ZifIwm2w4z
melrKDo4935Ff7FWvKw/OMUXYZPKqdatDFMb02sj5OT/yGCHHdOCZOSgj297ck/l
+LVPbJc9rfMWzyg2/EILVNHYvgR9UAzzoqBrXyuxC8ki4oPCtuTmYhbpRl0Tlw91
NdjttrL0IWZsvJJJtQYQu940z2jc6HO6W9dW03jN+ZEeRq8ZYjvTjxYsc/Ab8EMP
9My9Ot50ua5DjiQyH4koKh+M5VBfPO76d66jnmJhbfO6k7oaDtHe9bh1qfYm7Ekc
KHCIMaF0AenwAg8QZXUMoxnkCazMrXs7BYYvilWml0x3yWCeDBHprFZVwDeAuqZ/
W+eTdfncTtvA6IIo89GAlAWT3Pkk3ydLlOg5kC0+0UTOe/oY9lrVaSVoidySrbqV
tzNN+jDS0DNO9lrB5JvBrjHlb3WaA/5gghleAHF5cIf+/2nw/ROTNUi7QUjq4g+U
MczEQzJGKxamFKseVQj4pmsxNbyBqVBAjywbLGKYExSXja9bkdelipCHKFyBoD3C
+8t46mvNxcuWVDArQjUM+4gFqZWxbfjEIS1w0pAdLW7lQv+1CkgXsfMGdtbZ7LHu
yXY4t6X/WXcRPLkJBSfKIvu+pbUqGcnbUoID6NLUMaQ4vY2I2xesh6bYHIro1JyF
D00px6kRq33DA74eZ5vIxwQbPSuFf8jD0QIe3kqIbHe9o+bd58VvDEpCjhfmcEqi
DYwdlxBhGjuK6S/JWAT1V0D01I8A461X0yugjZQyIvpFjrDEl5TOSIfYjTHLtOd7
ybh3vgsqOTi4Sad5kTC4G3bd189kUrYRJgVcnH1UGqm6nHC42FbcpZW4tq9kCrrj
i9ysNgheFgsksF8jwRDjrDmz/Y4wLLU/OlAHQiYoBOBooEv7PEfdQr7pgudY3C3j
GHE5DZx/QncIRAAxeb6uhvWAOcNzjMHz5qcTeRZTbPDS84162LyyIAFxABcorw3c
vu8tXID/dPuMPYP7cl5rAuOeEVp85FuRs5WEzw0AWyIYiFXErkDGGzcS0/W60Ey5
Tg61aUzi22yHSEdBasySWTAEiiawpxpdNVonI/bvg5IJPsezBhtV9BnK2yxLg5l4
W5YcTV7oZ5c+dAUHNQTRYqZlqrUg3geFkYtngeP0LzYXeWSSJaqhCFdSGx6CJTxt
jG9n7en3uqsdcxJhpXYPCQ29YwhcDs4s1cJZaC2M2NOkv46Iz31jF3pClelb81U5
opiHt0HxYjwxEsbG4c3qaVyIKsv1ZBLlehhpyU4aa4TBlT35cuNna3Ncg/qQx+Kc
181cxcGkHO++7kQgTVsbTPnDRoyWesyKolCDHngwxcQrQSzEc0PlAxhkLkWkyB92
Q6olTKhVI73L784Qp/dt+xaDRvVlcwOBva5P8e26iOkQRbaSAG2txQJAf7lg0wKO
6H113BpgBgRdr2DD/WEPbko4CsXzo+Mq3s8FA+BjcKyMQiD+gjmvdASKWBYr1Bat
W91cXlZeKEgtFDotIhMkLTnjizWsj4AW6WgJWyC49jSTCjGTjJDwybeNA67o13gT
aZtwGaok1wezOtCLPp12H4gcJe6O4vboGhSeDgB1MGrldkTBmXrb1d++YDgVnNgn
sNM2fxayb6gfaUKw4s60X0CX40HdCp7dktJKhApTr8hNaWlcLtopRUfvoJJZmmh/
j/jk/wHO9/x+5XBgfiw+XLPJd2I57rJJH2vLvIHWPYYZwI8KCaWbLT/kDmLOl/48
rwgmM9sz8A+Hy6tXwud03EnBzfg6cift3Xr3HpIkqbZkht9jT4H/UuXBo6qTBWlk
PaQeD+1ucl/CWoDosGrCyKLfWrLiwpeGUWUrfJwSMsXtxPQNR9qBK93rROCmOybD
HdONClIO5dHGvIcns7fQNf7CD6yFastaxB9yEZZzeVdSH2mDoph7v1BzIvApWZOX
FNfhkvQ1o1/osi7vRsqNZRMHlpV+ryI44SCzVswcFX5VMk5sAeZIuOrnFwRTN0Iu
IvNWhcG7f4hF++0oCqWBqc7c9cpI9T0dc/70Lw2Kj0kKghkNdcI8BAG2VV35Ew4q
Tkr+cpZ3fEUiuvIGaoLXvVY7Uv6BQj46BPhPhUwvQHWEu1DIew5XByKUDVhGoO8U
bQsQnKncz86nX+jjMQMQJBLudvorengjp74cPEKeNGDvb49ilNXoI+TGEZ3X/Xqq
9HsQZX3YJwosmM9khNE2w5X2XT2MiMK6vcUTSf/aeoiN6ollNR0mvgNO8PnNdYw9
eAj+K20C04sbAWN8jRv8pKkiNuf7N1XtTzxH0JGvmuOsMXCKaSfXa7X3cKXuD8Mw
oU5/dbpNjl8982hgZ9X4aqfbwVk/DcGNDUEpWrs6A98lwTZuohtnvyo9fI4RDFC/
iZJI1xPUCqBZlF7LYs0TDC6S6Pu5ZR2qqpTg1DXKKWzcTHEdi6czG4m+hl1Hh+NP
ALcgXLKYxtWxFMZw4Y4wzRJFxlI9nl8KPkPPM3iZpTbf+odKOK1LgZvSSzsaJYnq
tA7KS+a74f9Tt4gHjQoh6f/XV02uI6it7i3RTw2JZwkKERWRKS6XSJVcLCy+xwix
OJUgYIi7CmpR55L9YXtdc7kiBQ4VjDjaNtVAWvKTKhdenJPSEd26r/iNYhbU4AUB
PCxZMACS0r1l4Y2uGLjJY2LzlrzS2qj83WRRoDXkeLnOG4oXi4GGis4z/BLhnTWX
cihubc8b0fcY1LzHcm3zYh/Q7fB0JKutYuH4vXoEv3Pg1/QmAG0i1S68ElWnGy9B
dUiuteN0mkAdvN0SEdwAIOG9ChHG9XtjVOMYX/mmlphCUogtrDvDv9Hr1yxSYO2l
oW/p1I0r2Z6XbubKnHTkcDt2mxuOwgHt9ROvHIkKHtshnJCwXpBxLln9FVYJrTAI
BzDeGkavSYdbczxkQR2tP4iM6H1fOKz03wy8u4lHWKgdK+5IQcfDXUPnDLUYxBAR
eorytLPz45opIpgN5qYLfjB4YxweQvjX/OdvaNJUeIznEYRBt7w+YoYNlkOPgzYQ
/FNgiV0CSz5EwxzHgI4MvqyP4ArN32BXC9N5qR+O++mBJpdE8zt0hsYnhV397M3q
zmD/7D3ikAr7Q4YHiqTdzQidNRmlgBLD3Wynl3fjSoeSObQ0urpETU6uTCB4yIks
+KOIQrN4l4W4Lrb5Y7BBS9Mi8FfaPhVjrr/iYLPhj7jBXfzG+2g6seMc05nCW9/W
S7M7iUcvROYFZ4rHCLIg+czTAryjyj9a3dZQP3YkkCYJAl0G6RygkrZs0O0OOIQq
20yZKvdXaoFsd5W3+JD0851TLiTTODYh9EbH8OpKxi2vQuWRwvfjQmL2b1RNzskT
7ncirrv94mCdPsdozxwYH/YCGj3C8k2twKe6/xD1U3455bW61c1B3IZwFRXOj/x3
1ACGwziBfV/IOi5kigE1W1ZpxCvwAW08yQOACwwcwkUkw41BGSpdOD/11I9t+2uK
wt7S6ew5RnN5ShDt3zLNBiVQlyU3ic2Mjh0qYgkzmNp7Ii4VvmQntrYcbGgs9R/x
h6xr+l9fAC8V9hKOB9cnunsnu0tiKbEcVhER9sdDl6z3CE00J7T5VMNlpIh4giTa
PD+KsqwJ9fwyQrQAFP1tg+NzkUy8ag4bGvadefh4OOxSFa2cEBPACkd/ymYdVTRZ
9Jm3l63rCcjbH7I2BHINVatJwh+ny9W32Z+unA6dTQP7KB1zs1ZHhWxEg1srnYOA
Tn6M8LO40CC0Oovssh9iY3P8WZj6TtJCXVCXRoDsoLHMKGPRy2bZ/Iw59Z04+v/w
PCBP4ZhEAQO0d/cN0ReW8G7ZVMRHUGHHJxQc3G3A/HHu7m1+3p67xETE4OYSaQUf
H6kt4JcshG0ULjhs552X0q69gFgKd8QBBA1AZuItRaiMZbWyou7ulO8rKarFMG8b
rZcPTrI4qt0c8R9F7npmi3IcU2Qcqcd6s3+IqeaQwHTTZG46MxUd5xXrCBcuBpPI
rWqXmhwl+NR/wG1oIbX/T/zcF/RJE7iCTrCgIJPDC8peQ1zT4CV7PkZoMUMouX0W
coSjV2FSAaFG2ffTbmXogk8f0U+izMZ1VbKvE9YPTPhKBRKtVSarx1cTvYdm+/1a
YAKhSaplrYhvh8ySpRV60RQEmqO6IfxbfOdcpN/plHIwm0Brr1rKVph/aMV8R+hj
srCn8HWqc4xIh8Y2tA56Te/q4db1nc1bX6+/sdrdY+h+zPzUXM01FyLx/KfYJ68S
JmDKF5ex1BGuRoK7vrMOezb29cd1eXDLWKFwWCSBv0v0k0mpgNPjUhkuwt4FwtT+
T2rPpnG+uyazVCTvPTVwMii6EJxSN9c/W+RfDde6fnbL9lxTbrXpF0pfk8DEmood
TxV0tULoG5EexljGx4yZGvCLK5SkcMQZob8LApX6I0QqaEJSUNRZ6k2zTbFufLx8
wBczwPCHQgx2h5954DEm1yIIwTxR/ZcK9P59uUBdnX30w2gMCJLLPvrc/qbxwn43
hW8Gv9KrbzDKFVXqLCgP/VpYfwIJSLcltoE5L7wx48LEYHXpRs5r14V4gdKzgDl2
KgSgsLFQEZFeuZzzH2K9hjzWjB4sJ3QYNlrzYxjcyR8r8iuJYIr67zDU2ccqH3HC
WQbFqnbgRQiImM6L48VJogy5T62uQuZsFa6CNSQf2Eyxn2rkVKyzyB7vOydMw/Xg
+UzrH2+VrBrB0sz9TsmdOHRSny7COL3Ankb/JWZiIC7d087Hi+BgJ4okcXhlPviR
+Z5GCp3B0S+NoFodsG0OC++TX1uAvEG3/LnsQyljwxFO5Y/CGKZjmqA8desNeCJR
R1ME0BAkahtC4MtXKpKQ0+vk7k1OOYPRiMuMLd3PSMTVyjrPuJGt07hFuNc1kGoX
u+mYCk5DR4KRjF/oo+qwDNbJ2F0I/SbjeRDS3H1bHCaY2NT7yu1y6lbtkwsn2Nap
cZWt7x8z10uu/niERvRVyUdIVWYpbNhygFi8DNFqmilwMoQJwXXcY2kss7cK41hB
jD8voFpemlf6/yrsI4241CoDUGl6XhLMz827NOmy6vmOSHKwBoo6sPJtJAjU6Iok
C/HSm7vflq5g0bNA4FzhhcndAjVqN7m6n16PzybBOG2CDBaWm+M3NDtkljW/+xy1
iLXVhi0H3i9vjVIW9Mzi+XzgsINeBpBecTpPrI2gzXgN88MG0ElTqhwnyCsC0HLY
3UdfSfmJE15MRRs4WAov3jlekeWhUEGe0t1nq3rjI0HIIqpFClpa2px7VDhsfqU7
jl0857nzU3uFTzdcW/LWt6ZvRDgynalWvkChE7060s9HQ1Y+iB84kCw4yyDcrAz5
LBNqRlXb+7R+IbMQb16acYxzTchKo4SgcuqQd8YklSa938D5NiUfpzs11zqN0Rd+
+8L7sFe6tYAdyBJJdVPtwLOU7Rp0dAUjqhOju46+yYCfHEFoIBpWa0tKthz9znZx
VB2ArL8lXPCVeCASKpKcED8JIvYS56rxRMtMlBodOFT5kkr875ulPS5RqA8XUsIJ
mprZATqX5WjMeycLzoSe13/Q9PChFluOWH3rhgYgBLLx6YNQeVRsQ4wdHfM49w6K
RLxAYnuXuCOf/XVpKlr2TsPUizVcG0LQC2vbYobUVt4QBqfuUbTFl9Em9pUiTySP
Y6gYBx2wRLaX2Go+6/dhpwLB+YEWRnWJS+5Pyn+F8kCO+zS5Z0FyuS5z58rUSKJn
zUvoYqInZasPD+MHXyADxrTXNECrMlFdTztBw0Ay1LX2P9O74vMRPIz0zrWO76V2
lxC3frcHBahsdKfo6uWLdlITEm/GpVI0smaFu08sRSLWEAU3G6kU+bkA0Z++d/DM
SkjpnQkim5OZ5dhfl+drD/zldeSJiuAmR3WHeCTi6x9povb5qYAp/eq07OSswffg
jodzJF4stF3hsWMz49X5+cbzRbofy+WXUdtcouAQWLVoO1mtLOwz3x/5YMUhmWhY
R36WkTsmJoUD+kDg7d80rlXzBme6muElPOR7BWeKALumzjor4xtz+2+AjqJ3VGBA
lOuorP0e37YE3Od8ewZd0QwixKTqtl9i3krm6GHPcPvkxdXs5oFO+ZRHjG5UKgyO
xbQz0LaVe+HXB7mrpRZTRT2uOvqkwMz21iAlw/6LqG0nunrCoyqvjfUrBM/fijLG
GvuhYwDVi8qk8tKzw1Um2bKlkE1lvcB1Ko5nN/1EfWulNaEYUqgo+UH2i9RoqqGI
0FgGLGC47FnhFCu/4xNSoqNBkmP1WvlN4HZzie86/eBwYr3ZyjIaicsCTn9X15Ei
bN1rdLL91CoQsBTpsqyl37hAaIOY1L83X28WW90/mjrfP9YXPHPKxIp5ZajfhYT7
c1zNgoUtY1dJrJdqFnVJqT42aVXsSvDsoJCSVL/1xqzw07zEv7gn8eoy+Q21JUqf
UOVfWzhrnj6joOiSt6HQ4z0YkwVJAr4ET2StT7W1kYhXe5+OpiNtXi7fSpr5PBiI
dTPIZKyQ2sFmHyLU1stFYIZEMcvX5+5qzeYN+TEqmzGtwLG5MPmNv+aIg1nm2XL0
16ekbYqTC0wAZNagV/z9sA2Z/KUUUIjqB4hWmFWWy9Mv3rUGcA4I82Gti0rf6iyT
cKMXy854DgD/1rMmg14f6wLERcJ+D4rjGOCMtw+0oR3IrzMRh3MRUT7UrgahzBGB
su0gb6YNwjfFPM1j24ec8DDfR9T5z+4ejiNblkL1s7qllRHzZl72XcnCh1xRV49e
asY5l4jk4J8XCeziOIpMeCrrOFwE0rU/cQEaGtDdtoE/z3W6alIeragGcPy4Qjx6
jCYmhD5IyNJTGch1KUEJPaiVzm3p5Cbcv/fVckp9dzvICXw2Qa87wUVeOD/KVI6g
sYx08y0+QH4d8vhpfQTpJKs22bBiBoU3FcKmKm79Js0SWdTKyeB3AQfqHiuXz7oC
JssAZbpatQDxXU/YoA1pkU3dLIbn7bHQrPSXykA44LAh5tyLupGjPTz16eSnk27M
UFxIyJVkDbgAdJTqfn/P3tsk8RprHMrMwjgh7R7H9M5dW2lXyo7iwF6wTyCAiwWQ
/v16PKbHJaNJpJ07PGuDHHnSD7cG8eQUDuAlStkJES5nRKbB8ux1rnxHx3oeRyAp
UUMhxdbJnlQxX73ZXTcCk1AoSUk13mqmBSrpEUsIN8ix3AuoRkgvHwQ+KGuKU2T4
BnuTpwfBz7hL9feVatWRaN/x5ua2qPUsxq9lhcS5PvG4tPzFbl7M6SvDdBOdR3dH
0RJZt7Nn6JM/BWm4a8V6Pb/CKYp5fHALSlKWHcPmAgJ4yDJgKJMUtoS0p4N5B7XO
AsJ0ti0cQIcM55ESQ4PG4czh62DoM5K6i1m+YbMCJFm0iccB2R+0h8saJDj+a8zI
D+kjhv6KzAhM3fGylR9JTwNVJ8CZNIPXjWpHtDU/ubhB5eeoNu5mbDXwOid1hO99
ZU7LpIHciLpaOUr9nGTCKi/hlMHPLuHURkiAKGQDVGH23OeVrQHtoqK8zihI6jxJ
zGjhV9AX/kqVJ71teU9w8HH89nQx/aNtq0SO14IVDopx451YeHZba/D3hz9Gg97V
0DA7U5rOdh6l5C2Ee4guEFdN/4nILfIqvVLze9r+Z+ajYO10owtTTDk55WVUkJue
av/YMPZft2RG+PEAKhG5agL2e6MX7rdX0BZ0KYtX2riBPvk2aYHnVx2BQGnUs40u
1zEWfUUk5T4OpTgcDVX009h7xPTDp9ysA91kGqAcxn9tv5t65CEZCVyAkxUAkOdY
xpY5iuMgnwuvCj0LD2aj8RytFIMRaUPk5kywI6YJ3T2Jw4PbM+0va/bRFHkKFOic
2AIrY5cC/78A2aMi7gHUxp5AaYhhcDBeZk+2nyBBQPXavEsI/RV3rZynoeTDMVYL
73fUgmZfoQcovJW5GOsNX4Rl7P+rX8xHlvZrIEEWoL7Fh45go2xurbdmUNjsUoGk
vJKkvHFe1f/RxsJ1/bq++crVDv+mEKw7UGPkdD3k59ZV6UsLtxxa53ceLG5yKDyG
KxzazoP83TqyOc2Yq33EAQ6x4lWy6UPM++7wjb+vPhGhpqLF0EsoKfTA4dmqL5GU
VzM575oKfIBTGnIJgm6UNHNbIKTfyizs0eLPeuzKez9vHOojTrzyTRrYHWlx1fF8
E04B5SDOWwhi5ptBvaS6T0BPmNSDY8fwjlNAPH2cZYYI2iTO/jUegPakdyg42QMz
KbySRZ3DVMSE/3X+Z8Nt1uiy3b6WUJjnix7C7eLM9ohHyw98NH2H4dFm3indhIIt
n62PuE0x/veqazXLbhvAQZb5sf9fR8ieE/wHCGhosd3jGIXYh4kh9BEcBshWxria
7HGU/+W1b+amiiQvbuHQ1krpfJlTudOl9s/6KpL44F+0levVKwVXh01egPEkf/5j
hsPY+DxXAe4oaQSGSz5wYskgsnOOnNX+coltZb6WMZJHAcp5tgUKKFSM99szMrS5
nGZyVBy9j7pj6aV7Ky14DWHFWUd0g7viYGw15D2K+6TtNnHBXU9vRdKHUOisikiR
w+eGosRywOA78wvRHgFRB2jsV0VfK5okclyFxqEw7P2/ALYy3SUL6l0DbQazVR1e
xaAc9HBW58/9bsEvvSgFzSTQDU75kIwNNmzxqT3vdfDJo+Qg25MR8WS1GAPfum5V
A43Jd1XW9sSQJPuqikzm5UxoTnXSLimhrgiIF32P2otahqizhZGU+CqB/NfA1bic
xJZjxyJzrFTss9C6nZ1GxK/7fqEEvjRtQqD8UWQvTA4ALmU6wpf2/Rl5Sv2qrHJX
wTjEUnohhHJ+hzSBbEDnFp8Ii/X1b7obC3FVpiAanhqmlrnkNWXaTnDd6mlAX8bx
atfLAaibMP3D0DKOgtx2awdHrEO0a2tu0RhaHMv1EVcu5MS1VqwxhVyNFnY2BTrQ
kvAue+NRmmzukgFa9yYNnbz5rTAs7ryfu5HcJgnMASKmC0rmz2bXVrOEGlEtdHKA
Y3uFXXzPzhkz5wsr0SIOWPKEc7zxGcZDoR7tThpn3mHeX+rQZ6Nen9Pm5M685TyK
m51s5xGP0yXdA0U73/4VVl12JgrbXPjw6HCv0WuTyHS8oGWRJyrgE+npSRrULCWg
6BwpJq2cGTKbIQxyg6IYLSMzaTvtvsbIS4CLysbYtcl2uskBohbi+hp/Bfi+hHku
QkE3RlAuzhTnnsE+VvivypeDFwPDTquv1fzI1+05FIpczOu/89hcxK9iprmZk1mE
rnvMQiJfRRk9VuGdtukBVbJjn/nqOjFnNQRnf4grwgad2/UedUDVA7SNxWwprLoc
M3Lcx+K+f58QoPSQ0TDNdWLneg/yrfFrorz6zdmXZDsJUEZZV/oKYIr1F9PgMyEQ
ZaQvyv9MoIn7eQj7UJejZML7b+esZ6Tx/hEh9bk3thDi7mn49+OS7KAKzTpNSP2W
TZuGjHrCEF7taKXs/l56ktaXVVRVABM6E9q1CRZlXMpfawwyK74F8v908Uhrh4P5
D1zic4Uj3ROC1mgl0SMfNpBDwPuq/G5YgRgRa1nrHg70EcNfTFFwHN6pw1LH2vKp
q/w8eyBJtRc1f/WJRYDTfOofIvG1WKmhRyeXMqCmaz5G0SJTTC2e3N/fonaNjl6T
7+lGZNKHrIq199jJzE3e9qYl1E8rRKR2Ozp4RHE9zvLVZUwsP1U5ZHvwUzZocTkG
MsIajCovsS9ZOWnp3vchG9MqUXx0fkrtP8zTEWhuhvZR+ql2VLrlb2x2rAjHHT0K
cNk6YmSokdqE6DRONcxD6cjdJOPINxPpk64syCnfGcyAFWKs//5wa5HIw86xASq8
h0dkg5ipbSDZYQoSHMtxTLKvs/2T3iuU/7+NZa6vjSAGxtOqOkDkGANoUnz016AC
UMjkXKdGgOiNobRPsR7IjW5g7BE3Ly0Aw5nmysxlC8gqFKwRUzJrMsHJ25EwdIiu
oSrfzF4I3sDmnWuQHmV0f29WcGTkS1SNU0EveBAbhZEgTAqAvOViaujrZTm0Z6S9
VJ+Z9KhscWQRWEms8HYbxELlRSZwv4EIAFXtYYYuH4qeZDY1ywO9hFPerAUgp4+X
GcRei6/U/paRkbbrh/5szDGW8p0ml9QdVcbkay987KdTVqQOMu70qM0nqoWZdImV
yD2pK85bPWrFEsZDKZeIKSn8x8xmHwy4bQMRNHbfi3HWgFIsjSzuc3sCpOok0KwK
kPAtOwUOoLKVEfxl1FcS3UWknFAOVMBeKW68mxkVYWRn1dwoLduwrfwpS4LbeN5u
4T6ebGiI0+rmXoB96KPCLcfVRt/zAw66edyhr1mcTpDd62ySG8m8gaetBLWPsssz
wXN/zSbJFKvuJ9QuNEzpFKFWqdzm7EyImxDmldecWYn2g5JC3/oM00OUqenlKLKh
bq2mF6xEBeUO2j0YM7lX25zPWVXx09ok6hNwX5yCVp/z4WLBO3I0tm6HYrUJEBA3
wFDBhpW1fa974jTNdnQt3rjHuC87v44gnt6X8rMoo03HnQBfqiRpHH6Ci+PsJUDv
ynWrVSquwMb0YsZJyxkfx2bQWUVQicuW2x0nlnNinq1pMQZmvtxtGZbJdxzf+xqu
8HrthunfnCUZzthaQOleaecNbSnNXrGesin3AUrIfVzv09ad2RAMGjPMRVF46K/c
42j90C7gg8uHoSw/7prQnW7b+TMRWlP/lyKtpaCQ7MAHJi4l9Yj2zBlko8k0eRiI
B2pTR+rv7U6IacAsmsqkwEbvHWqpAY7RdOJuCkrYv9ZSUUMZyxuP1eIjvMF2btEO
cQKv4Z/oCOyqZSXi1jY1sjLr7vlnJw/iXFlceJb2Ewn37BwpKTNyz1LSS6+f9h+K
DEiVNJoRk4LxoAQUga9+QWPYX41CWOG8QigNRGg8I6ZgF+AVM+qQK03950XjqFxm
g/Fabb/XHIuPe2dpIH5sAwhDQkyT2BO+Ypt/eQEHKbS2z48pN9MIcIqz4v0DHtVe
MCccPd67jrljlP/sASZcRcwkrasDjU1yLdsS3hG1PYMl8mw0uXh8CLCPyapfPxe7
QusYHfPVrBZOOo1UJU0040QqMPNc/D6txlxvk8kmsxBRV1KzIiYKU79I0SpNSUkf
11IousXu0gQmq+aA40ooTF/8Xc7gW2zQrpcR0OXJupkzMBY/9MYqE/MNFdq5j+9y
Spv7mLlHYudvwNBkdplXz7PIBiIs8MML0lmMcGNOaMp6LGEWAAiDjbGuzhVnEv8R
t82uIAvcHhoOshrDMn5SDanSsK3+SLywDTzpWBP50cVd1nIrGLSDcU3BeLzmWF4M
h+TVKwr22TC8oS3y2gAW8wqmlbdjnBKZ3Bl22WMo0Jt1rpvzNI7ULaiR5Pi+q1a/
mVbDOmSXCWnyjWuMf3T+HDzBJ5Enq7LjDAPXOsJJJAn+Yi4DVD4m08sSwnXjJnJJ
RTaWE9SbGwBju+TZua49co37D9X/Ckhn+v4iPJuUfZedDCwY9P3qsWUp4COTeFll
qf0c4E2ynvHMzsa4EsC34aVP9AOkmi3ISRuyA4gHw1Elzr92re5dFHHavBV6Ygzi
yKdK4xpJMqukFsou3vDqIDPbRnFLz65u7rjE3YIFJAz+EA8jVIByUPpQX1Imxtcg
lfdL5b76B7XjjD8omw3PJTkiGQIQFLeJI/9WXVJdfuNImNgO0o2x8x719jj8eA7l
5NwyDPHiupm3/3pAuKxTBhGLCNXT2yHCBEDUMj0+8QqunhHyXRsoFeFo3HfwTBmi
Qr2scvk/R2USX3eqBjWUlj3SkteeHtwOSW1h7fcZ/Iji9nrRzDnSpoy8/Acd5mUE
AfUerCZ/jH6VyyWGmu2bg1V1k/EUsO892aMP1Rd6z07WLuD94woFEMbktyhv/YP7
AuaIbVN9pcE/XrZzOMnnd8GBkUjGeCEOb6B54ws8ss+tPNRZNwBP84AcPauetOJi
933GH1XANbLl+6eynDgfjVtS1JEZRhhyNQcCrhkBYValltsbd4YSAhEElQD+UvtJ
mL7CjjclAitBZr9ikef3KsZk3/no5udrqhnBxRGRRpuPNNj/ggsTU886ATBRcmcv
EwRUhRRW9pTVkIs9lFLuYC/h4IthBuaNCC5Jw+kKiIui637bbcQ/2ffl1S2rctHW
P1jD5EmX8t7oNsWr0gmKRx+Skg6/H5VS/pcaRJbanPCOTi4zmmMGH4oYVjjpHtUi
Y/Vcx/bxSgPe+ULSG4Bkw5PcE+rFJNYw75C7SrjO82pkAbYX0bjhN2rjTE2hwUoh
Pqbv98GPXgHOPaT1pnQKrauc6BdwNTc5zRiSdavmK1ffUFqZ/0NVbfqIkhLxtE76
4P1bcUxfvl9lp1zfYEORalILkP7CVs2CEyMy2pXDiLwvb3Njw281W+twi0/woV3b
vFiUVTgtOqflMLlq3VNnJ0Z3pdINqRlyNTAaIUwlfrthBhY7m3h0ljopsjI3fTXV
Uk5wUq0szWXvLP6UfaK7y+ewpiGco00mG1t7Bb/UVPVZToDJSKS+1Fh5tB14trRy
68Bx2a08yM4594FgdjO1IZgush/VqEKlqEKH+lvYC+4HGxZ+dwN5CMC1LHQYCxJn
kpwowunXazIKoNBvKgBjXSkkzdAZ/xjKD9EIcMqQ4/b0hfc/uMP201eABB8Uln78
Wn+jqn1fUgBxm7oFZBDq9MCPksNBDNCB+Us4BwYEo3KLCk6AtT6LTShzuqYzYNPk
ynkrCUc0LLH8GpYUujKLhHdTJ4sHVLJQs+x28Ksv3l/Qop1MzYSOvm9PCT7K32af
9nrJrAZXN9YvlIV0wBLSww8ZIFzvytIB84e4dy/AI1PaxdY3K9mym8TqQe0x3mhM
rluxx6CnD3eqrEkkkY4asxafbPrcRyS/4cNKW0rz/hR1CZZQvO/JqZqz4CFCC/BM
c8JxJDt/JjkcD9qbRELmTOUVgLqmftAVnwVAdbPTYWSwMBZoGh3roDpPE3kuCJEj
2TKVXxsJupJc5aatieSQvSbV5DNtbqvAMMMhl0NhO6/X2bWBgZu+lIuZiriusB8P
L9PkgMXDVXv8Kp8OBAr1UgjnyhuNhtfZOFISENTcZ/IWhR7Dpd8NVCSwN7bdeW5c
xEBSQVrIbBwhFiZJ0aaGyx9AnWQqwb1rOnJAwiqW4S+S1XdUNHAGC8/uLMG8f8DS
Dq4lND6V7TEZdkaIS7FJ+8+/r2kulNZg7oPOHUtzj5VfE8AMN2BS28UyKmscpINX
iesfGYGiQgTVBf2mRYEWq1FHvrmSuhecbueuplRTXjYN/N5b4AanOIQZwGQA5Lnq
SyvQRv6IyQjP9o8Njqu6oStw0JWS9uwH+vV3GQjwC3j0rG07hPXACv8G6RtpFlA/
lhhBz/D9VqMiIH75+Iq0JrK++rw+xB1L5ehursLu+fkWysFNdw6KSDRkX8Hu7h5b
Y1YG3zksjtc270AfqRwXpCyyMmQQo0BK2/47oc/uE+++eDsp4TqlqH9+ibuX6V9j
enFNpoZS2oBKbNTy+AxbV5l58KvHymAs2m7BfG/j6Fk/G7WyBzcPhMbyHCZD+Mph
ir9v2M7GQ3whE/6CfLp58l8N11Fj9yhAAL/hjsV/uiMQC4NLquBJ+oOkajpGAXh7
g08zXrCK/yCOHGxgG/wrX/RPQ+e9KJAhcplHRhqjzKmz0wHZIy7twbu1Xm4NEW9s
k4IY+oYD1cMEBO0BUJBw4ccqaE2gaz+rJx+vKYoQH7slWZAp1nqDpEGrUDPTWsAR
ZA8z4ojv4YHqVS5VaHa/TmDzlEncmqfWYGhk7pjA/scs1xBSNTHBXdBnZMgGsLz7
vLSqNqOMW7dPQpYSD0KVS4DpQUaso8kyDzrbg+MyotuLGnHpszgjiCXMRDmd8rnX
uMedpAZBkn4NfMCJXsf1dOZR0nIHx/EKHv26oCWegYY9yspz+PKtlvp9YG/zM33k
J/ZbhI/Q/982qTjyql70bCEUV+slQ987dTFfKiRHPOIOzCjAghbfowNSj3REIYjw
0R+2sisKLaJOYvMfDkSFB6ahBa9MkiJHonPfa2MKzAh500I0wmP9Im5dqj1GqAO0
GKxS8OC7B8Rrn373Vg59/NS8cSXOSLSHsXNP+ygy8IIT87zeMafePjXRAo5e+YP5
M5Pk9d2msbTDfcMOllg0dlC45Kr54v41Lt8t/UZWwQe1m+nPCmHVHPlW28h9ebNn
Nm28gDyDmt4LuALFzjnX4K6JPgckT7XjXP3CvIBEkB1YjXuw/UxsB6xs7owiTg9v
KcEMP80UreChm/J1Mz3OavUgNpql7yIfoNQXvP0gQbJQmAXLq2ws27PdKkNTtlxT
WHpr9XDTUyFvowRI57tr6l8jcTFE0+S+gENDnjfwetkd5yNZeCFf9fIbFiqBqKEh
yThfLB5n4RIL1EQnoUzOTVtUzwl9Xnyg0lRYfSqShx0bI1n9L/sjreAoumNH+Il3
mX43qdofB1js4x7qv6Z2CTmn3jAFfsA9yW4ysdkzfwCNus1hrWMjCQh6i9yDc0js
so2nICdXCcl7K59fDmm4wjBJm6xJO/LdjliPMHaScuy4blFwtWT3oUJzJolNX9Fg
3A4Pj8Ydw3ukH4r7b/Qec8yIUiLX1XksLxBaTpzEyfuzwqdsN/OPokmLqAOysXAb
zv29G0yHjzK2UIchoIiSInJhfj9KNnnnfkxwMy/viG7uyiTFdTA2feOYuSJGhITf
XVXEJSqdVSd4waaIq3cStKlEgcj/H6UfJkpe57v5HSSD9CWvgcWBfzaamSU2uAHB
xBRCPopezGKfAxWEewfx1xZTbM+jT3chY9zUyhlVQdOghmi2Nt60lUTPgrk0RGpU
rEd1IBHDTplVNB5D29aoaJFaVx+ov5dVuZHa+r6kXmiQ1kJ5gP6T/zu65pmq5hre
ePHld0YT9Qa1Bdi4nHp4KLILE5Rl2Owvtb1nok+IM8jXMTVDqseqHG0sNZcYemDL
Y+8nqKXNfHChKMKz4LnSfSVdI6G8u4GG2mReAbGq2qHea8GtWDMB+2xbatvgx9SM
fni1g3uMvfBD5EW1z4ACBrnipPQIf9ejB9/DLldBTeZVUFkYii9+cbslBhnH5AIx
bOUstQEVS6vB3q0StrBAOb/Q4zfnG0Ep8TlIHkEYuRstUnO/8ByEg7xzG0nLtH2n
jZN/c1WQxgWTCSb1KpNZ+ZGVT2XquZnHx8E5ACD140tsZjgL4BrlNJdXsJEGm5W2
NB2uTPbw6/NEBtaThsqyEcNTXwo5LO4R2BuXzWz7nv+x7wBaFpmzDvZn6yR3Yo0E
+JtWlD71AIvZT3y5YqqIb4iEchl2MWaQ914iUS54gNIcLvNZdgG61iIb0TybKmVl
462q2cCYdXJBvJKzqqA2tfU9Ugl/v+eJZN2JboD7DyaYxNA7UhUZCign0h1OvqwV
il9hSxF+x2Wn+PW1Dd+YGCbS9T7ElLN7elbjhqG06YPxlpWVaZrOOrdi+z45edsW
ipZ+AxFAvUWzeoYdLhYM4Zy0EHjakopLoOZbVQKWnZOsYO+PZ2M8DH8141aOrBFj
TIP4gQrg5NF12LZHn562gku7KkJ/CQpQbj1URz7AdbgCb0TD6TbzsAIF07N2BxxO
eE0Dz+aJRDtTf+N9juoL32a7XzOtGg16XrmxAMaTtjfOmCnl89aDgY4JQ8dH+211
u1YfA9CTGA/Nj+1/Kk5XmpcFE9MrCMstFAEq4b9y/Nl+/WkByZ7yzL2jcIOneA5M
D7goFRBa9uAiYRvqL1I19lsGwcKlfKXrvs1XBwPuHMAUler38XOp3d+2JgO4DVY6
eoFKEE4qkggunePK++ra1N5uyUkeJnmso4omQDKjU6f+SxAJAQesLBGDFsAZiDhN
wrnc3yUYlobT53FYvxLyXHK1cX9bGS4mITSbiWwE9FmY+c2VueSre11BfJH7FBji
ex0/zrTkglozDuMbvJEQ88FG0lLBDGLwL1D/WwTII4YaB0qspJ8ExdJV1CXqIN7p
l7T6ZD5Wh3D5RpOcDvmXZ31ITy+96JQBP13L/ejMKWsysdeMk5Td8uL6vK/4eFk+
yADtfs9jXBrdNHLHEI/lDgeHe40jAZIW9vp4teNIMO3ZJqeTe4zBEfQIzyAlDlph
XRhTxejNBDWcIGpxE70x9eqkHUDWl7U1VZc/kvy388BJZv/c0hI8Pgn6jglvOx2q
z0huREjJZZqnZGTGOGIDXEG6QJBYWhHXFhIiTgBYkdZUKEYJjb+jw5Y+bukzSIKR
yWwc2S7dDDKXC3N9TognunaoJkPr3u28krRO9rtGj1xwAKPy1eRWfAEDv9EekssB
cVg3z3ai81/Wie53rVxZQrK9KkvPQ5xsYJ4oY1NGYHWygJ9+4KusQiz6yAeYLSbu
ehwUPR+Qm1LC+DQZVQsjcZDLY6MXPAGlpo1mrLlQSPjG/wFgBMWMZkWTsadGVR7i
L2HYrfhwKhMKzo4hSPEinnEnc/6s/0gBVkZNhfHsS9bEeDJN5wHfYYTxU2ZYvJw1
Pb/SfsnbWQ0pt9lbmWD/CCsmUuYtU0k1g92BxEHQb9HFi6x0LC4N1KnTg//aOob5
IqY3xe7KNbMRjgrz4RE3wSQHbUhWWPEyGo4cCTDClr4QMktwNsP5ESFfPimf37FJ
+giofSvHw0Zodc9q9r09i9pPo7Rte+3SUFxhbg4Vyt7qLUISADif3Hi2DNKtenPm
4ibStSIqvqilgw3s8hHYgLgQ3pOa1KCUUnyWlZpEOumRnEbOVvjFcwnC6+AfhipG
2NJteVxH+fk/G8TcGfSOZKHUs6vp8XnPfdbZkIxRRO0R2S2L4pUmkmOB7eCSltkm
eRo5H1Q+YEi/DaXG6Sk7JuttKH2VpRx92gaAAUpiixy690n8aJwnp+JhdV9XxDk1
Q5W1CJpa2aO8ljWcRlDXmXIKC/uYHeTc9f7I51/daNKsUnMM2b7dctlGlY3po0+a
yjaC4sqlv3tqsvTaxHHTX2ZFEvElOK2uXITQ69KYr2f+L4niGgxTAlg2k3rIfAO4
LaMJXq1WYWhlq4H8gE0+o1qizGyjFn1sNmVbixCavnahSS/sCM0zvcq4Whcp/RMO
eN4b+y9B4T6c1uaSoTeaQdktpEJJVg2F5n2lgIQ1LlpnXYNvubdp+4ELhy4DPB80
V2nbIh6lUBCLAGT/+Y2OPxqrkKBMO0XUkXvyjhawgPaxD3XejWs07f8NGK0KqwzC
a8aVuSB+yke6d6lMhh138Y9cQ6qohIX4UA4+ZTniU4GZty4rY5QBkPHe+6Yk+Drb
WXWGvJipEipRQcQGwYFFPq1KpmqzWlIQ1axtdXhq67aKcRm1l1Npu8hb4oz/edTa
X47JfJBLBLVVr4goDjTqcsArJnFEGxyWcS3IfcQMSPRDJ6iGEp8Qi9mIV/j9E+Uz
a5elVfSiDXynDMuziepAAXO6bPhZ5KY+i74WnehJoj1Q82o1sYiGSjt7vnJbABa6
GrPZhBVN4Kak32rkNhAvqEImHkhAtZbiNipoxMjG6OxQJ8MltDVU+gQ92fZLW+sI
/Sm1ijjDw9hT46tzHUzR4W7MyYzrTBe/V99ms7TbbLw0GSNAubk4RNNtLklzE6SZ
dZEF+84Xk2J4/BV8mT8cSmDoYkDfyyQnYBEjOPgIq8h5TN20GabwW/PQTC7eeFnc
f2i2GW2Kc7i3L/bBH0YCTTh+UYGNNzSjYj5HCgDXkfm7IEbR3dZkuac4Y8pf7fTj
SCOmRcMf3Gbe8ALVJLo7wHgyTPFgpwWfx3WydiLbm+d7AeQA9JoSn7CxVhnUuG60
6IGr9GuCmq+Tm+VQbcCNXHzXkuU+8BMYziV4g9jbpPxDuGBk0SG7utQs7i3+p0YV
maIim87JW0HQeLJDUO9SSeJiAqp42b2TolM2SMsB2PfkPhgWdn+uggHbG/mzwbtS
nf/mXhHQjU2/3L4btNtruc/mWkAKUvF4KRlR9Zn61FXn+EUU6Is8vAYSwuE3DcHs
2Nl9jtX1UbExUz436Rdg/Pxo9EYR7dsfW0SCGeIMHu0O+xyAHI7ZGMKZEMMgNNZ2
M/43tRRaVetFbhmBRZHSBzUwgWAbh8msLNE49/5Z7IovMai8ff9VFjIAF8hFoOIX
P8pBRQ1c3XN6k12XQHt2BaZQhFkUcE6cXkaa0nn2tcsGI7g8aRfHdtS7Eh3syhm8
E9mH48d3k1UNWi7xln5V2is4PAURe6+UrxndhrdPw+I7PXQSVo7ZqaGEkShWZzwU
S1mVyn1dqU3GzqVzg0Yuq3D1PUTumqdp5ua5HaNFh+FT/lgcWByoklncvAxRFZDw
SkQKd7Y5DzyzIkz7JPIEeL0BGuBYMUlaYuGQqXn44quTptlyA+ktN8n/8TH8YqLw
H7c6J0GcHs6f9j/eOdBG6V2kKB8d8ANbChZf1mdC13GYtpqKfscXg6pPNUKksuOa
TBwfE5xvlpwPD4QTOSXBV8jLVucH7TF1HwHz8+Yex5UVVUSqpzhq3YGReaWnMjdZ
/DUouCpQTSqdjVOBG5fa7CGgW13udZWqKkF4VX0zyZfjswjy7fVZ/WyYbI9liW6K
LDGfLSp6De+PomGaLburfN4WbsIu6MsqKo8hkpEwxojnHnD0mwZhyL6iZmrPrUTA
5i6xfbslLXh+yXhrXW/sjm9EBx5fcoybXJbnADexBpUVZB0Yex5dsnCI0tqQSXXV
o2XvlJLNg0beiAmPOd24GMdFQyiautRWeBdIO9rbizJ6Y3tTyajjtByNNODxfxyU
DoFWqlJbI8REh11irJOi+IdCdJFKSW1CLYnavCYV1gDKCPoT4pTtJup3pp28SOFL
wlC4slLJprOVq1irKpXBr6cTs1jbAD2QaK4956m444GUc8MwxX6L9bF9lnIIA09i
iwFTE16DmwqOdH7w6c+pXJVAUgkX3e32faU8yss+zLQVaP0Rs+lYkydJTcsLN3xn
IZ+0DLUgPf2hIceP4RhmsdRnfLKA58xqwFqdb1dldXwXPqbLPeJR6eFEyUwmVtgZ
sYu+ots4vbVnYQiucSqRkvRKaYxq8X2gU/6gUab5mM8ZyPndvAal1PE994rsVrfv
hVGwwwPyieThpaDc911CJynLAMpZeslrrImGp509JeD8gnB14LSDiv9TfF0m6Sxp
VJIEPqEfR5Ll8sqLQscRTlBbgg2P0Fo0AYV2JeTDSibPTTrTRAkOaKFnkdsFN4uT
mTLbq6g3xaGC2RWJGl2fVqfdf8QGa3n/v1WcnhinyhHK7QFW55+/aSWXM26xU0t2
ByQglP+ItWHRZKzCOhzk86xIXXVGfGj7cL2YFe7UxqXUG1vyuCakucCOEhiWBUTs
L/9+GPP2cZC79raKJDzW6s4L1r2dS5RIxYoF0bwZqkD/OhqXm36baPSOlyfRpDKw
w8dULqcFQTsBPqKIO1eoqFNH3i2sjcnNivsklRZ0PF+1gWEkwteGegcMe2gQQgeR
C9kap6SQBRj4rJLAQ/hA3wVY4daMBsIX7OsvLeMIYY9zzXAGZ1vw2GO7OEPZvdBr
bgNKtjkuhQ5DWUZvS0+Iq6XhC3HsSlc5voLjHGFORQGOEH+J6+YE1+alT8E8ZI87
Qo+F6PUyYwCFrlfHxCs1lRfZAiiPKduLX3A28BwqiCLg+GLVrGVilMUq5QrPhi6Y
Fr5K7b/CFNSr77OqmoDRYOp4fN/6CtYI1LQhO2LRWK+nqaKQ1HI89jsvEUNYD04L
ERcc6hqzKzRvFDlbPLGit9qf8gjUAoGeJ7jdvvlKZS2lKTXbX0PRL9nGnQBJoBoO
Q+XEkt30PtKyxvM6iRoOaww8F5oMAGQJ1pEY6GwpFMtiyz8p3grKi1wqGe7E9n8b
B82sPE9gUTXq0EIFSEqdeBsz4nxmI4WUVQsXOCIGI+dI9a+DiZAJHYwR35mgKSYj
v0DrY8LvSw4lBDjSHxJj52+1ds1MjRmlS2Q0VEF8QvM2/rGrOGIaHcRd7DWOjjiS
NNTKOcZKfxIA1Mpkedb1KdOb0JVK/hnGALhiGVCACx3K/ykxIH9sdiBpUMtSJ+YX
gs2x/tlqKEBTqz0DfwaNNj9x2eT+34gmA+MAOWYr9xcgIuMm7ccPFu+wGmS378MD
7cNjxxzkYndyoGOsLRKK8kmwS+bvkfis2Mn8k+6wYNa+g5T9PysnSFH3a8v0LaTn
PSBsHiL+WNhqspGR/dbgk5l5HmRz/dDVFQIjVCVe/gagM/Nd7cYotKhlFrv7dXlm
FhpPaNhhjVn11AfffQ9cFHB1RiLJt4A6/uEiSTXswtFHJR5+MDSHtSLjySWbByFL
qYHi/qBXzBxI52gYo0MOYSIPKPtf20+2Gri9xTFg7lmY+DrWXVuUzFnAXAs0g/Az
/zDFtULzZGo5hEp5Z0Ysw/mFNAMIYzcWaCUlLJUv+cwjncax+WWOW9Rxt7IH2tUC
bPAAZEUFbxQFsp6cHJKkXuMCy64ldox9OBWVRwgwkGiHCA5v/NqdzpRM2mE63jRR
pskYnZ085R6NlQFwkjxqHRMKHvjFeEjlLoihpDE+EbQrfgkpdtKVgT5PwVfK1Lu/
yhMedEXctFNT8LS9N5+hvdxWuX66YeohydGjiXM/lmNHBbGCpnIPOVynKmj2m4/A
5kV0+hcoztnk7DFwm8n5YOl6JFwZncA40D7WL4Swh6y8I/MXg3hlRMS0nfxtldWi
dz09C33nc3Up0znfnJRG1fzE036XknaDJf3iB9FgrEEe10LWl5UO0HLmMHVRenQ8
h58eYZBSpCPT7G5QGmZ1OY9AXNzXVXVoRqLRJzruxpm7Y0ebCjV0NSlXs0L8y+TU
f9zapVxzlf5QCNUhA1G/qAyPFGqsD3zqyOB4j6XEuQJO/rru2G9wXZfrG9T9A8k7
r4jaIFOuSWr1PDWxuWcJG1EZNse2XhF0YsGBMge6gDXA3bPPVMacYne5GWWtiSd5
9PddBepJvLxt4NXsfxODcDaw5aXOukT82tO6yhfUPl0pxjfUMdGhQ9QYPRktbDRY
bnuaCv0q0mfxCjLjSg6cRRHRlNog0U3PAOSmj18FK524iHNgO2/WmRE04/exFdhe
havDz3MhoiZlvH7zsg2YjSCQGjRWqRy8RhVrxtDIY7r4OLv5iupKvaoBcWYFcxSW
1BRZ7hcGyv4AgA6+TCSZydMJV/QMlUonKlaJowEso8WuP0bt14PvXrEMaYBxxiQQ
/oXwGZw8UglcuBuIJqrTH24pg5pWDNKfg4srsW1GEOa5s+ckTk5fu3hc6tgIRVYo
1gKGP0uDKBOBBQoEEYmlHcHEuf837W1EbvFbTDK8cKBlqQS9FNsBSYjW1hzBV9m7
bFoEAP5g2JrqTVSZmCBnCcUczgZCqkTdmlf5YHNM2DM2EunPYuxqTfXL0J9fgxHl
xyvhNQrw82CdhS0zY6SBbQfqRHKDLljArGqGSYNJXnmJLC3LFE9eBbN46XVCYpNY
0M21jha9wAhrQ9LUuyjxnfvDBpoGHyhWXtjaKT5iZXCNG/CXXlZI87qBC3mvBOfY
Nta385OKeApeSoPXNqcNHUUmlL/3ZIahBFEu/kkr2nCqf7KJlTvqcDcHslTXibY3
HTQ366r/jfrDN3+mLKIQD6PfYFotOiS5r9BwdB06ntut6B+JJyAuIWSGUGx8wLXV
Rfk344ifXIm1/YGMWKw5EsNnsyvqPRKM1cYlFMw4Ltl7iBWt5fvGxolQ4IpIMw1n
uo/y6YSfOR8nZR1XS/BsHoNTzY+9McJNZNk9WE81gZLuz8CZ0bzvcdLpOFw8eHwh
bB9YTMZTTrhKQ8Crk4ea8jGQ6RuVd74yB8Xz1ipYpTbnhyWB0iCL/OOLbf70H6fQ
96ffGHW7i+Lp5brkWmwme8SwiEFPPEJln95VPR5bhs/9Os/1aRxRIiMCqpZuQfk+
pDzFsjBrYDSw+XYKh28BSsuYFu/3S0kmkW/ZE85CcXrR4FovXyf9EAbI+lWQ7giV
nCskPezLzI6lYfc5m5Mv+WRiJwkhXYzB1AoOBbrPXmjdpD7eWiCwNSmLsKqceKdu
C+/EXZlNL8Z/HYFSnd+vbsKcpbsVkO7hhdUEBYPiRrlmG2hXlACJOOyTAg1vhwxK
nYD0wpG0g590Tp+Pa0dpRNHQlgij49cBmlm9cGSu2LEV4+/D6qkKfh8PsceSDaOy
wUxrSQHqPStk6EjmIrYsm68SulIt2ytOZPnNMQsrj33Cual4vNwqvDMiWm1hhtj2
PD+2saa5a18tA7eSbLcNIvTAJ727VusPIqTeyksL6uB8q6BX0OmGfQ6jWDq+JGa9
R7fcoWGqtA/HeWiF1gvEV0siXX/Tmnvs2cJCfRQnrPTDLtLPgBN7ynk+wb0K4X1I
2SiKTqOsLSZblbX5RMXa7FzWDA2XQ/S1GVfeQWsLEo2Ni4iPRmWYoqW7t/zCiUWR
EKVu8MGDvVnCvTU7whm+NRdrMvlPiVfFMKkBG5nT2TGLM54MrS/9i3Ai5JswFYKN
peoyRH/sARH14NNEG6JQ2uS8DnlvIH6i0nDToc4Ty2jz72YV84cIDwrPe9pexo4d
Rx2vNIemRZkJ/gNMFSoBxvPGjvxgNWQh9QE26T8iw6x/2S8bJ+IUW5NcyYts+xko
cWbuKQCtdHMemeAwMeXkCUJDXx6S4GYz0zyR9rMqhcYsrFMIyNjK3ywZ3uWgEqkV
7FH3YCT+IrBEdahMlMckRjwpLX4qrEOL6UqL0HMxViA698o37pbkNd5tIqaKOTza
oxToV1LvLW6alObiUvgBfoh6gWrqjG74YJn4zdXEvTr4sc0bGqvbxqROr4asZtPG
BPTez+WxrpZjqfneu27T7CkUL7iEji3qtwzDm+P69Y3+ckxTkeY1fbm7AbDDJflf
0vSyz7ztx5gWYQAstnNk5olZK9VQe91LdsGstIteLGbyRO2VRGfSkGt7xmQNQSWa
T847GyrjxaRWhK/Hnx1Kbq0lgPF70l0ZoKn4y0RdE6BezQcuK1WTvfCS3Ht35UIh
aaRYboW2XCJAItArPv+MMkVJEDOqf0X6VSVXUt8Gz+cy0KiR7zmF13ugyZBHoXFS
QjK3BaTWkISWTp/DNQKWDl8TccQtP5jT3uftNqcpGj94w+rV1SYb85Hc7ISIMTd2
Jbp2UGLfNNuKNv5sHYtZ95kSIQPKccBx2ObDeA8KHDorm5i+ARdqd+oom+kK2L9E
k3bNDZm9Byh2tzJtMBrDtzeN0OMrH37SYgh2XTw8tEaR3tFvTviomjnxZglJE9cD
saIYImDQVdHcgRCPwhCy8WnUxZgmH0hBsJbT/czrDBY99U/YBICdKiYx4hU2p8vR
MprKaCW2IlILgMENs65aItInLfUZZuekKFdKCkc/pW8xc2iOfU/FZ50hWC5A5uX+
4XP52LoOymQwb0h1P99h8PImqbZ1SzJjs5ueYLuOwHmHf7qDl7Dhk3wjPWWk5B6a
8cqUxeFGNzpiOgahpp41FcEEB69o+OVMJZotrNURDryW5lfr2t3Mx9/hCJkGVbsk
pqPgeccwE6awG7/OTNN8E8i7Bf8bHoKDilo13W8fsoCYAuupzfy9sB5fwok0jMcN
in53vExNbVcNB3mo9CfouN/LIPGy/53TUaeMUUKAsTBlfyguaxhf03ysGqWPAQ6Y
go5r0leedVBfEflKLzOgGy7ROzfHc+4F4SNC+da/OrHVUOLGhHQZqQRdRFYtiInz
6FpiOW5O614F2q3R4wg9ETCXc42w7TtEX9BVE6CDOEa5BuZ1ZZGvxW0UYN/20TRs
ZjIJPKonTOqBPBPao1QwUfY6qCYM/TZ/ITON5/J4rI1W2DVio/1QuyOM4ihL+9le
zxFsGIazsM2hS8Hx8GiZKGM576GvOI0Dw/XrExPiFMMVf8LF4IxTJ8Mg2jjNJ24u
KCEYGkL9Ce9QZyusF6T5junkDt4uRRLnZoqwIrqTkaJ1dtEqJL2Qdp2gi3iRYYeY
ChZZBPbJ7KNe4XXUL4Bc+hoq4Ib55sAZAh0nEiArLQNkpFBY5LzAdqbjYA3z+4It
GvZkyq+nJ601tzlKFX9OUdrX/gk2Km+JPeydZk/bxZZUrliXtZcK+BK1cSCaDxaC
FGqI+RnZb1/eoGIgSZt84QZr+j8RB79rFIpkX1dzxWlm/sjlq41uRod50Dd1/ni5
uWem/BfQpYT6xLhxo/6mwYCP1tAzOmdlbZTYIrmZ92o/d3nvGDnb7KdurLyDQSVA
vW7gLa3gpZ8C2QYL3VIk+zk//lMiRU5PvsplhRiFNfSyAMqGwlTSBWKUcy4Rb43O
SEAC23zdNs0uG03a9umsA9tWTeClwwXmfE/1rrU6y5HHYvTBqPZXfT1oqDLUL9aA
kdbe9rV31Bddee6n7wVlTwhKNnaRNRZz79S/9XHiE9Z6ThU5pJAGnYTeq/GynFcz
OAcm9o0PtpUViXo2Q5I9fxBOtpqhy5D/Acp7xhWTWG2Z6hsmhxb7OFe8sxdCYFfK
vbvieEtQ+XBJ929fTMSCVKRLCMmLcrRyeXinV45nJ+0Ys2ngm5uTUwP4hlG28oal
aIwV2eVv/Jj3+PNOoD3D6KigdrfYRPY5kmXnKJkOs1A/Hq6hhPcYt5mBnherUHTu
XVtQkNWmurFnMhP4KRW2rWiKxvxH2Cci6Fruen2vWVM0ynmbMKI6Cuy3LttEvKYY
h/1PDTjwqeA49FccsLc8dCw6gqc80uYpzY0XraFoBSBp6p6AuqTE64L6hsiGCxaw
USKiNFODGL/SiDxfLy9CcdKHnBgsmuwjObVC/GpD8CxioMucnCGztiQFPDdNVk6V
6o8WlpCSvJPev6h9TSLnOH3TdiAr75ukTZcXOv6ZvF03xvnRN6HXxhg5G3sV8MnQ
gXbO7PMOqnAGBgcyz7Vm23+BovspwlUlHzwTpsDCnJNYhzyfmLSsIPzkOrcUC8o3
CDvbPEx0z5Iikz62jn9+0RWg467PPiVzcSPfzM6nUOsVg6CwWWqcJvAUvdm6sI4T
LcMbudcxD6adqwg4dNnn7Kaq9DHmIb6ZcbJkEYIpf6qyRTb+qxQKBGb3UUfFbciA
iMeQ555hRB7ss+qmTHsSkRYwNOGO5mCgws+/UesZRiDdr/uGNncKMF2jvmMr/xtL
tYAr2w1lOp/3YYYxgZZ7xKjWJhC/icwSxM4hmDS9Do8S1f4SJujoxVJ0zFVNin8D
kW4p56MDWnXTBDuvExrbMYSxHN0RBnkFyz1RGmEcWVs6bb0/Fa/27mGGRI0Fh8JM
IsWRSe/aBXaDDY+w/TiqkGorLOO0lG33Sk6zFh12eN3CX0Q9cbG3lFV8E/CBy5t8
asNcImVPECle8t4Vhoeijb7wmNIdNZfUejz00VaAWvyfYEnK3TzvKSw/HkByrSYa
FxirAaab59Bp8OB4RPzucwlQ0GOinHZmFrHR3m7f/qcHYwixOCC5wFHtQ/O/bgts
bslGdOAr7lts8qniei8iz10tTzDakIZpg3WWo4xxGdq1ehl8Kl6b3Q+Nwd+83Qmp
bxTK0XdSu5kklsRVutNvXfrN+tMYejGqSWRAfRkj2RItEEpF+7kWU6HbKlIA3XVD
L1vpO4SxiZ3B4J5S/e7M994Q5Q1C1Pomv8QvkHNrWq+oHlqDULQmDv32QcECahiP
eckbESNkNvO30SY2iIdRbyZXAA7EiyhIAvstLISMNJdn02zjzbrAMxdtikdBW59s
xAk9sxJAjwTc6iNkHRaRw2aWnGV0DlRArho3UJls5bqHMkAxF2x6ZCCJQ4TU1Bjs
8bqKJl/Cvz03G6bK8+fcNSJzr0f7kkwpiQ01H3kYbmzgwFlTtd3q2/OZkYe9+GPa
Y042oyCVfxBvq+xetpm+StbfSG66L5LEYolzkqp8CqT1PHUjCHNPaam1gxqFnEXj
Ot/cTgcGxtPOq6r/x8t3O+arQvir0Reib+wgqdFxNjEziSAIVTOIvBGOtBJYYGBq
AHxnn3ZA10yes1CskYFlvkX0XbgrO6kLkoFj9P9OX9zH5dgIUUeciMNy9K4AcT+J
Yo/2RseISsej8e1zLFG0Gigld0Jq9tOZG8KLxZROo9MkY8ewz8W1O5uVw0jht05+
W7E8iM6dNad6w+gBrIvWo811uoy4V+pmlGlnLQsFapT504S3e0BgooaH0rbckThM
sVlJG70TmFLavBxKwg14WDZqN8GsybS+JTwh+DwBHeKHpVTxz2V41cI4MYYJwNWf
c4ROY6SvfENV2tsUvrs6cVUYkdytwGAWDBS2IuzxbwDHNEr8K93JbwrTf2Zc5xMt
sWA/ykjJMCka4KNjblejJwoxihYk8bbEPue/yKEHLRxXOwhA9CUBk/lmHEdJi2wW
CuLJy6FCrAuAbExi8Q50URMg0icwpCaPTHO6V8cPz6bfKiv50S84usA+wnXbqlxZ
Ervlji2TwdM7c/amo8h3xsdGdbJ47Sf/SAuOMfbU6unpC0al0U85SJtgNXSaxTnZ
k+Er21EBbNRdMZ8Er99ZZBuT/xcKGZxn0FVImHGDvGo0qPe5+MDm5nUOdnuntlqY
kEGTlQB8flbaOH3EB+cmMZQGlf6c0vHXHjNPE6ybiAWtKO1Tt5gmMJy+KZys6YRr
LOvqnjJX/WRJezZE67jBybUj4hclZCv3lxOhHx6DEz4stzfjc3bjFTCpLBZZCAYV
E84YBJOCdihK8UwRe6ttoap6m0e21g9XdHELQvP14YTtPA1hVCgzBHMqPi1PFHWn
VN5nKs0Da8xppZ1Tx0Jp7By2iljKdN5S3tyXgFK6flf61Qz4wH1vFCTdyCb1Kf8U
TdyKYwi4NV/r1By+53JN9t+0ibIQLVkntt7k+5oeYuGPTZYNAdAo5UndHmTby17Y
zkkulqoANiYqdZupMSdhgKu6N4JvgprTi51ht24W0qmabaF/McKoD/B+eTCW2hY/
Jhx3LgMdjFInXocq1s7FPoAoWxQHRCvEFXwEkkyYdUD3JxwLCWxCFrkW3Wy83GEH
XZ5wKrOapqaWskTwfa5ShT5do1tlTvI9uPkXgJ3I7i5bHUpwRMyr4UYhthX1gLcg
7Lm1lGtWioGE93TpTQkMJ2rIaBXmz5RVNSEOM785YihF3zxcSFhImlm196+vi5af
ImZz+RKt+4J2VPazguvG4/bcXjFcQ9eK7R/nfhXINgDQVswyegK1ixn1ICPg4qIT
gqZf8ggBh5/+quO7vLZwbSr3OePwccxRw1M3ZJyBsNIU48S2tTmU/u42Y85lWTcF
iOtukE0EYROW7lZwv2c1zraAVee+ydLiypm3DdMEyl/4ILaSA3FFxcVyzhvedvtA
SS6rGHIllX0j9CBnAS5jExpBwxTjU5fiREn+v6a4qos39SWL0z6Sbz13pvSK0JO6
b4w8FFBFUuOXQ+mNh8FqmspASO1iLJnuocnvF0/ng3jadjv8uG0CNOYb+D9rCafu
fAd8v08GNApRbyEgsPis5ErfSUMWoP1XUysd7k9IlpqvvJrwtEHcTXr6MCYuJUxb
YgMhxyd/siZzV7fxd9/NIXH8XB6A8FNTq01C/trioojYsMSMRHV+vbez04ZmdSDR
CX/wdaX/7PhH/+OfS/Td93fdbeU8QonsVW1ZOwzRaJz2x41mWfOOCN2MRTQ+85O4
lRA0RYTnG6aQ8NB7WGnW5nIdyyuYc12BY04X8WqCIX0aCRhitZd84iCE7nR98VZR
jRdZFJdKWoNLAoN/uaF4Ahn+udrSpcZNLt2qyiYeXokxJPiwev7xvEGHOgOrzy8J
ltueGpqUhACThyWcU5smyEFh/wsRW0uquRQ61hPBL0alRfrcblrz3TucCYKttiYW
SBIXzMNxQEBeInl249U29tQJmo8Plt+qF84Sn7jEieKs9QDcV+uOWXmkPRhlrZXR
ZfGHUs80kM2k3ZeSzAksv9anI3CPUVbGM5QsDCRZ7YBIq0kEr4LYwiJzomSR+Wxd
funPtYpAKZtW9THJh6l++NtgjaU4LP/YOTjmGY7GpDoL+2VSOVk2dm6tUPNIdKA8
YBdJWnYktrS/dI6rHesZ0VjCfUrTKLtj6OtriZ8GSUDpRCr/gf4D8l31vXU3im6B
sHOWze7uQfLl+IOIuZSbpypPbE/wLNMqEN0QITp6aLaLRvWLPgkZQXPVZgDuNjEr
wlpthvXQnm4sIWnDzJO2N8V7JRG04kau13/z4zlJInlBQaErecxM9CkVBvYgICrG
Au5In4jJGITnqK1NbBrBtpFkqxz+nzH2zF5MRxRzMkNhMn2SXGAYjb+i6Hbj474S
sZXX26hnNF9DtBud/KCh3ulERBjwLgVQUbZFD8nIkjmrKClE+9XQ3CrLkV41WKM4
cwl5kiZzfzty2lZy794uZOrhOepTvIyEtuU3tPD4sbhvxqEQ6TR8G7f923+GDpdc
cXCb4QMlM5WYt+ifl6PHJlm+0gLNQGhhKoTpCwX/zemhQCk2ciq+ZPoPp2UJtKXI
r8vZ3DlIDrdsweJWp9ZHndRx+UdwEAFfbQWOcOAC2Bas+VtOOIQtTAPCUa+N594K
DNWPWmDbhvuLx9zOImhBilsgFueY39pEe9g71bvWjuiLLuE+hdZ0LgBA2b2VEkoz
/liDZDb+aiTL3ewMQimi5EwPyweJH1l+chi1axmy77OXX5h8CNdsEN1ZtGw1g5ne
XzMpcc+vCXyOI5ObFByV23ln0kTQ30kcAER+K7rgoekA876HtG5yxYWq6VvxjSKG
C3nnBGkfxI6ScrV52tuxDYjGm6sc/yqX7Gied7h/nUX5tEM15NprS8+JZlyWBbnc
azo0P70oSZsrQ2i8hbmorJf9yTyxfkIAOtsQ+bKsFLr431lEjKa0QMy09O6p8lf9
JfQqPdLZYJmRK0i4vi4uptB69FjWFBgLPZ6eZlKLCt2RWkVDhl4dXeHLz3TRM44I
yR6bXcZZR5dHJwSS8UqIfjzahJj185DMIMkeIAp/EkEo5XZoOFA08aOXA8gIkW9J
0Y4jmu3uSIUepf0SfSkkRDX0981pHQRjbJyFi5z1RLX96wZ8hlYPJ7G4coirGdEY
v98LuoOuNDfm/ljNMyN9G85ZqYhlxRF5Ho3oU361KmQ7Dj76x1t2nkKUzFzHIGE2
7sn+oqZH2FIpn3OSLZwof5JTtCJ4zbhoE582FHE/HibyTsKoFInFjrhXKanmTJ0v
8ClhLTaIk+rf8GQ8RcGwwWYJTobt8rst1fnWSNqClfys5efP7zKp8xuaQDFwLxpH
nzrYub8ulQYZFYQ5MsSrzwPa6/lEtYCwBSZho/h/l5tf+5K2JBGbZrgFN0duIqLS
c+rHMC/yYIOhvQ9pEQau7Wn+6LnGoPaEbFMs8w/6I2c5JgWJBStZY1EMDaNGFDRu
eweI3p0fNtn4uW7+yTaw/UnDhBAvGRw5lR5z0BsHlVuhJMilAi9dY12Vicj7N3Vz
s2bx5PsPEE8JSP2NUY3N36oXryzKTbmbFfUQXxkf3FhUVN2ggj12IBMvliifSvUk
UyOlFI/5wtsCF/E6R9i+j5o67d+89jmbJ3zOzGWdmtiebqadRwnqkVgb1lOTk0ka
tgPQ0DGDC527IjQwisXSljhb1gnBMl4ZG+CJqGFlbuCTYkWOhsVXwcArUsTvPrKJ
XG52hoYwXmKxSyVfzFUi2fXUtlCvfmOV6Ix4+pf8SZBeJB5VcGVhgU9jKd6m6RKZ
UCTP9+c/7Opu65EE62JuZfttJhVgvP8rBuLkmk5qEFAp/+5QZTQXjv5DDNvh3KoE
jh6r4h889Gx7Oi7eXv2AQS9/GcbBepIbzSKeH1K4m57jUqyip+7Kwr6fQSeYX5gM
872kWY4SBt8HWOjWucWFUX49Lp07K4sOr9lnYC6A3mQjRDs4Z66hUPn+c7DMXlMc
FM1LMOi8lxpyotgbfJQHUkfzt1e8B+ee+2CU3kmZcmO3M/GFc4PkQx3rmc1KgYHv
9RP3Qrrxg8UsrCvn1+0Qb3INlGmvyBHelAjTmKMxPIuEstSYP2CYbCRjFiJGg/Z4
KHl4dqZLteg+xxVarM1rXc/3WwA0LCX3+v7vhKkv5v/+cYFfPVkq3k1EUmDynz5K
OcAJra8RD9xyt+R2RfgbOMiigmhdluw4Y4xlEbEWRQBIG3RkQBGr1H3K/ggoFS8M
IV9L2lmqmcLjZ2ikHPtfgYl+QUQRjK0EpBE/UGozvbVZUP0g0V4LAS1eddIyWNv2
vx9kiXEy9IlUAVsHVJeGjEWcuoq4hs4zf+yMRxcHoa4rbX5h5plJyj/iQ0ZJSnvd
Q+MFoo6AfClKAT+W3fTPboUupF9GgZHeoXmDImaHgNsl9+wXXwSXwlajfMPVS5Tu
kGcnVlb7NQ6ouw0zIpossKXr6/3eSaTdlCfJidM9vSypzufwhYx4lDNFbhAQVr9l
a61ANEztVj6ewP0628T8qABscuNbs1OesPzXT2RKDdUPp1JO7x1lA6rHuI5vhxnt
6jR1X6W7q14vCETTpsU7VXQ7rI3DNc04RNb+6sPg1XWXty5BOsxZcFSW5Kbs+cYv
pKqVL0obWoWamuzW00tQhLtG6JelnJi50Y8qcaKnUou5AkgCpyLTuXWwDO/d/S15
/kLBdrSPyGR3jeSLkK5xX7XHvD8NWS0RU1PSdp4OxhBGkLFJ222wPGshkTyWdbx/
hDA53wiwxowptT65skX3GtdRw8gri546X+Yi/zaqkn56bV3emIz1tZy6b9P+VUFP
3F9SMha7wIYKH6O5jCBv3dviiIDib+AHsED09PfEzGxF1ErUz6HWQxYBPgkN/VQ8
zp38MheNICprpwQ8pJ1/J83YymjoEiQHr1u8Ee52GYkuhthecL16oB0aghoN00O5
+qGvghyUkK9bMi3436ch7g0SjXiP5yvFqwQJit40KMF/yqMUHE470Ydrzw54Tn+Y
MpX9IK3mIOSD6vEEKKPtBQbWEBqN4edSHxS8gakGePK3cwOGkPitJA7dMTP2jTRs
I/aO7x2yXD2ZVDM3uEmXslxPTA3n+tne+W5ga0xw4nYFf3ipKDKcehWyARv8qYZG
eqROknDxmw6aNuWA4CZ09PC8TOq6HaqmdywQ53EnWV8GjGvOV7aDlsY7AijwiosH
l8aUYfiPtJF13sTkULMYgrI0Bg7t3U7gjQLdCEGr957AFIplh8QFvzbH3JoH+I0l
tmJCLNcA/fj8rBeK3eVUvS9FfLOx7X/f5Cj6yamTHbw4aluMOrz+6myEWTbH4QJ6
PD82P7I066LzfqzS+FvkNbRVm/OsDnBug08M+Yv4oYLt8qoRPYH4nXZRJ44ZfVQ2
HUNI0Wo6SEKgMk9LTShtIiKLfwfvEtOZPJX6UUpijOAcQbRXoIpKhmMBrApX7ntL
3ECCFNQDXoot/Ibtrb3HiM+MscvQ1Il7XjJMAYPlFzZTISkuWnFDxzI9dVl7XYgF
wIYfZKaIEETilghpEeu8/zj00Dql96BUde4KwA0gCjRqhZP8cEvwhGlyZo2IGmBo
mhr6CEX+t8UP0WEwnc26eLtuNFitfRlx4cVc90O9UIqfqc0nallLGMDMGbJHdjIr
lRf/yGZ1mcEtX8mNb6Kme94pFwIRxK0KNcI0ZgS0dOCw+ZV2EPYJ2CRoZYrHeEdL
MAv24QitKK/7iPiw9YWDvUEhOowck+WUmCC7ytJ2GbMS/ydmRblI3DoiKf5aDb5A
WTSjB7ThDr07AjpN/XZIUcqzKPfB28y/QCk5k8J+ohh6UCTvIV/OD+Hcb9Rm8dGS
MJEAHT30qjJBEp9DW7RVXwfZc8LIAX/3UZ1nwRtNh6e4dvGy9a6MR18nvJhMxRew
VPeyxt50kG5R8jO/7CXNSJIgMZ1TG5gMQODnuzbTQZxvnLgKtXzofHuObI3ObF6V
8sKXv2qC8hw8dm1ZCJXSTi/g3YTG6moNRlMLb+KyT++sy2hlo06ztckJNdOhXLn3
fs2Ta24yloh+NXao7wPgqXh8yzymmhmg5sFC5DurJ5qkXEhTWNiekhWlsykFiP3v
V4MDD838xWjA/PNeF5rPDjP+uaQ0LD0otPlz2l3cNFTmsM53s6sq+j9G3gcOy4T4
GOxJmwUu1LWuHgbcer5Tiz9Ce8Hxg4pYvAX2YCYf9/fDNqGnuFZdEXjyHHxIkMvA
6KkiWNITk22mnRBL1zERuFE4NTJQbaDHYlLsVuyk/iqKvq6rBNp4E5wgXKy7p2BM
Q3Q5FWPr5oWBxLwLiTlMcPvVWTnovBhLibnSZW4niNJ3QXg+X9SHGViT0wfzq4Qx
Jt1ficyCK1iHa3zLKkj1cGf3mFGqm2o6m8fh2VTblLLNs8kgWHT/uz9f/He0xSqX
FwqGnMcI7OCZpol8cG8hsvPc8CrLp/qMBr5y4uG5xhSlQ+Y1R4TkiX+IRqy5Zc5f
hRB7EkZKwRawJbPfsJ6uIu1N75b1CBmMsUgdCo8jPQNoGwIKkxV4IIJB+rPitQ+o
b9lalcrmBNyWtMHbKneSuuMt5ijl2+0D2NT8g35OCkbDI6a/xNH18lTBAG1QhizA
yx9XZiFap2ZkMf0u0vpNWEC/2dG11ljuHa9E5Lp3Iulew6MW9r+gnAi5dTzZ5/C6
LucYa21aqG7b90JB1osjCHETkJ0hdIAkNPCaKkHKLeV37S0SRofayAyusGbJeJAQ
v0F/zjUrJ+aGHgYjxY3kzRa0ZaAkPs926Ci3Q3nkYjHBEimTozNK6FU3aSByBEgV
y0BT2v0EOFOsgSWIqt1B3wrQOVoH+Djogn6NNmHVW3OicZ6JcO2K2y3WGARTkNNt
iBXt45yycYeZAMvMQZkJKd16sOG1Ta7Pb1OcDAcoEVVU2iajeCG7W6oQ1Dhxt9t4
3MrT9RTv7Trb2NwL6JQSh1IsfqjkwrOBBpOEqs+Erme7ITWWfIOLokJrcz8xAMWf
4I968bu76G2mSa6XPmUflN0jcnhZZuINJbwSnRGyDuJMaqh7vbg8HbpJZT8NHJVH
HdsaoQBW9lBb/qVq2PimuZRe/PGMo1UuM7Pt5N1mOq4yvsUrtchkhjonavjRJUi1
ujVlEmncHASIWyVVYI7p/GDb83GFJXS0qPBshcwprABkYAbioL82mZtR/ZBTdgFH
V5Bp+mzPs6WTFXe3u1gUtKqpfzmBM+n3/wDDpv33JY5PcbH6tcIgrsApfD08SzfQ
+rc9UuEYkTT+rJold6alLyqze+aFeLhWp2vX78H03g8nATiBu+kSI4eCnPDAb3lS
vpinlSUxxk9d3y6+Co+IMx+HHaMaFpaY7HUEcX5z8FxYgadu8jkaka7DaLRH9Uuh
lrOePbM6D1ulELVutII9kjLx21YJqP9WQ1MoofxhshxMlD1tPcXeE+j6ZEjN7UQi
gvvSjgyTUQyHVfiYVj9IZb/BnlPRZqDvhnP0jCPR0PnivAKSudWtCAOHWulbfV7A
YbCg9HIZ91Q9VpxMJtSZmFFZr/OrdDjGQM6P6zfPN6raboFaFMcDjpEjTq0mMqM/
SNhEcpflF//p3YYNZ2La+ip59xKkENXmEoOu4SbebLhyPiZYb1nQQniI8vi6xvPO
6vBfJuz9zDtXlw26EQZCP2DhUfPWlTPPfEMtBy2Cv8bN53txFdUJhBT9bnSF2GYD
Wvktpz2bNEdv5pywBcIaC//KlswG9jlIqJxGlggCbpPeJ9besLBQJ/8nsXjnBV4y
eTkXze4PE5N3trBlnjGalTcZ3gOpJPxVLA0sGSF8LDlKtaC0ZVH26rh3iSW9cu78
R/sXlLbGtR/G3TKcJRGC2bTJv5irCLIgLv4QnJS+IAABiRpME6OGYgtdIcdesj6w
MDEbsJeukRVx+e4sNDiXddUtT/y6Xy588eOJjp7nSEFzJ6bhIVDGKL50Nq47gOGO
Xj8dTdqlwJOf/QJp9MrhIYXf9FkK3krfiBWOdwXJCOu+4BWjITpHYtRJdnFE7Fw3
CvGV9XQsvnmTQOC0eGt05KpconOYQ24FPqvLNIGK1Fa9SQimeM/0mgCGpR0feNpb
lgeQ2IsBByWgCY0f2eyAaWmqN/Sj3ZiSMPFvJReMs5oSvY5tzt3YVHyYTyAB5+0L
PRoL7q9I1NP48ojiKdFKVKuubNUqLhBtIkUWS3U79/PXinXT/Po5G1+hE/P8VEEP
zD0KkbiJ2Pxn2Ozwt/2/9d4a+fJGxL6F5qwsYy2i3PSPxXMijeo0rLgPhu6eoCTy
osU5BC2hbwZPvwzTrPdIiz6DrbVkGYh+nhHgkRe4YfjEhiXMauURBCsUlT0ESlok
vHHxG8A4im1lMPD9yi1jw7y9YlesEQyUZEEWbOf9CgJJ19YYBKBU2aAoOCZoLSb+
lxajUsuQjpKM26lL4s4lermY+cZEbElndZmnyI8tpF3CGmX2HBgvtTBqsBPhmlmI
jrPIsqX4pM+iz8nubwCjZ3BHcENeJVNqN99jl6i3srxt/dwY27+pKVOOToes4Qj2
J/T4UExkuJPu220LqTF1VWZwKRaDRkECoVKxfCqM8Q5vuQui3CqWgvMZUCgrOF6U
m2jaBRaY8bIMOJ1KZoSadFJZ4oggSd8NNeK8IxNlIdxtUsW4PIGfdhGkDVaMJkmP
pyaRNqFKhxYlZgF0p6trfdjBtj5fQhaa6w5qeyochG/9G4dHH5M6rsu7FrjDbHNl
Hq5f8GiRx3FZ+3ymGhkQM6Az/EBdugJ2Qfz4sU9AR6Xz1PlRzUU/vZ6DsSuAHApb
+WGUFaLs1SqO1lqfHxitBWd4YqSt5WR+P4WOh1oGS63vkyQ0G4Lm18nx3U72R1dT
Kr04AvwijqT20gM0MUhd9BUHZIf/RoiLlb+Ts5gZXeYbAnly61oXSERNJ3D3gb72
mz7IG5SJxAIcJTZNCxDEXCtFRaBRr3L5736zwZsIcNpVmkq/dHeUfRinDyzAPDSS
vrHZwjvnDxMgILDnKG3Fz9RFlOv3NsZhdqvh16O7CJaQNO9EGgI0xBFblAeCrzgZ
zupT242TjtB+uvIkLcv1qIUTNKXOY4k7pmk2ib4KTUQtBftCP0fyX+/7EekF/P1p
ocf1WVqt2/fgqiNAya2BeqNjSivxZ2gfS3epgX8pLoSNgU1e3ue289wY1Ddo5WYg
XiqKz1hrImYQuxMgbmIPRXIJjucFzCYgUOwLOulWaDjPFLoZx2Qe0qsym10oTD2X
YMut4KwkPpDdn2v9K5WiIyNzub4SiuN8C8XTSGuszRmNh1QdipndbM0FEM5F/M1p
LSguR0lrw6BelToJW+nuQ/UhwHSTgU2NWk600XHPIQvM2DKldA/6qOUNwaKMN7E8
fHdSR6wY9SFQsBPqjPSY/HLxCxXApNVcz7JGsKAaor+Yrehu8m+oa6i6O8wlu/Zr
7C+HPdudOhKwmVVslPdUNrEkGV9MrZGPqYtgJcqEd5T+uI+2R8ATksZjQUXsusHQ
u2hP51aLDVSgMiJwrK89NQJnIaUnuXe69kyz0Pncdh+MwtUOF90adAo+vF84/BpX
IXCU86yRN8579744KUisToJF5AoNCrHBybn83IHFhfe8yOrw+rZbFkbA1gFivPMq
s7wCeq0JulfRvhIwHqvkn6jVDZOQU6Yo+E88AYDCub4Nq6bdPGsQxfrQgZqQAxh0
1bA9Pm1l6DnlocZp3Cp1DY32SBX4q9D2gJK+s6ztwJpZDRJ+7jp+M+5wKQu9Rkoc
dyMD01CvuQtuY3lIs8YXaT5pqXd0CNFbgVI9YSQ0GVfQW2aGLzLlfqZRhgM39F4R
EHoe+z7dhhLtXEVquePcEy4pNuXMA/uoUr+se5T5QSqRImgcxLWPojYnTef1GdfX
yDK849O0Hun5sDUqIwCqM2Gc71nBjOQOCQZhtjIoLrfGhyCeJwA5zDInWFIUZQTm
qh8dXSFDLE9G28j1y5AmrMGP8TPeXW1LtJHK/78VXfMR36xjWUZ6xs+ktdozgZce
Hwb+XsVSWTodBDtOVjwQj6B95e+Pfz4Qvk4hRRJBBosq5BYqJXGvDKmTKYfCLhUy
Xghp00HQ1qg3sdGk2IB1kxJMg0/8oH+unjY2l5Mc2T2f7IULO2+Eg8eJ7Tcu/JfZ
StEl4uEBr23AICvL+HWegUISFzRz1mRnv5e1agMYHmZbIRf/c47mnTy2B3Blijh9
vq+kGUdZWB90G3hKSfvCnRwUHoKQl4W2LIoZJsNq2u72XjwvKehUphVxsv666pIi
SL5LkSvFZRoDHVsekeG6qaTKtji26jy5kARg/yZhG9k5Agk/khaGWdDx8Ag5GSft
GFIfumo22NG3yNP+L/oEacbrzC1m9iHWAVpcgqtbFun9kdYLZ2TrGul82DF/oTIN
0vuwqIkrZKKNWlFu9ys3i0dps3ULYo2ze5+pm+eiGflnw1sjp5GQnmyR1I7mOkac
+4qNd7gnGMTMN4nSFeH0gVMonJbZUy86ebYgHRYa7OlXX9awv+U2DwPMREMMQw97
v82pu8Bkf0p3u9N+jj6bAQexlUMzQEIbCanZoEkiEh0CaBGXCorLY2Kpd4R1lHph
y9UCpXAOiq6E7dkR+MXwwKwkUa5OpIAZ1Ztk7djjhs8MsZfbPfxfM5ZhmLTDxIgA
iKn/BQaJN5AEG+GJEFaiysAU3b4z+6hgwciDl25ffQYl+ZuF/Gs8zq0f9KkvrkIN
Eu3BZhVXU5/BVcIBy/RmCJ5OQtJxb5dblrwJRB4h0vCtkx8qpwiUmAqff5ztkqnQ
FMifGJSWPUkcBaVSgucVA2UMMoFwIlYYyQzxx/WcFR7IQl9e7Tf5W7wzCpf80PMZ
B4Tl8vgHaBuzizkPO1vXNCrkfQUyTDqBiC46HE5mlR++NLmSa5kRXRdoOvum4LEI
QISdWUstEfKrWt1OTcHB3fj6AwV3FkC9WnmcNw50BynrLi+5zZKp9bSwK9pPrfa9
SpA/u6MDUMywVgbwfcixCg2lAw0ptW+zS/DaX6zYLy5l+ouOmQCODqXcp34YNXuK
srfC9kqpvAK2tDx2sZSNd8HL4g3CYKZFnTf3IqnwOyNQ7nYCYDp7OB9FPiQAFgig
xRzy3F+61sjRdLSni9tMMqZy4eVGWARglbLixiMWj3bwJfgD/8yx8erM5IiNfvkD
QotRjPZOa+xtOF5V8mxsYKll7f+y4QtPxI3d5uyNGvF9FbROKOdQOCZG0fwzkkiz
Y+x542gguONKamvdAYYaEFu4Zkg1knils5Q1io1HeofFI3KTDRrpBf4xsiVRAapL
IZxFOzhcFOQXdRm5VS1KrKpXQTGwtD9bu0xr7vhCL4QmRE0DDTFMSIMvq2T3qQ+A
rXCwgl0i9vCXOlQ6I0a59Mz+9PQrFhXSRZc5JezXHHTWtwGBoeHYDPDLWOesLNju
clEw8ARf0v/sHrjWhvGKIRPvBDiDjRjIaL1L88iEkwVCkytbS8TN2TpCeImnhO+S
O0YC3GdIiEoT60xiqcOhQ/PwGf8cC8woktKbrCJGXn4lUZK7g40zvvN20Q3kVzRj
TtpPSBzM84lIxZBoM0JH1uK9N3wedYYwSbsHUaRzXpmKvvTLu+OE35R8tsE9T/Ec
/GPrGoUd6PSXZJu2vlozKRT+82bpMJoKitQZIIlns+HclmsBojQYzRJ6YP7p3L8Q
rsg+f0BPyabmDJ1wFIJWA82hJBknx5ILC/fLtVKG4A8IMawn/peRPYNyfslwHiBj
HnhwSpYIsbTnI3f15+qVAb7RgffbnSTpoKFinfJX4BRvQhBMQ4y905pJ8vFJYm2W
2b4vkK8gAzMmZlaI8fQfBUfuvSAymSl2ylTr+z6o5SDihrZ18La5QappHXHHfdke
tLpE4+PJ2LJPbQVsJIrM1koYfOgVjLrw1IYYrbQ9iMBbflgKXy4jKREYd0Y7k8dS
nL7AKKjpc/6U4SZ7VpWqQeTZZon2JvqahVVLOFnOhkoQ76Ro8fjnBtrbF8nMFkaX
yYp0fBfzf+5dUx2TPY8rlE5fR7GaEg6+sr2Yhq+b0WUtOAliCGje2NSIu2MdUlqj
kw/LGRgM09kOpDO6Vjpg80JDrtWXXoyG5jPcKaGJpuLQmvr/O1o8+OXX9wIa8tsZ
1Sh9E0mhSyJmHaoR/2oEn1tVNt2EbnwRCBzg9jpV9UyQRYK4l6hOKgmBJ3nPXRgV
n9z+OBS8eadsH2qJ+kkWrWu0aH2hP2FPQKhWaMtsTZRnlQfY0iF6WlloupQ9CDc0
O+JW5b+p+tssG9iL1kwKLJbSGlxsf0yWIeGizi3PirGxcn0K/tPIDT/2TK9LbThd
CqX9r+Sd9Ka47AnyWa7kga/cOS71QZSXmpiKYCHvk5E5CGqcI6rS4DrHgDL0kCTm
rynsUkly+UWAlVPao+DJjFlLmNlcDzSf35tNTt2LUbzm9HDWrlYXzi/TdEC0O/UW
h63W3fplJyqRtAiatM1RSI/atMe8LBB6drVajw8FVvbwCDU8rmt5R6cuxcOJzI0i
UVpmJdzCqq4CGKVC8VMdizuo1cu2OqvfzikEL/GTEKb4seWR1HHGHjYDM7ljeA/c
XMf4/wR8vkrWx3qDb+2qu5ctA96+n3nnlpGQmTP5WSNFGH+flKhNu3WfGGaJE9x4
W9xyGCDtOZcAFIfQW/pu3734w9A9jTkh4G84xubmE7HYmxGnE8fnFBuoctIvxbw4
isxGPnktiVODE/XUG3LAt8nqdhdAkPOVL6gfUT6nJyiChFd6htEiACBPOJY2njYF
gYqts75kfF5jtzFWZg63+0hhE43kDQY1YioM0AhR0Mf/YwmAxHBJcw7Tf7U1o7zr
a3Gz9iggkkGNT66nJEsS0Fey/bJRRfBR5ny8/PMp0qJNB0B7KGh8TRHoAjntNkpq
9NFUT1+OH7VIM5p0HQm+pL2rzJ0ZM/owoAbgFjMrMNnQ3Zpgt8dshZxIhGxF57B6
jk6zkHIlKmBjLwFtTrTr782mSpqR4TDwSeE3q5sbJbD7dCfkXyBxmbODSJkHe2JJ
OlUT0VtNSwAW5Wxd7P38tvRpr2WFSp09F/7WEv1VuxTnYO85goq2pxTEs7zWNIPY
WmgRvtQsxScRxYzTGsYX/SVWxOj+h21wK12mHwwUOS2ZtNEFiRh4rQct860DzPem
JUngYqor2g49Xj/ADZSv7Uz5J39eBAQNdq3A5ipGfrOFMSpmYnExWUW0rAUOeYYR
T3Y8qKxoAfy2Af96uJDrHk/9xvp6dp9vF6bcU/zUtuAX3JxQwA6scM5hkBViv+66
RHwZ+29c9AHWnFMuVmep+xZo09jm9CQkLOJzFMgJeJoeukcSkhOMCWNofgXZpRTy
R1rchfR00oSf5femMN5rrdYbUkJm6KV5T1+GAWz5CUOz57K0g1qN84bJT+0GdfDV
yI2fB2/408ML+KUUNDW/OL8N/ZWjwMtMdARs7wKKOozBM0NrIgbNc9XR7dcpH8Hc
9MxIJPn4uBwHh2O9zbBjRDyMbO9GuUZ7ku6d9Pc4S5lumK7O6Lz9Sh0OHsS5NHmR
fmDQ1DyHzM4G2f7rTcdJwqDEOCGAOCHKPEvlKdYWeaUyw5KFYFztZ8Whc9rT1gn2
olhprzrf6kf7fXXGVRc1ynFymVmHKuiliPNTC56SS4Lx3kz9hyPkr32mOn8yT7Cd
i96mGi1oeYA9ejXVM0odIJcVlsq+q2p88wDcFkNtiZ1AlobecbLO6jTRWbgPj+ul
0gTopFCdmUe8kyvKabMaHDVjldA5G65lktYPL8uodgRBkYzooiuo4ymnu3SJLf+F
B5bofjHhJ1DeDZdS9dnrukmAH42ggUEWahvX5BMwqoBBJY2AepnNG3ZzwtBl0A94
KL6/1V6GbMTpZ3c1nccF/Jf/cDpTq/FP07nLSItkzF+ID1Ra/Al07w3ScbZY7ikF
cbqpTi4rgxfUs5b6hTu5Awus9SDGaZ6K8So2SB4V3BcO2smOx+qJcAxW29DUeM/H
k0S/9ZynnYzttQnqSCFHp/WR5OqgpCJdUl8idyKvNmu9Q3oBh9QF3ycoxi0Fz+5g
/AiV2MpOTdbIjewMB0Om0k1lZe0qKIQo7UVrPbBe9iVr9yqlbYTpYpk72HOj/TpA
G/q8JU+AEgFIUanEFjXCyucq3diEuVNy4BDyCbdOFz73r5c3Ko/w4+mbFnDbsLW0
Cu427ISFrOLPuDBDnU4GsdwPRwrBJAcXA/VRNxnFGQ8W+PUnKPwKnzslUhLO45QI
U9GKoq8huy+DMYRPYa5SOG3PxY9tfOfrh4xvCknNpGPBAVYJzGuR/DIdqORKV7OX
WV4HoV4dIrzKiUuIu9TtHUqPwYXrnK9i35/HakrrwNRIFRtB5D/SQfayWokVDX5z
wa5YtyYiaypqPwVgjnU41G4R+x6RiRjYrHGQceCnh2b3CpFh4QZI/3G2RA3B93Dk
9vfR53lpVrOl/C3Rs72WFRn0WvLoavLgEWZbjPb/bEmF2l5UkrYXQ84hLp8imLUi
gzHQpptnVVhN8tdJawmxfpTTSHdFo2YIJt4/gF6FLhMXH1SNqZuLm3x+I0VzZvjk
ofI4ZGhXHZlFaz+yfK6zYyUEhjB4RH6OhtMqy0VSztjVLumxzVuqtdYeyTzq0R/Z
JpbwpnP9wdmsViy+gdw3ydw4awj/6gbTUnuY1AoQQpWn28tOdvCIr59DUD5NrWYy
P1yRYapbY17cSo2jRJYk2YQl5KSbV+HW1o4t++5KMtA44GfBz9PFYzboCoHNPnXM
QWIv6gyteIHVAw4Mz3Vxibi5VlwMiZcd0OrnF1XsFeNss+dPr511fQlfnhoeQ+fJ
rL00BAZ7s3ZSw9/fR2QnjpE/9PJolIfYC6O8CEmqPK/ysFCy96zQrEU1Q+/QcJ6r
15uU6c6F1yA9zYWN9hTQgOpF0w5PI2fSThruhEDYIkWc5k3ROaWRvQbRa3uJo0T8
JhaxrEtmwCdPBOfl3PuS176bov0Fhh0Yyc4lb/Dool7aBWF3dtbX4LHz7Eb1a8jk
C4GtJZVOoH+6sIS9NsVd3KTKq7g+zUjIII1qr97doACjOsqx0gCUPZK3lTMdSCHp
jsfFFu6v9OuY8oiB/txii3IllwNzGSvghQcAR5jaJswXlmYg7TbYdB58y/O06mXg
LIIDwqINZXPVd9N3s+kxGl6owH9nZ8whaXFvkUeprcaEViYDCvnozD5CejQrqADR
pt2fyU/RhEzuZ6uyygtIvgOQRrHC7BA7kgD1dmEi3qDEMZORCC/PGOQCs/jx+PYC
yPExUsxTXijsEaY9Yejc9XK7VIYBcTPmJEbW2KnX1MKQHlD/mANCK3uN6kdE66du
ZvcZkZJssRgnxdWpoUMKs3L8wCGmACEFL5cVnHLTd7MgYYQxUV+m4q1N5N5vZEaQ
AN4ndkwrt57FQDOTS9H3w+9tSf1eKTguVnkqbYxfN/3zWo7VdnL2UqkscEAjXeTw
25tn7sNfhHOByB31cBiT69TO7e43JpKhlzZVl4K1SBqRzpwcE74+iOckNXIYhRam
oH230wEhzo7peALEuIhRkG9mrzxLwdHdrnGWLSZIRON16MYDKIf5g3P2mEXYR1D7
EUvOfmhr4yBIUg9AjqI6hK9/VMDMrG768tl9WG3Rt1xI7ypfiQzXsU6MeSAiDomq
CbUe7kWlPR9LMPrziEZmGnD65XS4dv8zBPxD/L1f0Nb3LWwLWsCXG56LMDxX78lv
NuXbHE1cy71ER5CeGk2/ZHpyuDJdiIFv2SPSza0h6XK1G4d41YNUsjOEd4BbfFyd
5YBf2n29r1CBbZubRLMbhlyCkY+lOjFfZkPf9fWNybWjH3RGMWvt06bW4If0SUV4
dqliA9a3r+m8W8lBq+EWL2k6knzc4ucvpeJaL965v7K5fUwC+I+/22nWQVDRk/+E
fgv993RxCFIC+EqfuFGzYdN1lkvcca+SFZPzoG4t4d6BkXW/d41rvLBXN8oCv7QU
wPlpQCAU1/cgoPhAubAoLDOPwuRayYSZoFu+//C6TWqK7N/t1mspcw/GLib2OSak
IKvAbediujvHGAnRljfoONT0Se3hagzMXAQXJNI95jg92J90T2YhybwPBNcycMGa
+asuG77k5eJR+P8FRG/zV5pN9RnlLywR0QTXcZeL3hcjq7r7QMUhCGrTCfWa35TW
fj85vnUh72FlkIoM91f2rKhbrUNeF8HjJT76wd42fMOQ2XA6a+YMhKJJ/w38HCb2
8Rt+0nBLBctXIe3AoDJfdIaTZDJZubngQfyT4YhCVqYd4KIyWTZXoiXP9BHIEakS
/NwabJIRh5SSQ0gaj5/da5+e+/hevC7A/eWzS5cOZjuI4lZEHXvSf5MEvIRjBrQ/
ehslh8WTVmr3p7frxI77GSI+cMVQqpdIRmCCgAv/5MUeRNaUlJ0cGVMDanESC6zU
CoS/MmGTYedlfEubQz0bA5zk0qeDOecQFSe9Er4GR8H9oRrmS7lKQ9vymtTx+pPj
6W2b+40ZNwEsQyNDt+a9muyBpHd90LX+uNlnSpIpuvy/c8nFMAXFSXUiyxQtxdLI
XYyk8ifh/P1KHrqeJlc4gDzlMqI0v7pvNNO4fjdKg/W7Kwx8HIf78CbWmY03r389
ejwMSZ0Wx6Gaijy6Zq8yWJM1YX0QZBdNjQVrfSjZ51Cp5MDIwNsMTB+VgifSm5EI
dPVzP93iEKtYIZRqRPh54GQmwrcuyQD7D0YCUPys3tFckzvyUG0hCPJa6fVapI7s
ZbSlAxjAZ5+MA5ek55iZ+ToDsHozTx2UT2NvnkM1fXqGCk47cMtefYfsjHb+Fy5A
g+qAGccLh/W8Aw/yukKl3yh4ms3wyHUq3mJSuA/maOw4g5lg6ekw5BgXVSHR4MS6
X3iJalInXjfHQfZ3mQE3gOEGeinHO40XgUBSkzqBGLazrIT5lmAHm+2zouE1jwe/
GxYsCQjYCSgJqi8yHdPKXBg+617hqOeD5onalJKv7DbUEGkWaTyGjOr0HMJpj6ix
J+HwJoZWz7zQP6V0d6boYljxDaB1cPYdhjQfumLAbehizT36PtY2J6q5P5m9WeS+
T2nxPbtVcPqpQy/Haxfa6BPXZEPoUI/6xe8+tLYrMhn4btejSJEzr3hPJ4Y2YeJB
4GtBvGOPTxq6QfGGe4sWOTnxeAhyQt9p29TsrEDYRg0RjK6fTyuFDVSybEy0mOix
23jida1k5k7fk6ZkHbbak29++ohbyzGR+c8glwizOmGMDqQn3h6UnLlhLGz1pQ4Q
LpsYvfLuTQVREFFLn5h3wisTv5/Lm6qN4ycDEovbLZz36v8VOTfbbtH138a8oiQV
NjoTzNYDrWOH0rtQmMHDBSpXwX92i2VOJ8vfGNJzKPuI4deijCvwZzBc3JyOVQCY
zIfiJuMJCGDJwuTxzFhX6u5cOGWU8+Uc/pE7eAYWpJl2+ZBbN6ZAmC8Ccs+eC0jT
+rmUM4w92ChpWwRvj1bGtMZBLg/an6u3Ss1g9Q292LJA2mZPxAGBZiMBbpxNYUhc
yQVBtoW83wpSOFVEV8QDmCnwEMP1ZhzX17N1sEkzT6mA/SI3mP6/14vGBkVm8AbE
pSY0hWn4XJqSQjlP38T7zXMsuxFWdUttPv4JsiFVKXvZV4ARq6VSOf7n43q2oyeG
5ZGFcJxik3j4kzbcv2ZvM8YEO1NIsWvuRgBYmG0xnrZ6a9QG3rjoIo8qPv0Kh77o
TPIKTcZFX/Cx/vMvSYQ+PpYn5iPSIWTJ55k/eovo52nlQ6tKYdauVeEBua5nmjhF
VWpFeaBl2asg9Tw/HlBKkoDCwozZizO5YrfN15rYR89u7lvvDdHYvgwFjXUT2IHR
hmMCZIyy1F21sS4Mk6j3VIlNFLE0r0sykt4dY/RmqyQUvCONmhq8z6wlM218E47Q
lDcrCng22Ysn7ju068loeTCvVV1lwn4DyErITfRmDarYezTC+9BsK2FeZxEwBrh3
bY8k+mILkcjsDOYgmnyWqLcnwXDQp3vgWFOgLLsxrf2uab1iJsin/T9jYWaoOSWU
nSy9rxe9U+LMIBuCsKO9JK1uA52GrWdMqOuz1EySBSTaU94YWj6qCEictLHyyl90
TZKa/ZqzeiPKknz5yUoDcttRnGzZvO8dxJdprVtcQGX4fxoQFosCrJ4poSWv0Wy4
a2ov9pp4BUh85Aepjov926pkEuiyZwRL22adtQW7oAkwta5ErDQQHNasMKwSGqjN
AKhWEE/Na5KtJ7U/1aLSHApEydN/oaS9JZ4pMahgX3DRscQ7GuNQLrMKpFhWhd06
in62QKfy6o1EadFZzs3qXyArm1HloNxdKCwY0SM4es6iQ9I/c48nMyD57SGUjs7+
Ah/MDuY2WyIavjFCIGQobkk/F1z46gBNw7wLsWa9d4bBA+RjCp6ghK/NnZDEzzAB
O2OQo/eNBwMEUUpme9ejURCVqWLCqiDjCKBZSGufNypV4ZT8mWSVnP4d8vmIo+P7
BhTM7bPQ3t712SERvhxEZNUVrN2/HFuwXIZ5NIEAxFkrI7YsmzWqSaaoeqtRphdk
E9RIiejyZj9pczJpYMUaAWPlQFp/WcrQNqXLortDxLJHaNsaU8NPd2EduZPYBNYB
V4WakYWd+qlJTuJtKx2uUC/7AGYEXpvS/ZSJu+7vpjNonkuzHphtgyjXiMVE9QIe
S0OkC9+Rxc50eKKUOEBIp4A9ppENtpzSUdUhbn2T3H90J/+psMRYGpXBzJ8sUFll
8Sn3uzsqG+3yUmSjK5icq+lQMWHv4xJaRDeSPHmMNPSdPfrV+LerTL1rOOKHAWEb
nM5mn+NAr2nSAKCRac7pVzjwuvr8xvNNbYrl7jzWwP7Uekq34cqUcdHwLGRoNnmi
FyBikYpQmrda6UR9JFJnC7LiWR4qVMTX94KpxaDPwDI8yQQDB8SKeU2XemmP9DTD
/9lVG2OPD6nDWwetUCYTg/gZQcg9tB/rHHpeL/Y7467JZhzIsGeDXuVOssDzriiE
H5KEhkqyjyugpPaO3uMFkczRg/coBTWcP0ADR94V0S4J8w3N50fRuSMXFqa7xI74
qOt5JZgjyycqxBgRog/xRGfpCl957tqDgy/ofRY+cCKDylwsVanlaFcir82FY5Y2
1dW+4GDbU00Lrr4MMzfDhrjUw5H5yj54HOzn787GbKRXOJmibzU+Js/cP/RCsERH
rIWvfnZ+vPGwA4DDuO5HLeKIb+Pwc64RYbv7ThMabTfLui5mJHxlxB98YOZq8/ev
iPwOq8nDV5NZfccPU7dF39jDsq2IBedQDvd8bmuNZBEpAj1VUqjh1cEFtvdAvQh9
ysnGRZLCR9+XQcxeM7KFIfl4re0Jx/AopcX7MOspE5xpoU8FLNjIQFizUCmbccCA
ezXX4Nav4th21funVHjpoH9SEDfGtQZBmZy3Too7mn1Zl0+TOIRzesqTVpI6dfDb
yUwd1ivFs8pvT8C146Z+cot9ddJ3im6j6BwtbEgXNwkZjrNg6ltDBfRVT4m+hK66
1MvKZQFb6s6AMDZ2q3947E6n7H6Agqrdpt6MuRkWamPIvHgJRf59EWAILjXLbbc+
SeOXGpTJj3TicggUf+vP4VioWht8xLhJvcyn1Agyu9JJHjV1p51+k/kH12PK4lXv
eO3Ua8YzzqDwPRCGlBWByE8ihPGmlz5Gur7+mW3lIzktD3lGZB+o0HAqDef8KQBa
77vfS81wIQKwwL4gGsacKkxqC/LidUZ4+woaWkBMVXHXYUVtd4MfCCX0eXdlaGkL
z/jWYMGB3Ut0W57Rsc6nMdYN2eDIkbMcPlCUgan6obAudjPK7kyLaL0zNTnndVzg
cjaUqNJbmgzmciVd0mozRQWc+76r1HAxlM2Jt5hzbiKOIKBtWKxd9V6F6igSVrnS
uyMQuUt+znSUcleD/lY4WlM8cRaiuy40eVSyrpq2E9EIaOeojpVHdF0uTm9vTLN4
J+EYuPBnwQvwRg0QMfpVfegsL2aavUqdxW9eDXOHus2BIZT2EJX37EoxMTECJvWq
+EkIvV/mnM4Z/K5LNojzy6bP/7faph9sRDGatojf0kIvnkA1FuMhpAeRUHXUA27Y
9bIoc77pr7KWDYSlCZNg9eImujbkNU7FWGJ2HqA6JzVvY/Lme4ws59QwlgdPoTPq
rmaGBYh71NwLwtvtT7eJ/byv3pUDtjhdGvOIjhHgI4jgqnJVOEOvM2bka676CqFi
PLEs6RxUsEDUQQg+vqhgJg9ccaSIqA7rhTEqPA1Xa6N7ezUZMzPS8EN7woWgBqgw
oUby14MTC2Uqd8uhNxaMPbgONufQFCMA9JYNnwB/8TFkVA8AHNUtlzWSBMcG0/89
kItPdKbmlmtHUqTFmX1+DDCAmYRGpa75jmPwuNiRiopG3zfm346W0ir4siFITdev
50s0006A2tL86Aqy8s0ypYSWHLSB93tB1xxpledibtWTkGtXJlU9L4oojdpQz9aN
QUb4x7YthQ3HTO2gjXyqjaaWHQwFGQBFAsdBRLXTPyXORR8TndzO1rc2yTmsarBs
MK4mywTCP+t1OADwGPX9QToTn4A7YdzIBEifT08ZlC8l1GwD4zlzVrwaYjPBtlyN
HEm89OXDtOOKBvcTo/y0jvT70yI3TdrFOiC0h2ZxyzK/xY/3osQszNBYBYG2AsrL
PytJQTnr4Ul6qLlv9RVTKrEGDjft86cDvAwtFMhyRlU1UMYAY9daCfjfhvIh0FT0
Ozc8A1qBava4XXnRRwMLdrw2Yv6J45DuJEQd8N0Typ2UCaIle53Dz9OEZ+GOrJBM
05t9T/p4zQ0YCs7LtKc2ywbtjeNXBkAMX7hDL3pKLyPQMfYXcBfOwu4KdhWL8vI/
Q6p2qjWUWsl1DFN2NT7lGKO/KMZEC95ywGyOquywbKTt96MgNfwOXXqGbLb0LY8j
9wplBwsijIxJU2pkfse+fNUeRFr0NnjFl2CdJEP8ZOBmw9jXLcwxQ50Mwn8dnwt6
AvnvTg6rXZDYb4WPa4lFu3rSCEgdjRGC6oBte7AthSMAyZvo5MsnIspuA3v65l6K
qt0KGYZRXXz+eNk70Q701PlnpK3ArVtUqQpQHBQoqU1wWgowcsl6mUZWUGGIbTy4
lOvB3lbGlBMQ8IpqxrGM4SAyYto9+OB/197FagbxaM9OsfQyQFncMmiajE0LmDi4
tODfl5YZU6skDa4WPX/6zE4PGkGrw7ccPtHjqk0j7pEQhp8j+nLj7WhBuSGPAE/V
gRGKQI5v28R5yjUmdq1Oe9RANi/S1k7YUDj7GbQA0636UxGOEtVkI2QGFJ8dAqc6
MuwG79mF4E9va7kaq//l1fFAKqmBJxepFz54fYWMZjoq5Uogpn3JTdX6MI0sPj+C
zpk4zldng3VzJBlAV8D04Lc4vXjW3wiU8xzYJ4Cjzl5vz01f8jhtYLYtaSJC/C84
EvOFxko6rPS97ZRcg7denSnpHOw2DDF9kMfLCKKbx3Gxb+xNKUTODioKm3butTUS
3l4CYibOijj9Oc3POPxMGZDVKqEN3CAhd1bw34zfBzL5JuTY//gPAvqUmv4zRt6x
LxCfpKDpm+U4ntC7t3r7j5K6nAkplPord/zQtFWXK90l9DOcpiCOKIhBmbUincrL
UipOEgrE5tsdWUnMeIVJyzYiT6aks2XZ18rhmPVby7lNZfJl4erHBOrDSt3S5001
MsTWzrr2xOVCrQIpUpWJCMKMfFmEUANw+9wms1OLP7KbgXkipft12N+rDlPB6GW4
tqPd01lbUOhl45KViFui+9Q93qvh3IQuy4QV1keWt3bVcyJNzf1SdykLW0xo38+E
EQrhfM/Q+AAfPa410Vly5OjQs+mt0qdRzW+0jm0jzZOpGYpBQrmq/UZUoA9OQje0
qplp4SLILWlQxaFoixcoXbJXhTnEPet5ccLL4cHnQIYqz6h3XCOO9MBRTt+aqV6K
HB/VjYrk//m/hbgnFq2tuKxpo4FJRQUnWkHftqU7z0FjY63X8bd6ebVWgzMJHAkl
fcORvqkzW38Gz9A5xJF0j9mH95ayD12naxfWzf1G8Nrk4M5E+zUL4ptpbafxbrIH
5K3FV82ytwotQFhjS3VBJSQ3/Lp2/QGGBj2qi6J8URKpejf0tqfbPn2SpA6/UWlZ
bnmiqab1vVyBTquz5n1o2A0clnCT/2P/RI9UloDssMurxPwx7ueviMxkW5Rwa8QK
0IFJh+fouQI0Hfvnsi68/H5lpM0OWoRHZBAGQ+wa7TwkNnZ306w/YekoEhoV2tya
hhfnd08ye8Hbl0KFMspSCjMWZEBgO3OpALFCja+iifuxjwxWGQ4K0eDF18lhOH6e
5tS3343i8pytlhcAUeTLkzh6iCBA82cIaZBHXwcYB8moa8on35bFe2IluKUKgMSF
Zk/IIncrDylTLnOPXa650FdQIIwmZYtHH1rSuMzrvk6cvELw5pWZDW276NARL4VD
IynSo4VSu4V68ZGEsdC9B5EliBUOn/rOj2Km5SqzRKACkT30Rh0wIJmLO6x1kpFn
SHtGRFSpeK+s/s51cxS9kgR5e2Eaqa+5dx3XEcsnK1sj2FNugkTI2OGotzn/cXLG
8EXos7FsT7RRcByvuN0wABWQzX1ETcOwoxwmDvEjHsMWxuVpV9S7EzdRyj9yB9yC
0vaL74YKnuwU92ld5XvrzFyMjyFCpWTiBFX1L78BtJxfqJ0Qjd81EL51oXY3LTBx
8yTx2nGOsGssnrJrJIzq4Ra5wtbH37HCEZ30eoN+l4N+7bTF3icK7PLSmCBH1zro
l+qhel/77rV4O5bEdtVGwSWHYj1BiD7srgkMjFXAiSYSTTwO6Jg4hi5BRGOeeUl3
U44Q0X3On0X2Cixywclwcy9ewJLhAJ/glQg9KzNbKg81VJCZ+ow1/yEpm+txQHFj
qVdP+lSOFg+pt/CiaWxUqDjXNOFpbSc1FMbz1y+LyouVYulGtSSvshJLLBbGJQfr
HWVhKRVLg0Te/mJ3MLOLVzNlqUz162pVaBxucfq48pn2BLEfI/Pk2wY9b8OAc65G
BR8Pda9IBPsh21K6WPWJOEwy0ckFF0rU+L/iS6YOJylTGv095d80CYGZbA7WzJu6
SZKhLqftuSsyMg51UeBkv0YDn7cPq8nQRZecUBG5dNI+fKfLrRRCYF+yF50yoqLh
BRqkX2ZJ2gi5I+bRj8nM/peGhIpUBZXIGcYJwKDU0WGd5SpvaXLC0LXFKKNZkXEg
f3LRd6AF7v+1EWf6TQ6fdLDcNyTXMxgHY8Stdjky98i4AL9lADx0i5aLr3BJG7ZQ
R7skV/C8eMwwTgpUBDjWsL0TytUpfYfAEFET8fKaGQy8tmv14JFtHFiv28+9OCKD
jIy9XDKh45ic22A4ERGWitlg4nkCkM1u3y1mPM5lIc8arNHDbWHDarP0ejybsDLH
swnXYJUJHcSqUo2IWHSF1I6AHb0El3OmW17H1ObJUHq2astXht8HFnuQNUYv5jNj
AhPgCYBNKm6O+ydiCE8mq5OhKwCY6B6SJ/J14KYwICLnsinsQ6Af3MiHw1ZidJPA
HMa90tUjkp4YiUFwjeH71L8ou3/Dcw2G5CAXktkkSfz8wgZmGMlkASYTdgBJ4aJw
fBzuQ8jOl6bu+3Lqx0y5OxEe1jl42UKIj/+5mJflLeOX6R/xLBVOs5KvjilTolAz
lGzJz1Kbd9UxC8yPDxLfPxjMWVGqWFaJPZcAePRaJH4Rb56eeQ03/THmrDnefJrU
xvvM2iGq0v9ESvqdlkweuiXf2xhl5i5VzTSGCo+JkfhjltqwaiO4ZfLAazVyU2kS
3ZpPUdTM2BYBmc9n26qAGmJ93WaA6CMYEJu2F6REWT67cg3obGdSNbWNFH7UTlW+
+Ad9jKjiBzvy234JZGZPdXD8vPFpRqf5iez5Dsb2iRYHbpXbqimm6SXH6UibOEEF
p6JEzObaPJqLuYJjJ4EKCFj8AP1/x9vTD+CrcCspXG6sQxodwwiLEzrItJ7GOuBV
RV3+/HcEdch53QU/VRLS+cP3VOyJLrfN+woi0/RJNTAPJ40xXdW4QSb9VuagFyGH
CI7oxkKtKyZ9p3YF2NZLegCgXKIcTOcy3inLN4+kvzcsWD3nD3c94RqcRqlCVxKd
tiSDOfvErxnxFSznq8gzxYp9TFiC/Uz3Sm5hRbaCviPUIvEZ4yYjnP2fwmL5KjBE
nCXxR0ZTP5G8AAz/9rgcGEzmLb8Xj6ZSw9GcZEen9LpHSV+a56jqnaW90KMg6CvZ
o9rUeUIoKN5EFSP0qju9UiTZEUWRIHGa1sLB+BCkcTxdGiGlMR6sh+qfpsF9hXFW
GphMmgPwCsGEugUwe+BToC317JDk1GxKy4K162+/RSt0yZ8XkEmuk4qbjvNpJOC3
UMJNFdnz+EvO8QV02f/oGJO1L6JSJLosrEWwKJrj83aAuk2nmYkqr+RxlTYSV4Xn
iWx2SsKIhXWykXKwdyX/BhB3y3wGfWrUDv+w2KhRWkBvuecZaexEkkvU5H8olcfB
W8WYw2WlHlEbItZmbVOD7bU7dxhiOsYwe7NK00U9GoaQP1RgWjvUvXUkg/SVvZbI
glXhohZBLBGwUGM7DDvWiagv1mUU3+H5T3hxl6bfGv1QXpd3eBcQz+bqEdV9hy+3
G+30hwq/mu9CVKdypalOnvxVibmC46QvC5I8FhgDaoUrCk3oEsNUucg30sSYjJVh
aWeZ0k1HImXUFW6yU5h/DXqoHTwfV3t/HgkVuFHrweyiyLiaiQa1EH5uqTX9yYBN
YMjddC3B6fjo4g721nm9Sq6RXiZbyJRtiJKQx3zJ7YoDJLCju06zKJmAeR8bHERZ
H9yOKA+hr3zfdBebCMU7YLk8AEswoSxHuThv43UWzFTnigIQTrl4G7RKNddLNp/w
Bx40VozxlLVPMbuml8c0OTFCrLuACKqH7FffxsuQhYqkwM/X5lu+6Ofa3EMsKsDv
JxJ4FzA/6xQle0rVNjTb/rH0MXpUdpyVo4RtvE6o01R75o9Llh4OBGATm5JW+3B9
sVVBwbR6PfCw3OHpQl8ppnfnlRKuOI7CL6FMOf711+CijHDy9ep4xR7DlggtCQEv
Vq0HBqvtcS2yFvEMABURdW89yhnCEpf9+BwjWfvfK5d0AlkxrPgiXAqpZopB/2yC
qIdwjiDoq8i35G3bqm6EYD6/nWXAjIuOg5MbjZp7JkgFYKOTHBof5px65c2pGACX
eaYMOs1C6Dc9ACqzCl91BZ170t9gOc5VYsUJcBpmDheeDp4wvj2kNjRJRIeKO3KF
ZhV/e7SKmD5taFSEcehxTkBzm/uJbEptYXhDMLsorCIVxlpFYeJGy+Xb7YV7NS2D
GNXQv2ChLKWa0P429EWV3p0VcjmFelDSvMu+AUVO1ACcWXTe6gwaRxEeWKl5QoIG
zcSmNYx+dUxDYloBrY9NCNaCx7sWLkxlaLupJEZqNbCBMSrXyP7412i+kUMyEpCq
LGspwFvi2CLmvhaBIrckdL2ppqyVj85GdFWFm377iWb/MMCV4nIO2JsxZe3pwwXc
D857tREvVRqxXEcfHTY99jVetEEqjXamrgugBOUoBZbEAC9Pl+m2HuyM1m/NZ5IF
wZzQfqmqYVux4SbKoDuDS3/CRWKdX+kbBMKBD+pkCxsfXYj0rPKJ+h/ip1IdvjlN
lNzT1NuqaA65xUzRwn4PAn2Kd+PvtfgQ2rGeRLJLQZdMqy5TroV5rLQ6Cx3Nwbby
yL0zN5txDAWzEOFnAbqqo9vN1phuRXXwHKo5t7rXz93argRVLDF73rK8RWEhazoC
LvCJUsSD1pbXD35SN2BjWez76b4KsJnWLHLouUYTXqIboVIKEggK54yRUWz2hr7T
PACk/OFpSp8MTrqKeqtQfN65O/pOcxm9DypY31K7RGbpckgIxkDpTWGpm9Aafht9
nFjymayegL26tQ9DTmbZM5nWI1geP/zDoPx79wamy0YtdFwf7y9ZydmDZPuQoIQF
EjrhcYq6Nx7lX/r1hlE06OOtf54hJyAk5mJpq2yPAMZtbOH0Dz8Fpi+q3VRwAzB7
eA0Mr8ZKukRl5rWRsU166arPc6QZvuN/lWsxHlRTMmSgnRhdwi5wDkUcGDMpIg5/
liAd8ppEHRl4MN4I6e+5xr/TUQoW1sNxZOCScwTQTxpP0qdgxKRZbZ22HgXRbizn
uW/eqkyzbzmsBYJLSM/ETGVmPFXJMo43YW4a8KCkvITc4XWob1YKq77KgEM1KeGO
cafeH4xjV3YLEsEOf2Zv8OBTkOFCY13AqL/z8wAd8q3EwzHytAzoaW2soqx2R8eP
na1piRcerStEHnwO5WwXP5xG18ZXqLXsM2AhhPtwAplrlipdjDL3xHj/ulcYgvpM
+JRLnH2J4nk/rkJHZfEDj4jsirLgLri1kW/B1H2zvyqw53DvS3vPdQKHkBxJjTp3
ZMQOt5lKJkf29wsx3v3b9+cbqTGz3Ulm1g+C9G9DlW254sfYa1Ko9UUjRKnaLMsJ
mXq8+8RCIa/nmhMARmkyX/CWw/h5Md93Sat31l+jG1gAOzKSxvb4TuZ6ZWQRq4Dv
ACyNczRXYGfwO5bIC+sSOrnxdcm3W39zSglM9sk5PR2ghp0VRmj+afi00Dng7qYv
rt6qiERDNG1uwf8ddvGXifFCLu2yVYHvLkc81OmLyWOxlDNs/jsrIDfJWXU8NF0i
UGkTagbMUeAxqvgqGudximZcjnVbp9Ds+jV7h1cCdL72vniDOiuHiwfa5zNUmNJ9
rJlotBXet86/RkIwrsF+v8FxT4bhWJcpxhBwwN0X5z9iuO30BJ4cMP+m9MZqsF7p
lm16nBjc6cXhissSKqlCn/xI/RCDGv1cpO68GIO0yUtdsNcPXU7J1J6Er5vMBaIN
CBSpGwQ1ztyMyB3Lzm5LQgPqAk/VdbwDGXAMTVq8Ti3ozPuMzSke775N4mw2LXUJ
WdndfZIQFpe/EiiZTonRveheBBSA3FH9hoXjiKEV8nNX9wi/YI+z/PK7QtdBHVCY
iWhR0Dx84CEcp6kFU+L7DAqMVHQDFEczGP+Eagc81ynJAldtW1M1r3J1hKlwOCV4
javZmEWmwKZoQb8HIHq+M4G2KT0eAwKJXUr9bZXkolN33XoxcUTSmWpifgTBnn1z
NtNqK9zYjyiGSPT/3yqxDUcVShxAWFD2IzKYCGSkzxBktvyp0767r8K+XrwzY4y7
DAcP3fwDEuE437Bl5kCXWAFDy33J3rEDBkSttsXA7TmQjJt+FuDUmBvY3qXKglEd
B3cyuhjIRaTs2z684ZBqj7vOG4eHfJmWAOhNGK/WZEG3yrO0V1D/mmKt4pkDJfMN
Whv/S8aLWqQm7auT1YVm8Gd3oj/BBZkfmi3pCYxTYE7R/D+aLOnsmcS6lnIBMPv6
z74JwCPH01Jdtpo3ub2sRrAMN9aWqJ+JhVeA5FSZKou+Gec/PYc69Ck0AeZcbWE5
8xVmUMQD0kqG3T47EWjaMRT9oGPbDG7ZGUgTmoPOP3IatoV0Jqqmp8LSc7VN7H0h
QXpDr1EBPMTyCQWuK3z+4XVW3ksZsjG0CnDK9Cwf2ahXAkGB/772VGZcY2kh6lea
pN+Z/jNyauTXqqq+jT6qJancV4yB05bTt3TNLaFXooydnC+V60WdnRCxF+gkPjVA
c86gPmzMJj8gSHlZNJ7mqwLgBVv9VP71E3cWhJGYRC5WNIy/JuT44ohhTNDlhXwU
VSmNRMTubcBHhe1w9aIt3tok75J1CbiJ8FWzjM3YRattucBLHpNHRXTAtAsXOSMc
8XzQbZ9HI6upujMfECkkBkbG1EdKjht1H14oC0GSSfHw4ZOUkkP15GAOcwLOEP1/
bO64uiGPeca6u2LWiK6NOFJNikms7ETAMhttwokAXVCYfgKhCq39qipOzBHLSoxo
mLJwuN2C/GOqGHiVTEegPgm4RjavkhnrcNhjm1Xh3OlsmENBTQZcQvtZo7h58gV/
bq5r8JbJYto6Wsab7X/tUYYH+zgErZmd1/W2kvF/4snxLiwn/XGjMop1BX6fK75b
MxLCwL8B4EQEnD+uazxXx0sRTIabfgSIaEpFz341ObMAPFK8xiujhRcasKTCp2c/
OJfwVZEo30sLjGjYn98j4z/j53LERGcKo8xu5n6ecy7BNRRGvc3Um3gf2lrrvtx2
0ykAslVzyt2TeYOCnzJ04KN5VfZUE0JkMQ1LyqaAiY+bB1NOttHBiRwHO9MQOovH
LBew6u1K/bf4dj+lI8h2aWooBi7RHCOTIvFuMJq4VfNBQVCcWc6Y2GVIGET1Ht5L
tZ/6r3r57mcj809SzRiNTBnRU/BA8QLw1dommVcMi+EipRVv4Mu5nhKZKZa+MTCz
kpMCWQNZAI6ajMdGYaGfyJ+8YLBGo5xa8uz2s8G8qe/qSz4qVixzE3tBU9vupekJ
5T86SueqvLoWGLTGxAlwcqWiHh5OjkiiCHWxf4TJzZmBfPOLSHxCjqzROiL7Y0Kg
RPMQo0PuV0oEc45kiO4wZQOfktwBmW/S01nV73xrjBnMiO3HXHsstvcVfPAxrpNm
E4wO+zpue62dhfuuK+NV8ExzHnM2cAXz5qOTWFqqiKWgL3UWm8O2UpzWs2cCarWZ
s4OrTmjXyijvB1tJJWr47YKcjgLir60+dtg3RC9DOdEGuolKvNSmGGSiXm8zac1Q
VmjupFTAeM5pQnhJISMNND1KRTQ5fwHmVwWwCTxt+Tze9hXhooeValEnZcKiwcr1
eenn3zLNcghMKVIu1lShXHZbKHPHCmyG7+K55PoA6PmFOoIg+jYgctqeAlb7qJmf
w1DWF8w2rYXLXP8Q/IMoJHAbh31qe/rH0N1SQPTNZZCJCvKadUj3aqWU1KR1NLxI
B9a+6n4m7mcOVtW/c8jqgjEeaRQD3wIRyEqU7SMVmGNb8Jw11+GUdYqgmXrvM11q
7XbqJwvgyQ/c8vnp9YTNWG2y1fFxWIyfPXpevzVPqmzQGrS3xG4hO8NZTx2q7Mha
iKxoaxKV8ehAfnewgos0+KrKB++wqXXg1drHAqUMeRttcYsUT0ZGeY7Lpdqzk0BB
2PiZFrk3PlyjqaJpFUTe3fpa8/3/qaEWKbNIMVt0Qc4o3siJzIdfbkgjVkfQEADd
HR3K7P43rjQ/c+AKHLpxjzNfjma8EYyqyC4bzECSyj8AM36xmfOZh4o+lQ6RUJOL
KAa0uZ5+3FBpY2BWYkEEH1YXfGeb6qwse1DQJvu9H3XJ7/IiInd6Nxc2sUlygRYN
XgPU2BzUjYWbITymft2vGvpf7Qq6NfkK8n5EbD6iDUR6/SbN+goYXvPtH77q86Yh
f7rHQndbFJ6u7hnYDNehTgxO7GpN05AE+yHpVQgNGBjAoUDlglv9BsHpUoRAm/Wz
9uYRZW9LB3hKVbMGAd7cixJgm7uTY3G2MTO0czhihUTbjDzoASDWaL7cidT7EcnR
eEkv5rX/0RwiV7QX0bEkO2UltU09aXuxxPGJWoI5jNS0qE5yRevAxnL6614r8Dv5
Hk6LAdehiIRkk03tWf7U3e3dIq/CBXtOAHUJXfqS8FSMVdcYJ+2SmVmTduSDGfJ0
fJhQ8aPIwNJD/vGUC8BFFuDn/5dv1KcnSSV1Dc/e3wfr6JEao1jHRiO69BsWbPms
BaL4l7GdcPWik8uRxn6Pck1wlikgqnXgE17FoTwSVL67/UhAa7abOrsstzlb5en4
ILU6tYgLhx3HRqaYv+/QltZiDo9+fn34Kwjmw69GNwNrXRyljSS4ci+3JOZsFBZe
SMq+2Mnmto+brU7mDogz2v5T0nh1cnOPJiA5Eg6dt0ET4vXZowaO7qFbM4AbDHAg
3t+YcPvzxwfWvqyROijQ3ISQ8rVD9EbfFQdPfD5FD2CX/yU6FD/YkgGEniiKOb3i
YGbaukE2MfZuzXi9eSPOqqI1dwiDcWvQd9j5nYgoMkMMolmEqVnm3qQrIwdCvzh9
Cy7lGDsmGBxIPkkA7qo4CnCYXyiqU7VwP0S0+4pfcJkz/yu9hp4q8bep67zBE+gG
iBDJ+0hV7RGgV0gah/1eIt4mjBOgKrVvJwnwo4uHdH73u0u/XIxZMsOjJcxbUBjx
tsXrYBg0QFWu5kvzCNAKZQab3PAL8nWwepGBz5pI2HnNi1nOCgsvDp/O9Ie8+UCI
xKoEDaDPk0mH5LPSsbmxTGzAXegRoeJyw7YeA6ynfDjEHwpM5X41K7W8agujhtq0
u3Mi4Nix+MhSQR57PAX/UVCDm6gCCLlXvhzxThkv6ERtApaQVeRWfpw2QluhhLEh
60VmucE8Ph61uApOjg/rZKPeo/oit8s1cMU/k83PhhqwcUukKBQ7i0hicACBMKkS
VRVaHT47bhXR6MMgsFsz/GwEaD574nLUFWk9WR0JSXB6J/evMB/rUS7/8AwBaXV4
SMixOxL1OB91B8ygMeBs11HszvCkiVlYwDipueQ4tC72ajJODrCFXm7fZsvkZiII
Rruf0NsPntm4wwQcEzo/nsOgAOXSYGBs7bLWKQ2TrnSlhesqP3bWZ1exHms4qhHv
d83jD7GyU2QTYBdUnU97MGOsYbO6fcrGa9b1HscPUY9FFaNesirgH+ixA410Ik5K
RyE4UZ1kZgyvX3gO8IN2BkF9unQy8uBbjITYkEiqyVkEfJXxa5pfbdefhZmqJdH4
e4m2UCtF/R665SHulShLHp0iWOuxX0+I4DFmPOtLIHy+VWIoN8+xOK0fCH0rlqSZ
eLNrlwY9U+F4bLb3hmRGBTGEZaF+KnTss9CTtsIcAkHeU9A+9WLFsSp2chwT7s3r
a2grLcAsbVHX1pK1coejtykpRclK1q55r5rBmaKttrSs1i6iMcKmW2vneG9CFtpM
TmbJfUeo7zNOQZrI1lBRAOXDBOTGEwMqZQK/mhQdf4L/OeSZLoYs5UEN9J5qgaQs
T4s6Y9dJFzO5n+ChbWVW4B9ujrlIvpqUm9sfAttV0ECqqcXMPpLlhDQVP+5ajpy3
MeTUZJM7taaGxH1E+nLI0+Kj/35YFwjyX4wyyCkGH9f/7cJcJoFSO6yB2VvMMezo
7MYOSjss2NUKpWExBGsOYZ9Mahd0bc0ugroOn3l9PDZ/xCPOCxsOmLpOFIii8fhm
JXu7JR4+8IKpE11oC76PulfHWXTj1PGmy0Ui8v5f+EJdegox9baQE+dq0iCODTDg
Z1NBPnDpfew9y0xaxtcWpmGnekDgB404lr179fOCfV/Qlykt1hCHJCrjBM4y3AfT
/mIvW2+EJfW4YdjidzstIbHjR0jo1kS2ns+SYTihnsm/otIZEIleQEUdhPL4uDBA
TVbdg0EZKtC+wXvieE+seNZre8NV2hf3La+1s7n4nZMjmDWXRMztzJfDvnlJuiS5
SYfJO38qW87N2npT0Gqyb4Hg3hOq313g+xlfrxPStfvpuLDNF32dg+K9qKIZJJRy
OKRWXhAWwIU1qJmiEgV/iqtlQA7lrnjLYD5WwQ2K0Y55dCZceXoI/ve2qySuHaFI
b3Mlq0PZdVMdXTdsTlf2rM2CBandQIPH85OREIA7UWWkTrYYlwS2PcpeXu4qsDDX
Oxn+pA6+F5ZIxskRWWQAwtXYRfayYwlZfr344sAg64mbenHA+IKSXso23vyk1RWU
AJItyaoYGY03NWYns7yiiboTbXTz0FPvLviSiJDyVtgNrskXjz2t/2KDTx7yDjOw
fmo4hfQsudkkinYUlwWP+ToYT8SU4f0x/gV6fkI+w+ZoyHk2d6GgdEx3IcaCpATo
sOXIMVq4X7ihC4heRkOltO0dPHT4qGXN6VLn1RabhoAmvCxJDXmN6RZL9SHzIVbF
0hXuKI2b7N9MVRfjJ8eqmXPHp48NtDacY1S808KUdghURekauoI3aUP2+jH4oBKW
5TA4S+1f/stp60Q67q0IOYbAWGtcrHBYLGedWJrflrvVsQxbaeWvOvLprJPnMPwV
0cdLDUtMq2SOvxb0lqQC5+iBNJ2NFzu4fWCvhXuVtdA1w1zltFTsXXOrukRY1qhe
/JD8GfZpIicsHOEqX+T5vJNPco9+cDjEeM0vUeWBA5kxioBlvpDhTZl5tIjSfyvK
snjj1re232zz82SYHANXhVYi9wezwNSmiHULrhu/mBdTuANyOYqnemDm26LdjejO
D6L9DwLkK+m4c6euOVYGs31ssg+V1mXwNtvQUyKt4G1pJ21FGy/7csBaK/bLwPQK
K3hbxII3C2cyGls9qZWpTdjCPfUuC+P8w0/7gOHusCrQAYKcm2frl59W2gDLfz+p
ZDvRIagIrARHm82UmUKGGPQtCdgNpamYgMnEcQBkMxp1jSL/JkeRO5O/tyMkomuN
vCE4xhnOkm80hSfCEBzOBBI64DIlyM5fc5SyN4LdWWk0bLIBe8K/pMBbNWEJ/3Pr
9ChncW0z4L1byVO4GBhvQvAmPSU08QuSKKoARfDjvcLjdSTULMWmJIBAyIMYJjKB
Uiz5AXWqFBjLtbHe+rUqId3RNigC0Awo/eF/eLz8ERTCJhZ5gjRg+OG7wUcqPKnc
jEh9/WbwFc8yyhN/qzOq5zU4QXG6Yii9Z160XK+4p6GWIEbyLEMtfChXwegewo0V
R0WGohHtKFrqgdDX39faEasYAYKY9o8x4fq3QO1szS//f5hhtVbfyffVp099xijH
4kNH90zgOtTiDOhVI4LFiqW9FNWYoag9nVXgCU9yntkl63uL99Eu11dvJqu8M/lH
RZT0ujsCyRn7tqWvJDlpcO2EF7D+MmEczNN3MFWyKwJ9zWBpnRO6WQXMPNxVgJgs
hWNPKYNUPRdQWh3uA0Xxhkvj+ZPXtHzIowQ4k9IrQeL1ThYQcD/GxRys4/1cNId3
IlwT1dd/gEHUMzVcVv1enkx2QcmHiVNaH3RQLyRY845dUPT6IxBfVjJ2hDwwB3Fk
SWntuO0dTPh62gkpoKCW1n3pSP82HyIv34qYFsulFlRDgmshawfvgHVN0zDE6WCo
m2sXXVffSYGq1rUOqBm7stzymjj9om1kQqpSt6kbeuo2L29l4c5W+Mn0IY9bRycN
buAOayYmBatCmIkaYcBvB+3O+LJ7LISuZ1uiVGrsoBDELbr9ehn7P3WL5/lF7qFE
mNWWL5gTc0f55ZX8a8tuxWoX55wbqhujZ5HfVFDk2x7wIC70D3+EQs553eWYLOSl
izkFVYLlGY518WXNkdhgL3/yGuKlXPlPvIWed7m5pDISjyRFHbLhlmVU6vfwnegd
CEQH/q5dn8DTLQ/kJgvca/pgCYWnXZm2B7dKUL3H1JH6MsyHKrvliGV6qEEcXM5f
juwDvfAR53PRO3EPnpasdEH1Lvn0RLk3fdQI81f99S0oNouDrbOqS5rBqHf/wVHi
8IX9jNTorU/sPJob+fP3aDiRHIooKmr+oLAcKRV8rHXlzmldTgUbTc4pn+30Kxfs
WY6ZUapt/X7TQ0AjYddBmXRrLzawnIzFusc5Nv3r74LepX3yaGpAzomu30dEMQUh
BIqyTX0LLDDj/K5VZSVQJXdA/Yjz4Cb2Md0MNEShkIimYfPls7mvFqTZ83dPvP+C
Hf6wNgeDNso2R4OYqrT0KdMxWGnUY/F5rPSLzAlh/Mt09y/cSdOv2+ueciRvyVLU
On7FunfhVedIFePQTkb+l1j8xeWL0K81QQdApLfRyz9wXpV2GEHn0rwMM1Z64rX8
9/mKJKojaQosiOyHrmgwBHeLyQAnEDokwyzxjjGCQ1Mg7hQTSRx6nS7M5+ueOb8x
ipVvIB6mMlu4jmSsKCJHs3xp2t9tKTIstW6FaGKP+OxHKyjvCOAjMUsdN0b0+GrX
gI6QDeeEXxglNPTkVvwCsA1h3HSxhDt817KBrLMqGmci/fPHZV0FDrl2qs/h2uUk
+kSY3OeKuyyNti8IJhFHF6i7UjIz9Zo9AvRZvNYdX9d3Rw8pi+vJe+5CJxcDoUi3
IdTqSkv7x5ucQF9pTrmQBkYpjC2t3FMWWC9ZeCxdGE1GhrDR4uz3nkhDF8W4y34d
Rwva134HvUu1elc5XuRknpySoJtnTjOWlx1lwY3DMNYXpg1KtBV4qD5oovyUYlhL
3ruA0JQ6h3O2G3sIvpcoVlEdqB50rq0UmkHNVYiGaESQeLMHyzt5vYt/G0hxNH1/
y6SQGkuZkefaG1dIsrBA4SToZBB84pj1ajG94kIDZbt6gN6dGPiOwXqXyyx1Qaxa
GYmDv5B1IKQKGK9/Fql9S5D4IAYkLRgzC9P/CEFp4rnkbN1UrMvIRTGOZVbkRJNw
5cfb0umofiN6R+J+VTmrE/YFm+NLrlQzpaH63xxHahC2BHk9kuzM2DnBvNWWt128
Fq4uFFotASqh4qFhjjvNTnBXGFOKOD/QVE+QjQYgJqBO7+osFKZ71et8er5aWCfi
MxkpcsWGEzaj1mC68oFAPKc2oCLp0cVYuSqeOnGmZtOkxiYo8rUxgHgPhwkJE2wR
S9v5JVjksP3eWoM/asj8Xku9VCYW60pmbh3KIu2Ia5k+gS3TJneutbdKOQrKObE5
+SzKwl4Y+xxRJYhUze7LF6vBo48em+L4j+l71HTw93+bLWXKrd7BE+0dL1uqeqpT
JQHa8A1+jLEfW9Y6sCHfLGZnlt0NmpBL0EZh1Fb4eJ73gEzjdgbCx+WscKygt1Km
+aEL0C0R4wGPW6VMAO7E/tzrUlmAd/D2WQ18EQufg8sQ+/6dR8smTLe4N/djvRlG
XZ2y6+nniRjN+Qr/W1jz1oAb0fXAWNhOToypU0PqbhEcMC2jcXe8mErbEu27Ald5
HkpUtOZKqyIvNFeaciPvf8sou+5kBKS7YEbN3Q5uOUCSy9xsGlHliyezJ17Whvtu
0xgAzo1+u1rVPMHDF6UCYKlmUro8apW1oubF5myxkEYpSaOxKgWvBZl7X6e4rjRb
3IsMX+kukr0sC3uJwmuw8BgT/FEv6qy4RA5wh73JHfhAyNeB86wrZVWZqrDNvZYc
ADiRnlR801wTdZlwdzQ+DKD+qqm8RdCrrNxFq31KtPL0TyTHE7cu4z5uAv8gXxzw
DtO38Wn0MW/9E6+xrcZo1sddJTx3pSVerA4L/Ac2O+UDxLWa7M/pniykKD/db/CQ
VKqx5zQr9nOW6J4QX6SoldmZ3Zg3iLzVeB6Gvi5XHA/5WshYKBvUBQBoIeIKf2l8
Nh6RhP0FxJkJqn83sEH5ed4FBzXbQ3P5cNwEkdzxe7ZisCWDbDl64t2+ybMBtRw5
ehqiYyu1373Gng9AuA6oBaM29ktkboSKTjOfHoVQ2NvxynBuqslQC/FVr/5KdOno
yZOU5zjbb2Oq+mIvTDPcVbfbS/bY/bsX/KgpSA15mZ901+oogeDRsYcHhr6h6Z3U
VoqmJyDSYQNUyIunA21zzvbm//ofj7f5e2eqDpX7CZ1MRKvBIkO7mFfEF5qrOnNa
xBPFwGsDReRiYzFbOk2d7auIiU6EgdjgVgOtSwDP3JoJ24mWirq5PFyw4luamxMz
fwCXnYGY6CguCnZDaxtjzDsP4z+Ql8JAVqPmcIIq3DQscApr+eGa37IFkE6cBcXR
KVAhZrT/6QdAC6TPuXabp9AzyurEEA3WUMGB0EJe+AVlAJTegtwMcQ8iDEktZwd0
M10Bhw95lbakGEgtQ8+L4x/+519yLNjwc4rkq+EQ21ThPBWUFwwHhi0w5Bwt/My4
GPdKKS8WGiyRoCyQZjUL4Mo0XEyMR744aWPFB15EgKzjU6owVxADbIcIFAddHQ5l
8tr065McmaFxTxXXBf6GxNbgFpEONyiN2aJ1xpsGmKDXyvzon14TX1qL+PR4p/SE
YBHVb7B/euXuF0l/MRAeC1bTBazfVTEwQySrQfo9zMfKkm/lQJ6rFXqIqGK5R/S2
wF+O7AtpTS3NXWr6XBtz8Bp4VfN+Zy28NBgaWfbFRNbs3ZfEW4imLspEqzs0XAIT
10VUN06TsyderEWDVEPU2cskN0wz31B7Q+t2BAAMpD7DBJwuRdHuhiynZLmEoUwQ
kAyThUSqb6g3hH8QWLfMTdfEIoOwffvT2pidGhW/YbPlGZ4pA7Mn2cF21Q87XtaN
H8K2H3BIgfjVkkL7xWv2BevzD+jTpE8B8DPZBG8HqGOM1n19rbu/J2S4TiZuY4dq
sycTaLv4u8Af+EF8bL4zMROZvmbmT+bC2KoLu0/yLnzqiKYR6Qqr9Gso4oZLN5+c
VX5+4D5H7j0QNh3Ei36c8pkCiEkYUcf9R9pYNC0RHq5skT/L5W8YEoHykhQTBrIg
5uifVJs4tVqu5kVgo5qd3XOphBrn4lpmBhImcYY2au/RIl/BPZmt2D6j/7V5G3GD
s4qt9YCLrTraB20OnsaD7vLiv0jfa6iazzel/acqKShnXGZEOynLUvgDdhQuUGfA
Dldcy1UlApVd2UpjvpNQz0ZwvG6B/mvFl/4LOe8r1SChOdbXHoXGQSUrKVGTIm6q
mBkM69OsX6PDRvEOjKb9rqpQhknYsB5IynYc87BxqhcZY95/4qEDAOEhV44gtHuq
RUff3VEtaZETkG2iql3j5IR18wUmj2whROIy3yG748SYvWTHamQVmSbp2O/HtmT4
HH0wlhP6nY5adLnTWkPHETCQPe7oLS3OG1Msd5wG5JRmoBipZEYN+hShajhwwokm
48MCCLEVj2DIVlYgtORNbqJ4mtmb87r58gJXQugktlxXqePucgaJjs2b8WWMi333
n/11DlKDnx9B/NRy+lAbKm8GuUkJ8E6ScmVXO7RvZLVAekE/XSzv3LY/Cg3aZeV4
99O/8we82jiFmI0IAw/9AL9C4JIb7j2MOKY3bxjGToVxyENiOZoS3LOYjV00FLGC
7z32JUPtfKlIwztv+pHItqViluHTrFzCWIdLiQR9jJVMjQc1wEZRbvt8RWKaIXGO
YG31tD3bI658uANGaJOH/WTslAFBluGE1f1v9ZpDPEITxofgnwmcOBZSLxFdfJBa
182ajilHMxCNR5EF7XlRMt4c1Ad9S3bFwlh6nl9c+87rKotNKvkp242e4ewor3l0
bWAHZtSBN9fOa3wuVsWde5alFNzcKf1R1eb7s2Xr3hsWpYMFfebQ0mPCBjglmZ0y
YmUzMpGGoUhZfKVmeAkLrN+lwWw30ePW6xJ3YYHH8rFkxpOQLfHu7UGIwYay917W
Uw79d5j1uRrYbheD/4rEFUZT5wy7c0QFbCxZd6Bik+R3/n+HVUJ3qgeosKWFCb6C
ziDbDxIzb3y4rK9V6xnGMLxpbx+H+5w7HHYflcdh2pDkLwd5TBBsiT6Fli5CYz8K
5kipAOFbpjLyAFwS3ZHTGZ/NWyWP4I13OKzLhmWe0HNiaVOuKfuECOUYo4UHEQZb
lqEHrGwKXKWWmhe2UOMTKwXINkUTVoHfadNX2txL/I0ig/msCxLTIhZBuivHlxD7
dUkqDPHBqpdmW1pqZZ8I7qNXox4rj+N/+aL/xDLZAugCUvjuqCVJeVA4NmaVewso
ErGQ2edwPdU+9tcURDRHmIQoLAhKhO/+zS+FY+0uU7Cbb5H3JCM8x9BnbMXaP+a5
5UY3jL6VKR3nTrqU0WBVtbB8f8a/Hz+s40vBe7PhnR+JHrQHGTK06SwaeM8Eoo9l
1uWyMgfq/Nk1u/T+CqzKJQHZ2KgTdgjeYTlpDx+/3qlhfT6VoCaNcSU6ehNNyPzm
dcJ4ohFkZnSgewHX/Letx1fz2fnzWtGGOmFT/hsD4d59r5YG3rmptCAvm6tIb9f1
ya6+eGQJi4xhHlLGXlXWBRyDP9Y/U22ous0YZnsf/BAPqCQgzQnsxPpNUMEiAMJi
+ip5sodJEgZ9xnvrCyBIyEuCIlRroRzgTSUxXm4iLwF8kK/K+sNeibeXOJFyxdjI
8dpqs+NvhlTicQQ/6kFY2h5+vtjj1PE/0cwwc7/q7sxrgxGDrttZpm6iaE28XAVX
EQyxRq74cMrQKraEEJKAXXqlALBkTMDuarj8IkSlNh7uYIZA1nwyl5ZmmLoI0L3l
f3gUeyJxZh9bb1U+S5zJnRkquuJpIMbqdNxGbd7q0vIlcYzJYQcn1UptY07MrI1D
x8+SNF5k8Z49U1Q9SVFC0nNXJbIi4WNcbE6oJqjvhn/bflz2S4Fqfyoc0pMQ7qGh
Kb7GjqsaIGXjRgpnG58lVxG/zBX5vPxMNA2Lg4QQu/2iXhX5WObvmZnSGFquJdXm
e+MsvSX/CnOv28k42/aH7OomBAThMFE4ydJIMU+bX1mVu3QfVZ7fwHSjIfbv+Tzg
cQ99d76J+4dmeCHuQXiws2gDvJl3gGQcwwwEnto95W2JKvcvPi1OHTZ7QtNeLvek
qHclGqXKooO2JM996BpBZNwkac3XJIR00LrbRnsjzYL/jS2f3gkW+pXi2W0EOBkc
/lw+YgwZ+kV4PBDU6tdWZfuoO/n6fhE27L/2vMLvFCUEgoLIG23DQ37pRJ/1wElD
EykKAViG5jfYMLSLGyKUApEIpam3o+kTkQC8Ply46tNa0UwTpfY5dw73qKr0MevA
8bhDNPJ2vrXEKpJs7NqWapRb0z5HPE8+WbUyhSRKBISWb3MYYRrecYNu3kTeI0Yp
UmegaO7lpvMnt1n62Hl4oP0mf9o7zNmz6UNjJ7SGTKOEqy4sdRdb8cpFgc/ZffBi
6Qp3LIkSyM46tkHT47H8V35Ocb4He7/v9Wn/JCbjR16StolEI6IYdnEZmkNh/sYD
DPyPxNLtJ0NAC7oEJFpFYQIqsAkz8xaagapA5HjmoOAtog3CYp6Q412wshiLpPIX
AFzJGyXkVX4UeUYYETw6rnkU5bvQNameipnrr0YWxP9Roiqd3cJMTPbHRg3ZrMRF
6jHr4sZhfk+P/1+Tfm3SXAK6+JcecxpNkXw7+zTjucI9wgca1MFrhVU/uM0j5PU1
gn3qItArc0t8DnSGw0ghigWezgOfx+MAkAV0NrXuhgcWU0NTeQyEA0dF+RcWvmvJ
S/uLFk3076i83dZDqmJj14RoIBMVUbDBpjvL/cRJ78JFe7lWx6itPe89CzrZEs2t
kj/DIoCVCcns2f3wyp1yDGWoHkLsP3Lmmc63/NmuN6xqEEoJK6P7Ttg2L3CV5pr0
zb4AWoKrWyxmw9LW1Wg7axZm4GZcb00AHprffIqC7Xm+xlkcwWSC4R1dMVP9BHva
6iEPwp4qDNeVLNjsWC1qfdOQlX7Cxl2d+RGg6tafrnS6fGBqMnLHAWG6Eb4D91Et
ywpRpX9UbiSMXrmQRUR3Er3FE9aNPngXIgdb1Y+C6/YguxJDoxZ6jYjN5IDqwtLq
P0XmG7Hq19mRy7IqDEhfSyLuiPMvPH/0yRbAzYYTr5KL+v0XMm+bL7ePLQoTMFcv
uLeaYhj+kxsGZ7TQynPCdg9C3moaTGh9+xTbqbbEh19q2d2GlYcT8WLt30U43xby
3/89RBeNpDmIoWOIEg8RVEJMOw4AKchRoFllbqgLJ32dTeuX40H2nRPXDkhijv8a
pCear6iAc6afOzAhvkrTsVVJ0sG7nyS/t+3acJ6Zg8VcWwDSg470cmkDRluASUyj
NSdaenuZjNq1y/GKgREyRD3LrgR1Kne7JZ6yaBkOD/XwAsqzaqfWHUUOkHYUKqGY
sfCpJwlmrzbJffULPuTKRcmdVb7CmSMcdLn72ve5uKZoO5HkBqQuE11yg2uDw1e8
tq+bSvX81x6QSjNoZpWMnB86M6gTmMXU18by/U//BSJtK6VhxPPTLe5mnJZhHjWh
J5l1uEJwRfOvw8bgAuxUljT8Mw+1cQoHt0U0/SyweCSWdW+o1cGjMEySUHMjIi5+
JzGuxMZY+NowAQpL/FZu8Y5m7kWWC8LL8DXBB31S3tr4vaawGkEI9TvASuAyaSAJ
ZPQPyIFHHV2qPTH98TAw3DKmynO0ji8ET9e0fwdpOB/pSg1GsI0wCR1G+PEJ808E
BF5yjRL6oo57xdM3ldDunS76cCMOWE3AjCuGxkclapkRh+HzUtRYNjGDztsSbGuW
YsqTqlOG4Q6o9934bEoXJAOiEVFOcniuOspymVj5/CyAtKPZYhhPA4tlnsgNypGh
WZBymVVaVSO/BubarndXzNulrd0TZ+0RQp/as2nJNEr05pGtbdWMJp3j9zp2jC3z
LSpJOaE7NkvdH8a/ehN9kKJDTPD762Aq047nlBeIaxhLVwleWnlalUsOoLPRF1gW
Fd16eSIZ1EwDkpugslx9R1PD+Af/HCoXXhiDmtdkuvEx1l8UtPGeIANYJhKZlfNO
eHd0c1FnB+pwpHnFjLSU8sGqA4sLU05HAfRPLXA8RFUJAxgHfQruS9FSbb4XrFbt
97F6y0Ngik+eH7andWckqcpM4rrh54AfOHqC4NtpYJZlq8KpPkPPE19nmJ91MdCO
I2CPuGlCzR0K42Il3kAfW3Q839vcvVp8LiXiI6uyzIzeS/JinVVb1F78IXOv1Lmm
28KlO2RDh4NLTALFzptxVjJDnYy1oFG8GvrudU/hWjssEz4OJ+RmqZPPUjejdTOY
ZLrepca95z0t0Xl6A8f+IjsHn4RbYJTqFsm7eEDxJrGct64d1xcP+xbRWdwd77V/
SoKSau13nNkJtuqs9HJ4g3LyVZuuPlG1dZaiF3Xp19O3yvpvWQt/iewuezTUG+gd
Hgd/F0zCodBY1pZX4K3DHVwvvfyZe+dtXMElFfniJDnGwmvt6Hz15v0iQw68XPhp
j+JEw0K/NDVsviF8CnwBl5sFUAGWbKJSaWnuLU9FyJ/GpFWsqn7+bAluoYdCMvwx
wvkfzkj0d80DByrIPkPadbkhmusNBUPF4qHGkO941YpNuLXjcsBKKEiK3LuzrTnk
pxwSCRFcqY++KFMEJQwiw0a5Xk0Aip3PgXY7IpFIeHyg/hMCFYceQ+HC1dxF6Ane
uZe7Gr40TDwlqRgEUE/kfKxUKsOX9KYrEt8QbYuaVJh4qWQYVQuQ5ZcYK86GSCXZ
FgNpW9RxjrksFKHsohVQIuJn1CWv3kvRdRrexl+Hc2GDmKADlmK4HhDzU/rNeDv1
kFbZYYGksF/i97HsIz94L4/aW7eK5GkDvnumLreR1w4GRdX6gUWgWJ3MnqMQWJxc
b+FvxUDEZKj8p9lcDTAQn3yVL9vQD85sf8jTP68A4OzEFNHvvtLwWYDPPc2Y9tWM
66K+emqyfvL9/yoRrpf9ZVVXEF+855fWgbDIfV4SN0ITM/Zd4J+6Lo7O6of40xRW
DF7uGk4qRWSa57cs0WTyVKnXVnpNlogmizGmEhvkvG4Bq0bX7zruZCceyw2JhhRm
PEPJnOMgym7VvkQ5sR8cprUFYhIFdV9CR1bDdRGHs1NM0xPDVk6bKhPrvANb/TKm
H93KsrDUSJRA5dIvTP05TW6rvVNal6w3Se0nvgkWZU/jNrW7zrBtrFSDFhjlkVsr
r0ZdDAvDFg72hzaOyZ9QOMvrdwdEoUaom7HdCcFA8Xev04cowJOmiryQ4ZpGnzPp
diTQu5DSWxhtsvSkZHeSI6uIL9JrxGwpvw/cs/DrcI6U5IzBp4iMd84NX+bd6YpM
tCMSjczPO5MCNKqd/kolqym0M1e4p9Eqgzw++1wT9mOIjURUAUC3aveON3g5XNlH
cQH3E1fWnnRF4cDEqvsW+zt1139T+n2czlPTfC2CE0DzLfS067w/QPb5KeSVRaWL
c/qrY3f/aNyyEl17BMd/mb8mnHywv37tykbtEmniRlgoVHhjM4zdxGVQdSIrZ+PP
H1ZyM+SAPpgsf3wZXgGFcmnUDQ+KCiBxqFOMlQXldrSXpFpHf859bmiqu+X6eHHF
dd34XheeYahfNy/VDf21K3gXcWxPYxdsMMg1CCNlccrfgOju4sNWDD4LwMaFNwNW
Jjq0MW06OfM86O4U+0rhGh243FJEfFv4KOPCh9aOCTHm5sd/8oxychea2H5RDm/0
f7O/MmLDgtOmoj+L9Twqcy19t3Y5JsnGeHmko3vb3U8AZunoKh/qnUVgtoPNQ9n+
QMD5EHLxUk1MNik8Vs/+s9Mc4rbJ20mq+89oAAorLsheR7l/thQrUaZKHjUb4Qom
obgd7EhbP8zvtcOrPMFZ0fItkYFVK59FpbuXrSM+xOVGHBZctbBTXyP2TBLDOYls
SWwNUTgIWzHZfX2tbznXci4plx/m8ivn+fI9rxyQDwpqqtonfmuKsLi0m0k4Jq3Q
BEJm8nadLtrqERHZNEMaZIeLYx0qrrYSJw6V7z+1A1AaZIaNeRJrsZuwMKQ35AIZ
WZ8K6B2AiU4ED80qWnzk0z/29PL72tTPguAevil7fKhTFDfdx7BGy7VJFcayHFlf
9ar6FBZnOIe/cwD76ZG5WmM209GVkjiPBd0/rwhVXnZZKhLdyp5RcMVPTtR5gYaa
1W+v/4M9YdeCEbDjGr77iPNb++7c8XIKS8YPMULhxXhmm+qhoY63rJrZ769XqQAW
ecLrlpt44CEADMO+1gAK7PRxTBeyNO97E1h5pWM4sj0AHyxIpYDMWXGrW8JcXUk/
/oUeEj90biEdx6o5PtGeOyUY1fFBzpx6S1chwiB6fZ33KkaQTlsLGN4raD1y38dD
jdMRzoRW39eL+2sVwlh3vJi0+FFRbr2eBqsqTuWrLzWkfeY+Aaowu2Q9+LtSz77n
EeguTvoju6bD+KU2grU2RNLEgX4VEv7F3GjcLUXvoscIRc3FH06/n/hK3eXumujK
KYk6ChG6XqQf71VAI0cZYb7OizHJircLkgSLKFKAvzPZYvBF4OB0MedYVWq78t12
cZPar9KF11WWM8Bu5L0+ARWHj+6sZPk0+ndojh8NSaofemygaVuXgfvd8X0Q20gQ
qf6fh8q2v7SlNwjYGVgDzIoNdyxFd+HOnn3bZ2rPPpnuhVrf97E3KZW/s7l8jply
6ROz0bREqxp/+HjjL//7POa/dH+igcD7VRtb55WsS3DdmbQf3D0G+prGSIo5s+lv
P9Q6QMIqAjQAGkwscMtplvXknpqq+58/lH12HCb5gimrw7vV6nAXH6cdO1XEAh/v
vJGXHAVPFJ2YEEQg6oZiRywS1UJevoOZv2ChMhR4TmAn8n3J6VqaIwar4/jCfr0k
aN8bQgYw8i02zE6yySE/AfDsRndhlAcsPl/osQiHxGdsCH30Vin1jJN0bLuoZuG0
o6smK5EmQR6Wx6eAhKfO1U0Hz6KIRpVCg5twa3sj6MefgcpVjlzPjCDMknFiIGFy
ozs+9i5x8vmk6dQCU7X8hFwNZLSw4NLQScRKc+qwTESVrFOreDOMkzEbEnpW3f9d
HhDq0yYmllIHNMvtxndAJ5wwLPedVyp3JAissjAxoob/s72klZK95o0lvGSSvy+v
S+LP9X45iaPxEJCQtyv23PqFkwrBCIoE9dU0dSSB9aNAyNQuyO5N9UGa/AVgCfXv
fVnHzuyyVIZOoLX474wYvxRgXX0RT/SjnQ8F+j0vcTOhqixQJi/WqnC6CiTrylf2
pE0G7RFhsWijhnU4aNxi38resM1xP2piNGbE6fOre0waEH1RyJnp8+42mhf0eWeP
wjoznG0kqA8/Z5m31Nk4ZsA1ZodoKOc+QiLf1Nzyu72ImcqPuOtOsW5MdS3ATX5v
7H9ySmoBIHR9hP3VUehWqsqU38CAWJw11qSeG3EyK28ywzD7ZtNmydyFppykIlq1
SX/gTmPV3Yiki5hIFbhwKKK31lSlIcTBShkVvH4pKRNaFQSw6B58zFhN9mkPXAC1
kjDS9APtQsbBkKfl7A94eiyGQecj5rD5wfi/5VS5semB1HDUFVR9CRIY5CBfQczr
blHNxRsl+zeiknCg/45zXbJ27PKPN7jUspESKXzXqsZHgohTTb1eZmModk+EQpHP
AEfRLwwTnMVZuYcwBinef6LAJW4YUx9AIIPFyiB3zd21LIQEmL7pbGh3RMITxOC/
v090qhNOJxN6gDY3h+5pzqS4dPwHYvrvX9HhF+nmpY/BXQb9EfKr4S7Hh2AkqLD2
AdHCGJYOVykChk2yhqPAeP5pSr2hREuk93iYu30R0aKzdaAKlC+UNZDwQYSWOvi7
QizY/CgqwXcPr+udUyeRjrzW9GQqsn7v7TiMH5tGDFK6D4U/QK4VwlinlP0JM8w8
Ha+sYGs9aTA22LWSa42pn28zCz8qeO+YQe7cSpUfw5X1OxNeibYChzqdq84shuJO
TZYBY/XQ57Jp+hSXhelKy0kI9oTvDq0fgGh3IYzPR+ortf0FZL3OzWNq58v/6CmJ
hN9/YhTOGVMUtVjXwTWbrfUI7ikAZ/RSTpDJjZp8564KfjPdski8Vg3E+SEEGDm7
1s88ATsVxJu0YT7mBMTMWP+AugmpAJmirUk92UEizehJhD6NMNtm4KYBn9vcH3XK
dDCX6kS69/hTN2BKUQxXRBXSzmkreZRfcTD1CBHv2aKMA/Ja5fGh5RZOwZQYSfg1
yIKJ+3TMvdPaVZAGCXj33QOAwPjMWAd5ylmGUStLqcw5/tse2y4/UJJBq6gw5Tus
JsdAnsNGFAZmgVu4qHgOwmpp6ayyGvNwgEAFPG0Yv8kV4nQZPUDiY5XrZ+iK6c3G
KfkeKu1prF7iHXVtz0TV1oiJO1yWMrayJtKxCGBi4wa8kVnmQ99Hr2qBYhKH6B6M
w5mze5ockgTRqzYVlhVholPvJtBqZi4bf68dG+j7GCbWN0W8LbjpPBrOpuJtRl2L
0qeBrW5uFNzIlW/9SPefvXcJZAN8Zu9yXbpn4BaS+EpHG5V29W1Fc+zGJBT5vdX3
HmTmzwePBb259OlLaMD3Htz1VOYr9XfpWciWQl9qIxLq6VCfrzAuG4bIH7ug3Vah
c/5GApmmtiEbQzaYyDRhUL0K4Oioz2Kli551D3Ubw5kuVa/xdMGT0d77QF5+7uih
+RkzoGZOTe72//2OaFVes2dATShKk51d0j9Vp/kxwX4li9w2OhAdztJad37d3MRH
SnIEQevl9Hf4wmTgKDB5KpOK8wJzE3EzMITBYu8dKVX2XPKBGDgEA8KifO1ELgQg
U3PpJu8C+CdC4L2lDN08VlsLG+g5OvmiqL7k5sE7v3zmMLnVnf+DEfBZl/fTetKG
0y4ZQgcaPg+ddCcuJEggQXaFRLkLHxrIg5SGFxVdoYu1U7wO6M1k+zxAID8LDNwp
CK/PaZpwIzFl75xKTbdV0c8FttZd4zfIytYpk0y+6wbvYT1tNKnABsUpzn25YI9R
OpS81jqMeZbpaJiTR1U8dc9WngwTk4/XOh/Sl4c777QvzevDGugr9IXqtAbdByzL
FexejlJb8dvVnVkV1eqNK6crg70PxEzBQv4hHrrNRSJOfBpeFLVYqa02HfadhxkO
QQBlmofNXdEvGmL3HIGqxgVBKjFZbQCvl+GjjPtbum7XJ1zaT+35mTvoxo2ARyt9
m+7K5paOZxi8/DiDqGzEGVCmNL2Lueo9WFDVHI6dvUuKkDln1udegzdJulw7olls
CRZThe4NRawDnyncTtuF+M0opzgP+VrvxQjBeJ62Eeo1kTbG5AazKrcsYj1TSlEL
Gs7f8m3qFuYMAwfyV/W2pethz6CpWl6cqOvKWhodbwiviJT6laph4inH9UODZRPH
G9ZsfPhlORg5RUftAjLYfdVv5fqkyWW5OVFBQqL3qWoFsr5xG1mV8yNx7MXZi+PT
iRJ2AzMRpMZzgwvIF/zCk+91l4aBel7voJUxoNu3yTPZPpKkTv1FEK9FcoWhTOj0
whTu3LSmBAkBOdZbUP2mJQsl75tg4gFzubL8isHSwfvvyFWYVrUCp3mnw2+JE/7s
dlarpcvEVlsLtTRteq2BwNMpWtQmb9IBJdOqNcK0z4wsJkI2IKj8g2HMZePUE/x8
7x7LNQ4WhD0nYtcKEBNl1hKOVgYA2BzhHUAVNN3O/P0bMcjjlAyLFJOLsV9QNHBJ
I3nN3GM8npdEgWBnWxlKKeNzvBMcmbnUdWgC8lerwN3uVp+j64Iy2owC76Vee6fu
ap0K3h6apjArNNI8qCmzgLdHOUlr509X6qE3XZlX6/JoRTry7naRa+5BM13E8sh9
S2n/UnsLLn/jinV8uiLWzbR453nAYCl8gW5dzR9ROJMOzXWAToYfjcneb1CCcDOl
lMn4ilxHry7ZjGlHPA5y1K1iSu7d9NZwFlIhbb+egrQvAAbpAdjUDluzmMiNK8A2
VvqPbVatVMGvwNblTYJ+hfPVQBEPJZG6BN4YQ8Ev32m9Ohi+hfB1yKt5GTBzeD7k
7diNrGroZNZ6Vzw55CybjWpqm2WXcCKIjn80BPatKxpLIImxMNnGh3ZSeA48UPOY
EBrPTlgGWc+mpXc1ilQfLEjBo7w22L3IQ3NaZnE1x/lS9vJMPmOg4l0ab4GAMN1J
uLGjAhq+szgEOsBEP6Bq8DvtOWLq6fSQP6d1m8kxcUyP6HtrWajHcwUnhKi27otV
d8FLh+TjH7fHLutVgUJRv6Ojt8Hqru4qj+afrzxRePYiJvk/3CAyV6rmTg0QLOpY
pL6rhaQEKvxmSxlYIC/3TbodvGGY9ZcGQMdP2lg2eP/TdNgpIgGBYBq2Cf7+X3oM
K70cb0UePZeaI2sHt2fATCV5iL3d3BU3kZucBMf3t7+CgYpqL55UAIPshy8dhmGH
45kgtwlJLsgTBgW8j6oRRMVfWnNrPtK1Cao2tNnLYXpapZCtsaMxo8g3pz1pL0on
TDLRexQjyczu7K0+8A5bDL+XoQZUFUjQyWImH9LNtfsHbnG0p+Yqix45ykII2mrv
xcYd5M/21hzdTjXSiIcFuxpCV+VMZ2wsXGQXsJPxXV6nO8cFwUzHCn8Xx7Q8mS7a
wW1M8GEnlKKPvb2YFgzimmERGxfsq5XDQnxt+7iUKIc7BuJStfz5Bhjhh7oqLP8Y
2Ku/ke7WFxLT7SIl3BhSfR7Wj84Fjk/r0iVprnFxfZPaPMErp8PkBRQOEXhoMl9o
Blped5JRfEp9GEbU+c5nV1rnyZOZzXCtKxWFFLhNN+C8tPCFNlFL49LNp5za15j+
RSoKcsQJsFCFFI9TRfLneq9iR01MSPMFWE4wOrj3d4F9z3zQwfIZcUadhhjly2/m
jV/7H5vDCVvwxLq7hWBYKsWJLN2km90oGIPhmpsqI3txOJzCVmdBEXYmJZUs4mA6
rL82C5TyhXt0sDMMblnoCFAGYmWeX63UNty4mCtgFyUVWK8D4SOXP5YFs7ku1rcu
ADu1Vh107EjetG636UCc6i236O5f7an66+JijtkqLNr7PN1AUj45a2cezMYkGvBE
kKQFEOC/E715Eiy+EuZB7zIawQLTHPMNvicJof1azwec/lgxrIvocCY3lpChlO45
+nOZwuH3e2WWvPrXfBYUkVfRnbkxxGsHsbbPuZrdeQx2rT7hdVnJTVYkUUsuw+Lr
XZTqXTN3e+BuK5S7/8mJbCC1W8XX8TVg0U3YuGRdlxQ3YGsY7q9+yqcrbqHg4lhg
yLa0HMmi7QC3AHVFnwr1VcNtEhx+Ke2qLZFS95ds0XPo3Uwq4hU2znXQ0fDZLGNH
pj+DcX/nGZ10G/nqmOcHEqEdABvj68QNypsczfGOBDOCPGYDWhwFYNyVXqz8DYQn
8De+EXigeR+Nge/CL9Faib+NZEQwTpUP8fuAqxWwaIwuzZMRIw9icWvhtPUtSQdJ
UaqKDt6Q7UqionEG2QcB4MKza09ulQFDjBM0Yp78p7gdU33HIGKyPEmDTBCbGqlY
nH0nJjz8pWedRq8WYrUtbdq+e01QY8EH1A0onCQ8b0g9VzLGsxJqM40qNnTngKpi
6gEJIUf6XOqKTiEKgyXeBclnb7vIuZwhHyS+eKFWYZuyQxjqxT9ldxZQFXEQyEfK
TBjkAcaqrEQMUfAh76Dey/YHkrWZqbY4/Nn+JMlYVdFFddqJCtIKzne0FAhcpZ9Z
gYDXSg2cHf84F5uBsjDuUuy8kTxzucItA2xf6rWXgcWQV9xWco6FVgM5Ytuq+PTb
aYmBj389Mw9eObp9QwocEpxglJjEpBqJR2NKd6uFzyn/kRqrJ+1PP17ljYB6K6/o
GOZttaOm09kjvL/S3QQtP1M1ByKXgysaYZcXGS01dWb/Wh8LNUU9PuMyzDPr5Biy
KFier+9pSQSm7wknPeLo99oom5LUFXReFD5dn4b6bdbHO1vEmEdXX+G5T6QH7nPH
K8z++5/8ybDgXt6A3frJ8LEgJi2aizmQ35cUI1gSil9NzhHY50bOgMKKRguw4+Yt
kbRrOKCWFGf9ZSrpQpkLk0+mFlPQLpjEU1/tMUsQrEzFybBNoFX9R2Di2jNO3b3T
Bu4E/sX7ee9AO79ipg3WvZEXD83/ysbBdLxX9JX57kxJyWLnQMRNieku1zVjLxSd
qA0fL7REnyESbxGc31fXB6fkRxameMdQ/Py/4sDmVybJLb5xjXBlZYqiij1EWA92
XkUI44JJKmp7a1Cjw5J47+feQh4dNsSaoU545tp9r8SpeWZ7H98wFMcu8QD+G2wK
xDAcVTv0VgphjL3Y27/1UY1sDZuxjoAzVzz3SHgek6NmVNhUDXize2HLpa1mawJl
pPvbHZMOmlJT/gm1cX8MRQ+bdxdGeAhMnCXW3U0ZsrbRmQd2MUgP6X8WORUw99A7
m7iYVyQUzeLyMTxugmejHzjC4Qm+hQM/II2jYz9ja+g/iQdztDM0cl8W4Djit0Zb
9OGXfNCLDxNRVJm/BVzyQ8IFjQ7CpfLTWAI77GR16T//And5aL3hjr+twTMRVpjv
5QUujLfuyEqwYuqzo768c74OcH6yxmItGAL3PxFMh09Sv0kNL+lwj3HyDwnprjPt
PEUus5cW7i3558UD6LuU0P/jlqMyGa9MsrnO/Xuant6WLfskCRn4On0VqZvWAl0W
jzcPAxSPsCsRImojfeyQ2/9u8qXgkHwrdrp+CXjmCu9OFiYayRyaO0Gi3TWx40iC
EqUXI2SUgm+ZaLWHDbjBm/zywe9TP/PCI21+BCwwPunE2mExzKzad3F2bNYv7oTO
LWJjHp8kqPYuQZD+gNVMSN+bKdU0inrCuaj6sbu8VMTHlk2A5NxBEQb81knbDag2
1y0dGLG6HiRWGm/uWWCvuyKRAk0BeAAsX02vLjVIx1F6l13QjngDSYen6WcvJRFh
zUps/e6vP2rHIUrdzIgFwkFtDCkOFxosYU+OJjQeIT/vNTxvDPjZklOQaaQV5w0P
azBulE7yqUstaJTrycGS2rsb3emblBY0FipgWyxwMOlxggBF277E36q+H/vsKWEU
Mf1ouQBetplBmQCpNchNuSwgOO9bbflwvIHVLmQapKMDbh/F3xfa+PMQIr9mKAtY
v9eWEADFO/ylvWP/irIXQUIw9wlyO7v5bCRv1ox1WdmXFcbTzmooWseWl+Vh5gKi
Ly3bZ5xvJ83PxwAJrDxWyTcJoDBDMfRUw73yE6u+J1gUtPga8I4EWTfIA6DKGLk8
HG07eOXfpiMF06pVap78jt774OuCNGHtauLhixnxI9u6bL9UV2o5UMNzWhsl22FF
sG7SLwBSCWM3EalNnj/K30XMrt0NRULNTFGEErv8TS57DIwve+lK4STZG+/jDX6E
oeOrg5wwWhgRoax3ZID+r8+9ARaGWFWRehN5Ts/ArURB+rHISRYSunBwDFpDBO+H
dNaHf39JRlc/esrqrgvLcno4851l2uF/XN8X4w+MsC0F8sP+rmZLatzMmMJBTqj7
KngjicS5lT3Z2X0l9ZSj7raeCCkvOxFEmWlLPjZuE2OAxuchxoGXgMKPGZA6Y8VO
2pgdTF+hc2oMzqFvQ005s3dz1mRgOSiJwmuk9R5qZEIeClsCbrNjW3DKqJZKIhcR
AKqaOjmRhISN/wbsR8iONRTlAhfSQayjBWl8alqpDsigdIU7J01QUJtkW9ZxOzaZ
axBRTHjQRxNviOnBGR7uVWMVY03t1mEJIgzOgTsP+sRAlhB8hKbxpNiCVaJjZuU7
8ziqqglpKVcs6bNB/LNIASwCHnHyl9fW5hEK+QtITdJrfkoI9mABV9xkCO/xSssk
vFIZvYUluePVxSWJ7UyIO01/VZKFG9KUIAPRR/x3IgW35rzBKqS9GVoum8HTbPcn
PVYL2Da7prqrTc/NA8he9CpL90awXEyL0MUkiF3F9KNC1al6JO2Ab0IAY1RaD8p+
dR0PVUX9T7RXqEWfwf2UKJH0waTOsYLtXsusiaZjnVEUGNop4cgVkSuNErq/6FFl
zJAs00B8F6bEQWSr9YdMgQi86rJcgAXbWya9ArALq0nOFEz3r1LstyLRrnGIpWM/
8HkHs/wMaLBCARmf6EEZupzbh1Zpu50+lDgi2fSq1DDoinMNl4doU8wJ807wS/Wg
HPzh93CHy9xlSxVEXbz9nlH3O/JWxz4Trg2A/dDltda+2LNbzzqiKFyac2dE/DXe
YXRi9TKygQcljFIv6LoMsT7ZeMDg69IImzXkJKR+Qdw0b7tNPejV97Kj1UyHqzEG
gW1mMerOYIZdITUNrO078eBIySOUFE9CMXpG4CNyl7NZrQlX/Lx+cpbiwgaSPlhi
l0JFvWvhyK3/VuZzmlqdLSna3dUITjrWIdpCZH5VBa3YYGF4wWborlenjzRc+WvY
yAMmYE2coduUEN6DkAr7EKhUjAOI8fVhYJ3tdUB3cMJynO3YAieIj07La6l/gwe0
bbrnOjBDrsJ2whMU2H6n1FqtdryqlIVw4oz9tQUPsjwIV83vreGEFYgtuRVpekR1
GH7BOrbzaA4QDAfN+si0DhhcIQPms/1dtcS/dqo//6crvs6FwTvON8YP3CaVmJYe
i+poAkudYb8OO+1H6MZ6oNmHWxretTll3LkTIEFeLhAmKia1OrORlY50vuwuym1B
datnPP0a5+ASoPfb2MRiQt5A60EIWn8j+RlIHjHDjBTsqSnXd/bjOFu1R1DoTzCZ
Xx6rfdKzSk5RcBz/qu3xjRNCciQW2rHgnAcIuEZpS0fAr2gyQ2CmVXHV354Dvc4Y
GeUOb9HwV0CwuueLp4SXkfiojhCPF/q7fy0ziI8Xh91GF/uwGrrMLAkKfITP/qRU
ZwIEd1aNdVFYFEXRCu5KQm59xsKBorOqSaH84b3YywlJxmWRoTyw82v8OL0vzrWx
8uSw6A/tqcAvvvz/pG5eX9BffzQWjuPntBGpc1W4XZ9z1qd8nAIaMhOouHA7vopk
eF8ZDdhkIJEpnliz6/NMNfcUYKiZi935v6qxqBeg6lRAemaz58E1lS5V1ACtVd54
YYUc5z+VBODm69IJrpCJviFJjAM0JRoh96kQh753SCBqQ2itCqfgk0YQIJMuhozi
v//q6T87YMyF2zP1oAqmOfRqBh6vF8267vIetBATfzXlvBOFYvdipuKopFUdoAwC
oyib9T1QJWHTVbcUmxAc4kSbzZVrynJw3fWG5T2i/svigAFQU4nTP/efycfbJ2sH
rvi9noTLOXInZA33mUgsQbPbUuwww29QUh5LmloL2UhLFN3hyoYEV20Uf6rfjOzP
YQDLD7+np+jwb51ruXbo91PAtrVdpA1ofoPJjWYxA5QmH5j+rGn3P53hPqfn/XHx
KzPUq/FplueuvzGxcRnhR+SxSf7kYR/tR/wyJJGZ+EbtUQ4N2S1+8lwO8ZGD/kRe
CTAw65GPuroEBYV1EqWG+5JIDBcAh2hx8NQUn1URBFqSIpLRQjZLYa54ZxWsy5aQ
0hBYvangr9ZZJXtYSdHzmjUA90649EGCNofc+FqbZ9QxnSUo3YAAuc0Sa7FtuKHN
ZfnNMgO4u7E7c8yxrBDAS+rQFVPol6c/WJVJ+IcIOyzL104vwDMr5rwZ4tQovsnr
5rdeZTC89/hqBfB9Tfl2sxHDHWGKJbUerXV1BMSd+itbKobi8TaxYONVOLB+mbhP
QSwFmEjU1MG2RaCl+Ov9aVIHq2xrVr0W1MiXhkTAcuf3/phhpDDyd5SCMiwSG4li
CaNaqXdq38oWG90E0d/Qb+xbBvxd7wdJC/jSUKeKSlggYBHDIfSUm9OUfLe4oR9G
7yEBVydYcjXzBezkUj/b3QcqKRmwI0/seTldmnLyfTAmGbBBazA/Rx6EHqqv/9P3
GUYRxtu2ULmok984yalKn0PX2MmnaE0rupDyvBGp61XkQvCB3+LXSYyJjk8F3rg6
OezTvwdetDiu+yko7TmYJNaxzMjtmVCxPHWLL5UBZtnOgcRI2LJawTqNqlIBLk++
+Fg5SyDtVUVGbKCwgUGkQz+ujy4YSTooxTTMFL7kxRQEh3+Z0wdk5to/GEEUneR8
P5A3avri2ihlAcEHw5ef3TdOdSi+FhsNi/eJtw1bmJq1rTQTkfAxUqHdKR8mX5fv
BGXKybOUlu1P3NKzKgT6yypuaaAHVqPvxXqqVhXmB5cSd5TsMSpHVco4ey6VyO0S
EwhbwQMTAcri24+q0NJPgSl3NlGzQ/Z9i6WjlV+JqKewbDbaQIG3ebmRm5Hha6Y3
cSZh4S6hX2ttMhfLeMriOwiShukbRVySbp2XCvX6ArNR6nxa4ucBilyeov8vtVxl
tkIeDpvEBz/UTsbikAvOX33Nmkl/SYYaRZpFR6HtyUty2cn4nKnynfFS0VN4zf8B
lpm/niZGmLL6Iu+iT8+JzZ1V+x/M7tEPODk6kGaHqrRMR9L4s674lNABmsdZ1VWv
95IhTwXko8di8wOUhXNadHjYs+i53GK3FdT6kovN3Wx5uR5DBxdHO97410h10i2L
UjkHAqgwkukvcF4KOjbTHhI1Ibd3Z80dxLXuWfgJX8r051lnnpujpHaE5Ewlgz2a
UWA1jV7UIHu9EaVeOfEh2M4KBQM4pegSrIFyKQmbMQ3+gzjrZdTL7R7LiX7ifY+c
knc50wezMQDopff7lj5v8VI/t4Q+ngIP11EgcpdU+Ef5clHJxVKMQ56Gn67Mk/47
pgvrIENPq0xP4ZwAVdoQz/qqJqFf7NrHOCFgTie7d6gx01fN4YOfMtaAlzvvUdrU
cIiXeTUXD0QlI5GOwKqs5Z/p97a7aQtbCPJJ+vYpgTlj64vyyZ8tnVGrkc8h24ov
SEQtjfGG6VBhV0RPpNZ9/TamzclmWT18m27dYonIcquLXU3fccvoEPD+fbNJlPuM
sjFVspYLhhd9E1S7f01pbzDOHnPiR+hJTAwMS2PnsJC8M5FQE6MdRgkZlOX8b9cy
3AH/MBCQTrNIFKPtSX1w4IesFDA/ViJsKSdJzqRgufaaT4d9zrF8/T2aPxx9uGrN
ywiKDlyZo1ustXMelyMpqkTr4EaJqeqK+2+RCqSDMPFEqx37jGBkHLSz1TVTrzNb
BDfUFikBVFEDaPj3QZedYXKPC3PYHm+hYBo9NOoQxislzOJoUo5ZPdMcoki9k57A
/erhvHDPCawC0kg38TcBwfptyGcXPU0dbsTYrrEsmvb77z118pQEAtL0bOLp9mSe
vbH4aLzxWjEyxpgpuIki2J4wBLty6FuI8YlHe3t954CLijo/hAZK7+ltNR1mh1b2
o+5lPWNybimJuypzj9MLV39NpAjHj/WSjqZFoCFQ/NjyzeUxP/wT0Ll74fuhBoiD
bSzzP78UxiShGNJCK5UE9PR5QU1lVn/kQB5gIuAEKL1OH/hHHSeeKq7A39qpyUYH
waKgJdPlckvGCDSdy0WwOq46d3iKtO5b2mcgaqkbAbjzz44Cr4nST6DIs8YbIMjU
MqkcKjPDH3oyyB+gvLJ8TMpoW8xfyAeMrZfb2/+hHb55kJSdbBAYwRS2m6GcOxPK
P7t3CZk0SsIMNguVi2gKc7LsUWKXhRoh57BTeIfDQJ4hOgO21AFb1lWp3Zw6pTqo
31D+bb+ML/greT2J/9T5kb9HA6G0EloKwVxurfaPvxixSF1axX3VAYHSeQJ0KCCo
Na70fqSTrqoUi+IiPhezQ5O64kSH7furlE4QPXlzHaszC7moCynsRYju/N0O0hal
dSoDoV6TbIXirAo+DMZU2somBAIV/fWmW7gGfRxD9g2CtlKPf1s1xmL5cMRANN+L
ZcGBcriEcO4yACKHXn+fjVn6Ez7IHLUhA5+/nQbF7pkXdv7ckhMWcUHiB0WtOmpY
4cG+wi+mXMCQXr8c2ZLN9mFznnmVYA/HrsytPKuKo5sXqeRwC1N9k4raUAIihZ+B
lCe2MpMwLZJWAK8r7GFvWxdSYe/Tz+65JVHno5t/AvofD9h7vjqosZAamN+TYG2l
R62SKdzIyFywOXJaGMQg+fr13Qo6gNUwuNNsC2UY02Hue9cufBix6McLVVfqf/yb
0ZwsRHn2UpmF3AN8O55vSHL8acXUwR5lZpTwa/s2Zd+3Viw8mHBEUoEQkC4ZzqEV
HnN2BWKQsOoYKftdVu/o7xP2pfabzB4OUTZ7YMoDQB5LS8ES8AN0Q4f7lCAQQhXH
OHjyd8adw8cydopFT5Ea5Dj6js9rZ/5w1lRG/FpE9P1qcoUuNSQl3jWP6c27LVo4
8kQsC0RFkYwAgTPJEshDOl9i6g7p0bgKg8LftVvZKIm6ogfWrfgu0UBSJN3mR8I7
5o7S0f9+L4eTSi4H04wmiLt8dDY5Fe5uQ2rWXwp46cW2AjBIHJ22JhN41ha6K0yY
EBdNurE6m7TJaZ6A9hYh7rUCE+Gu34VNpR0SAp2Y7fm9I3jtWwL9qu4d2meF+l91
YP7nGHkX10FfjwkT4eTDgZt9bAi97PMF6rAL9qxz3bQMvoq7o77FWk6RJmFPNsIA
XPRRkhMHZlLZVSJkkQ/quZLd4dYiDhuPZwkYTTPmYG8XzUULqey1GCX1X2UqWZXN
NA8kQ9FHD15SF2z8VpZxEpZHtfr8P6wI1m+VTUcpXSwkt4AHdl+UKKMKS8PjWcHS
UXlvDwUcDAmGM1AS/OiEGyrYP1wkMs6Nj0IB+cxrL3M0lpnx6HxdpZoXJNnExMgE
AsbMnKvSYRNyvsr2VfWr7EoR2guOCKJY041AL+S9J/jdU76tBhgj46XQmZwffAw7
xw+tr6+rR2nHSdZB8nGbRbzn8ukm2nrLy9l7KL/q1vDpXxDnM5KGMyl9MnA9AMuX
HYR2mLgfnK9/cu31Swjgc901gc20AnkXpsFbjD2BT5WIxM8GPdd0MLOSXy5hCceL
T5TvcWEjPhtYMkyR1mHYQBYg3h24GsCe0nQ0FiaNq1VXzLcqmM8fvJMX+cY0/rlD
B4tnAVwtFc5tx+QF1KtkHlLALL40efsIN75Q9vrdYwkKGrosLch7BQlKiFjwKEZC
D2C5nyW2Tpz0mmC4okWxOiP7iOAMjThmnh9HlFWl+yWkOxzDnb8S5QXXTrE1PJBK
Y7NR6boUmhDmNRQuwnxSb67i0ilwQSQnvXZACE+HEvSJTQ9I+8O8VhPZ3JFWISA/
Cu9aTS0OqFsrQtCTJYu5YrOwVyzzDBx5w8FlutqI2eobFe1xeVYZ1vfZRBvIQCuM
uAfzhESLBYMMEac2978YWMf0oNahhqImnpGAroWqpUPChj5169r7tMAZ2pqHOk9r
u4Xt0Z85CUnXuxVXHDg8bGb1QqQlZoWE2XNTrxHzHZRUO0ofndYIQWU1QS95ohwb
Do4hokQzr8pSr4dotPXNCFDhJiekPUlv4zsnWwqYqBEskVjEVSmK1MrCTlGLuquB
gXcQjJTb0gDbaer5OibKXl5GvnoUFFmWly1ekw8PemJacgDjQvSw8+9jZagM3fbM
WNrjom+3gS2FlHncmiad2sMWoAKx5mx1XNUfvrUTfEniRMK5pGXbYSq61cwPLJyf
y9//nbZLi4U5sIvfqVfKkttH0xab0aQ/qSg9t0rA14FX5L8AjPXXbNaxMx/5rGi3
w4u4s+bXiOsFmOpjdFt72RlkNtNCuqpiPwsA3FPKOUcLv7yDiUQTO5ZV4ejsuQQD
HJT8nGhs4QHcHJJ/pejO58HdXB9yzTWgxZ7uhpTyDAuCFlyeLiNB9nfIA9Rjb0kx
6YAv4gAINR3cfbOE4vtN+IonGVl5zq2h4rUqBfKBRL5XWvWJkOQHHRpYgX/OV6cl
Gj+vZ17qf3cwyIInd3k0gOYf7NyIdqoNpjcc1libh6LMUB9or/TtBrJqeWlv1Vt9
lyBVs+2FccPcxq7v45/lP0/WsPjZuXkrAO9A3+TifyXHq75ltRtG3ifCvNXmrq5s
Kvy5zVWOkOeGNcE71swiKrPD2q6DPihUvYoC7JJb04HP/7AGAiCmiBbYYT8YNSaA
8+es/YqZhs2UDHdESkN3x6n9kvJdUV6ibY38P96GnvS6XKYs8baJtf0MRSkE+zr5
AC8jyK/hLtsaWB9MKjGx10pO0LEq6U1nWlPWLpiqFbHm01BIvFWmBMiTNAvM29wf
O4oKW/6IaHfHS60uA6etKnorVqCbaY65s6swHgf19x1sShdahg+sTwI/cZdOoJoe
RW0Jsfj8eRCYHBy1UNiPcYg18BveebehKLXVeE2gjgqskSRpz5sc6dv2QSr6oPr3
LGx64zY7KceBDduOnAoqtpvlBHcc8+KPXzow449znogH+CTa2OY8BpHSBMebgemO
mwqve2ge+AKj+S4bOkzN7DctOT5HEZLsZkfDltqL1TnYBAbEsQax861ViqBjoG5M
7UeDbKumGnFvELyAx1KcbPTmJq0Ehby7zAegGtbWEVJZZHyS22qKavLDs4GeG5QQ
fEAz4olZoxghXli0f/Y/SkTn/DNvgYMoUXW9xl+De8hYrYofEGlNmsJqlm7VqtlB
a4kD2Ni4juTl1mN7RdkZYm5Xz00AIiRaZ2YSkh28TBKhw8PxBBTnpTAdEs8o8RKc
OOWSYAK61TZms4KFGrVGNSN4g4HMBgHFlQ+rP2xLaEkfAGrrc/IfbRhxiYTq12uB
qpkOfyTC+NJwMEmbsfmJD3lRTdGh/rSyKeaG+OQKk8TElhgEnXex21j0tPWhUWXv
WOPGpWMmXfzgIjK4mTEx/eFxPjW2YJKO/S5QHDPJbByz63NaDo/nOS6jlYEfXQsC
gHiIy7IwI8gnCnfW2GLlTZHbjBVU/L5h2inGzFR6+sc3kUuISKvmhoD4A+vKr/xM
tFoG+lqoltdel0kPlFAPMdL/GYp6/A/fRF4WeXPOs3GvUWx1qKc/s6Y++teXfLgw
BiSA6jaEWJZSl2Rh7Xm+CtWduibQUgNBXz92k7hnVDbvghImTvNwHw8DmuhoyWFb
9FltkU8QomdO8iwV/XZsQnrHaUdAK8w3/9H0x3iB3zFSRIZMegGPK8yLRKO0pLyr
W9M50EMTzvIgEbUnaDnM385MnWp+ZADoZ4Fzd4wDUuZcOvcQIliJkBMejxyGvHtW
zh7bs3LtRLlM4MlbGtkP7Fr9sJzfztvdvy26bF1TXEyvgMDpNXYm8Ljlotc2ibXO
CCAUSwWQ4QejVDCEtOP+eQCkicNtLwFVH7AP1d5GzixXpfjN88GLf1J+d21Qxq2T
AgI1+lyNuRmjrz5wkxTXmhk+6RyW2goJQHtD0BqlDnq1yxewqqmjdvx7shrmMg1X
XYCPEomzQMABWP7UzZ9b0qJk7vUU+iylRb2q95Of3/yh9DTu2ATISjL1xtgwWATV
0g1YKj8p4QnFcNCfOSCiC5j2P1/pJdgUGwS3R6bY2j6Ipoway3XdhivA0qoXfYNk
KT0aLrDmQILikxCcEFTd0ruub58O7ZgCe+jpvudKDuYqThlyLW63AQZEG0tcTW+O
yEfNPIaB1xDnhuuTPysuit2nxBaFBjtzlphXG067bxIGBqgaqVAD/Xo56SsJk2d/
TsQ1ZhlwVOKf0kFD87CKc1GYIFRcxe31oAIaFlyfRguIZ0QICDnJwHjPBklh9ocM
HD08+WGb1GGcBskzltYuAH4qvZh8e0cVJ7B6/CbJ6+Bp7ejs7iWj8eUHIiGO1Chq
QSEyHnm84VzLumFMYKCjeBrVXemUiStCkkUFU/3R98EM2s9Gelf1kgxSvGRA/0GK
c1x9z7Miqr+y9L423b4NOwS5TGIeHsTgZz2LsiRLZr5h6Qe8R8n+nDbYo7zgk8QX
/lTATOfgnBfAIeDCrnFpPGnnjFVP11QJfBXjoEDK7WLaOE+5jEPrNbWNocifZbnG
es86okv/H0PRLEaKyyWgltVPzT4Z3J/zDvx+GfIiz5Xt7M72TvnRDt9XJBWFM63Y
aFApz9leo8JlkH+UrUShgzLRztrgKxzrUIkzD2QWvXUOjXjyJqWfznxTV5qlDCsD
RHEBPMAiId+z42XdJuI9j+RkiMXq+ASLkRiaReLbsEJAUPCpazPLl1LLYiIT6EfY
eHqa4y9e+8haEcSvnmZW8IrIg3R47MD/rSncBuMGd4XgXSkyps505aTfnC6Gi9rD
ZtWaVhSmNXvBIevNVO6PtsLFXzKZalwx18a6dOQn6tmhwI/RSzjuYLRBumv09MEN
xEdOuroJpzoq+8Wok/lZ5NBjvz2iMxAECW83Fu7NmoKWw4OylcqckrPCmhDgfMkQ
xpd+fmeqInVzdALP4HgXf5MnPcKtcAl+AtsJQ3nXLHvG9QovlB1oKPfaakEL8tng
RBLc84K6SnpEDmPxX7W+KWTmw2TBIs2virNEegmZXouSnkLetZt3lvbb/bxXTgai
QSU0stzBk55HhT11zJC2u7Fzj6/MAaqDj5Q+5w0/Euf4lJXwIVf3djkmDAdNyhua
FA8FMK/Fy8C1HpzWwm3EII7qiZA7XPtTQZDGomJ6uNsEP8u/JLe9RsYlz6yfKF/w
+oD4U+z20NCywgkON6I+XLsZr6/zr2QZ3U1T7l9T4J1cM30AAkKvauBrwIMO6t1j
/L5AAom9I7qdgpVPmHWOGvD8UhjsUH0944Lh2FrEY/pP1NvvLdU2051FhrCiCYVH
Lk+4mxWu85OnPSjxc1f7g3pQcCuSRkS8iWt8JsvuqEiIX0o8p3aEWU1ttZp5YqTK
/3eRdzPHmreavN8FTIo73IoP7ddIgsIE9OLaEtkwtu9CgjtMrjp32wPzgcBlG/f7
odCMsme6WODW81IuUbWaoQ88U2/l3dy+dVrkNBvodfkWl+GBCBpFbOP06Q7jrjxb
EsTQhwlMDTKRRiyKqd0Ca01vXMW1dhePqiVuS74lT7fPDn6Sftoa7w1dNWYu7XP1
LAqtZkiukibNGly/09l1QTQW1TLlPs3DhUxHUrfz8vnl96qNu+cVxG+VVEDgGCBt
ZoaJ6JZaKTUJwe8+PDkLva0D2+i5yl1EF1WFglQc2vD/FuXqlOx2hGTKkPbfRfFj
Qw221H/cksokvLq8JvSXClmN62qEVomH/SF0PZgbadg3RZjQfrlq64PyZji6XojW
MFJVI6cHbiwRxIRm4R+fgAFTJ2Wa78+sxFWFSr/ceQ6Gyz0kMuSXkA2oxRMyC68S
+D+cUrZn4gCjBSdviG8FSJceycLI61Oh7gmMSkA1nmsLl5npdu/UkP5+sXC5cjvr
ncYN338bxbx6IcrwRTWCO0mmy2weuHrl1ZPD7zwhhPUtXyRCwVBLV2ael6o8q2zh
KemSOmSKmeR+5oOBnOFHE0NP25WT/F6nbv4tlNfJXHKiMRpqsASFkheihAG/zKiw
WmjmaipI8pg1KvatoSxUPE6C6PadLnNMHiFt7MdlHF1kZnK4dhXvLmBc6abxXB6n
/Me81F5bh06oUAOhaLUMLcDaQsjEPHHJvk6cfn81FPCEID40l9l1W6jMS58jCnL9
yRxANtbH1vhTFSde8wQpTGSdHxRPG4WCnhu5J5Pdy58ciUSW+x6EJ9YZUVY36xY3
OAR8Rbb/iXR/5ABRu6X2BiFNFbXWrm59nISFs4ewYV9V+q1Nv+PdSQHCOpLHLJi+
iWmEtMzShf906/vgA/KkoQrcJ3oycitDn3MqBccL6eStnaodadHCDt7H4m8N5Mem
Y2Zu7g02sJ9KigdZ5274jkibndzxQ2IL33eJa7hFG4YTtaewQ7QBSFc2LLy2Pqil
Fh1/14Te7HxOBdlgRTfrPSIqsLzxTUtK38dMNDBGt3pFkDbdx+NapLGV8Dkq7qYD
0oXOk+lB5th10HV5gniKDC6PKConia6aAClUgaPOiHCI26QsdW+QGz8Zz9UnUHbO
QKkBmwymXXER613Vr2Vp2rwhMyg557GfEQCSfHiRLPxdZTRfZJwOv37oguSe2fEE
LhwAc4iGXU8Bb5f8LnBUXMMcR+TTpU/JmfroAOt/T7jMsPiKYlHFO4u2OttXlhS8
V74fQ8spbWKv6N1/ND4ptcvbgGdrOVl4N4b3EtYPwckEpdx04cs5RfIERVf5cMf8
Fc7JeXYnh2huKzXkZxpL8nhUHzLzCBBraUTScKf9HXf+YxkLIfZNUwFoi4Nc18wv
Y9VP/8gqojHUPkQcgNrQq+L8OvymiYic9wDUxL+JQUSwnXZiI+vNRrhRmUiZnUS6
QvbL4e5ky/QHSwmQuI29jaB0jbGceUhNQtQfZh5hAv0ergxS9nIL/zBuuQ5LUIb1
TMG9eIh9bVLLWsZkhfQhZzYXQmbHRZ6usbOQS3xmBvk6vBqhgyc712ezRwq3DUrR
HiGTXvds3gHxnkyMhTD1Ip9H2fA8RHXj3/PwkJWw0sdxgp8ORxqbHCqk3nRTzUy6
DXZj04N0JxgbyKzfsxFAXcmohSyuz1+0I0NKykc84ti2SzJgnJb9a5ANJc0H3THd
Gx/bK+maMY/AohIy34wF6oHMKazrLujSbNf4r8MYbLRa5Nn5vcGsDzWSavbK1Qxh
LxAbhVOkVGAhzLcowNqwMkpIh+mJWtYakk/nOsu6jehg94k9wa1YWIF9Fet45HH1
Kv9qg7Arwj7bKlLJ6V/M/h1XMd2yGEv1wwmfd3cqqQ18UTM8KNMXtMmnirXTpiMy
I1Qjn6Ein+FwTGbnHFzanv6Ei5mBl0bpaPnkOs68wOjbIoRBt/VKBlBE9sANNrqO
MlDhJJBUVZO7MhTw7tg4cGoCgK/6StOzneFQ4rnE4QofDztAqdpMJGmiL7lxsHdx
+ad332ZrN98j+CgyvYf5VMAHkVT5Y4dWTLDeiPDVeHRB1YbvRSH+fWVHei/yo57H
fEDmg1h78MDPrHGp7CsoIXDRetpA1xN7h2fwN6hB17rfJ/orjHktBaXxSndcE6IT
hAcjiGm8w4J0vGWCEaT2vToEIozugra+mH1vy85i79v30q/BPRbXh9tgOa8yFkpO
ZLIzdOvOIadNGpv6oZbWjAycdMokrL7dee4fiTC7V/q9ObmqlGfUaAm7e9o8A/DB
diVxLwSBilk143jNbb69XBKBWu7RvL93O1MqOuIanv9c73+2gvSTp/uAB/rV9OpZ
wG7BjtDNwzcKOdKaCeJf8++zcIeKSQdWC7OQVJeV/nJvYVrA4det5we03Uldlntm
p7JQb+hEKtBQ2nri4d2TvjvE3MenJGH/mwP6LUPaxoA43GPWbHjw2qBx1cQSig1g
nG0DMBiLB5UNrESPu2MmtGwZaSFMYm58w7Beo1cA4sTF6pwVMzP4lauBvXpWuSE5
+NGqhDVRbrnaU+hpobYUa7HG0lPmNJggnemc9cQqTKQGd0X0dCdwb1EYh3hQPjL+
UWNwKIZdL3IrVfwGgL1J1toaZRKLPgKuPS1ib+z95xjdmGMu4VDxdYAMVaxAZrLF
OCmcFUNPQ4GeaCzWtDwkGgBYtBjvia5FlRC4j3t+5mI/nR0JB5Lze3LyqUucYn88
Lp+f3iP4dZdop5g3CenUrOaTBlVDba3JBsXMPAZ8i07olJbERpyUIFCjhqKyFpLy
1PAn2MppXO7+UjA32/snboRJCphDwpmsrM4OVMMx/qb5pr+FJNq8736rd/SZFQ7i
BnMraKhEsTTDDQwG98ojEJpaXp422Msniu0vAId4HLtcGk6lkObS1RmrNENfa4sV
3nA4QygFInyLdVPWjQaScsXqOrRN02/HExlB5WIy0u8sgLf6RF6FS1oDmQyivuSX
4+IIlYBldo3yAo9SFMnTG+ARRGUb1GW5wnvsoAr6bQNa7/G7NJA+yT57P/sT1+vP
qJNR/KkX2/TuDFQgAIFAxdxL4WpCLMEFrWzUsa2IhEG8N+LVE8QCiaGK7xg1RB3O
F01u/I7hoBj5GDVRw/s/jZyHJeoCb8tekq+6BlCPeSP3SIlB5mQ/NDwaZjQI5ij2
aYdpZpSwdGVFYXSWjhGG1/Hd6xnCyLwIQ+RMl6MLa7hCKZqpy77ASqRCqUHmsn2V
dhdKAVZz30spjK1mBAEr4aqDooXihZWIqqebKLwS4Q/3jdItnKxaATnv/7N4MgHP
WUt/HgB6plI0ii6+/QZYDGkagdvX0gpDgcRVFm5lTckwKVcl51zhljBSI5m/HvY9
/vCosXeRs3XGEkRfWD4/I61yQvsOwc4d/z/Cf77VfCRk+dksF2Utsj/Q6xDXknCP
1xCI+Vt/GD6MGtueLE+IBSS5xVZCJwEH81z+dt3Z8aXhijhm8kaiCPxmriN1/SJV
sm3AN/wuUmuwcG9hzEqhEXeC2jWt5axLdtTZE42N6C4+sI29PKlD6tZZ1QR4xCxN
smRB/N/akUWPZ0G0lgVJAku2Dh/FS/NNx4cCUS4RXy+f/kx93GfG7WrqOPTDTbG5
2st4coru9zux7TX8hIRYff4lI3U0zWEvhnnll8Z2X8bFyQOGq40CUlTYTU+/jl/h
+DVZ0dUQ0dEX2fzOHe8IPrYlIsHDDSZr9O2gpekHRN2Jrt9PJMQNZUfSeP4Y557I
vqGjSmocFLOk8ZW6D5wOerh8UI493r7McXF13I02LI26FRYXnRSQgQ1FZZ3IARIv
WewdYGrxa95RfiWJFxlLDahp8TjIphRi/xld8qzxmHslkz+aDTteDPtyR350wxBO
vSXC+WSFqiij8XxDT+ZbZaTwRGzceUmpvM5LSygnaknUJqXRPfieZhKDBQhiBtUZ
DXpWhJcdNjY5IRPeXsyvjDGQKWZKhUqSdpQx8M/JhFgJLbRuKu2rLs/PyaPTZNbx
G/wjBx+Y0+Mv7T+7/KkETAZvxeBI6xWCOksZepmVaT9JiAr6xQBcvgrTaluFTh9K
B7r0AFM9c1ajDH8WXBhWS/A4ej64XYaHEPP07IWEm9s4GCygzlkhPY/i2Rh9WHIR
uwNN/mtGDJrW2X+XLNTnCj6PPKKLqWRftKARHaX2+1bLmkSxog8h3xqPM534t6oc
re8YlpGxlQGItCnT5XPsbzExaTREd+2L8lDqGkaFRX/gZ+UedTAtx2mOQAcVrDGx
2coImoEnEqeLU2AQ9r8qmSmo4uwGOg3D8GhY333hjRxrjXtT8EjQhWB6QP6QEIUv
00Z+6A39Q5+uQ4M4tAY0DBf80X/Artmg4/0SVO4OEuYFhm0utA0RAx9abE9Qj7+Q
wx6C9Vfc9Gzhlw5KQzfKQSEQLZdSnNq095YFUMKRDmxsTAVOBitEJdZM9JkKvhoF
/5plLnra+wmboKzwujWfpwr3OoPKZFexmrTygv+jUICiqdkKThvGijKNWn+inbLy
kiyQlpL9zHl3IC0HgEfXhE/YuqZjpbkIby5bW3h9vjT7N1wg54YvSqMy/zuW6jgw
GI4EDV3PKBclWkFCtiUaO/u8AJXtF3Jm5UyxNmzGKcTM8Eu3MZB1O2I2qTPu8kXT
1POrNxAD6sz9ALKIiNxVpu8FAs8G4fRtgUyd58BxF1S3Eq5Jxzg37CEX/sDNbp64
tSLuSSqdBeuH37h1WByTfBbsD/KUJO2Rgin/ZVPLCXYKrrwH0zwDPGs4lIi35cxC
+wWd+fuisQC7Y1vHoPWECFN6R/icmQyQMBjIIcObBwySBPhnxIRHcaHvTMDRTSak
/6s+CMYi+xp5wlYEXKqAGUTJgOAifm6ElQzCpAqw9J6IjUtryf4G0Si5Kaljsnw2
ZnLZuCyWQvrD98c8U/rLw/uavkL8wmNAAfEC5HOUBohuUxFuKfpDxigYCVOby5w/
ICgE+6aXEuyUeQhTvyF/4ooQmsq6hWIur0R8ZN03iw6oGfh68nodEX7dwigwchOa
cVG2lob1oOr3B5vE9Frj6Hq7HHmOtIv5J5uDdAWy+lZdVVXRaA7OIhoKRMjeyLiT
xCMYx+jinpA9PLm4we0YmWVhFGUlH4TECTJV8jASQ/1ddu0qyyqlXXX1d6YdPPKB
ajdRvZyPhpptCXPGXb9aXw4wpKasW+BSGbn6uRBss+kPZ1dTCXhNvR+mMMA2d2vW
oF/BkY5Wx0+ZzLQ6RA1YLuRAJ7QiItKj+VfycZqAPLiZGIymLZGj5TPSwp6/6W9h
48SIB0l/+os89tlUnVCafjsZr2xvR4QwvuW3cZCai2XseQbEBGV7BRQR6BRUa1KT
mReAQm89CPoPm/IGiVIokNNgrhy9poDYR5cOwMlqnRNfde7DH6+4BmFHn4OYwNwH
r2o29Gu5QvwVqRfmhnryBR6dBewZVLX8cqrk7/jYcnia9H4cJdvIp7Ua2EqlsTZe
rSfunwVJE7d/X3elzoHqr038/rFcAwPDAPqpCKPzv0BMcxqz77VDeiYEjg32xRUh
4f8YzimVR3biYd40+aA8oGrVYc1VysvqgrtoTCi3FVSUlvPnOQiDVVUvWQ7jTn6z
E1z5eGuMzlzeo/1YZniAVReAFEWnRYJWs0NzImZptqZN48421yap6f8BPWwbaIBE
V4E97/npO3elNyXfcFRMsroSF6DoSCifiUjrebcfPQf4pa340VF/QkBC4Qm/LoDD
hRdDybqiorDA6xtFm2WNIj2hwhd08JKBbuVvCbonwHJgfD9TGQMxPOvYbt+/zamw
vuDNm+swO1UqprYImjzuBeV1R2TGFW7QexeOmjxhSKqlQOa9vzpWKViPheaufS7y
ZKFtHkNF7zWhddXucDwq4inMS/YPcs9kVq4xN/YbFpxul4A+ElDGsD9G/Gd7kU4v
7a46Ve6tvyuPu0pAtFEpAVv1lhpL4GL13WUWlHBLBkzcBdkolRDePg3FC21RyEai
HpKUlwDYIWiM34gjwl+GUCbvDXKIzRFEgs4vTtSwfftrA9nJkZYS3O/zL4px51/4
Ph4EsA/io2W5UbxCjL6NgviV+6hD0KxJrA8Sek0PJZNNBN5/+warKNVzTzcnAtp3
sVltxUXickisfWcnU9zHXFd8dN33p6E7HxHPN8yZNVEacAC2hU6Is8hbBuPumsdk
rkbog6rluFjR39f9XLQ7zdzL0YhQBfUO76mj6LtXw6/BXQxdE5Ec42YWesX2cw4I
p25wD3yFwGMXemUxNrXIp/k/xa5PP9TGjVZcJQaPlN+kdlxZW9kIui6cFTsNmWlY
P4zezozgbDSrFuV+upT0slgsnhwieJHBJ494lEKesn7WrB+OFTbiZD8dzCcJu4Lz
rIr6bw89AJ3K5kuTKO4B4Wyqf18OyWG7tzMfHNAbfSxxbfGEmvtbozCHjAm6Ooyu
zOfti34u8lkHFSkiu9MYmTrIPN2Mzjz38UBcisJwIqTFz/kkaW7TdxunZvfApz+q
Py1LDJIjgQpgY25vY/Y46ArFQJxMrzQ3Ux3MXDRJPNaXod2Qv8NlhmycPMQtYOvt
XZQv/OVLckqJp/mZE+g9Ko5Rt0UZgtfGLRkkkP1co/fKnIbRMAeQRcrDg5FDt7ah
afF2m9cZt5crN+x7IlI0fvVBScImphclxVSNM/keFTtDncEBvG96DM250235TCkQ
syUkwEccEeq5s6VStrMXiErY6cnYT9veMmN7jOYV9wGuH0u8IhJwZPva7uI8/urj
JSsreVQfqKhIbPpAFN3fAGCQ0mwJodklBiUGVOmxgTXEt5ZVshsw1EEiqe8PmqUe
jfPXrbYhrQFNuTmog2V0hSIvsY3imrFbCKnMJqDabpM6vHsRxKqpebKlhJyEhH8Q
23+hxDuMiMwApSOphHgxTpB6lxSrKMgmwJXHyiX3RZtBdOBWtSR3+RHdI9jxseSB
U2NAoiW1yhBGlG/SV0tvdy04Zqfa93jCswMgn7iC89jEBs6gzcGysAsptLCZ2Zuf
6Lr5dwzR9/B6cEnsvhmYjr2fMhSbcBEW0Y5LBMnvMMxtMjSJ99BIiBUgqtzbKx/q
73UPkSuZlOaDSXN0lYZr808jPeWuI0MJnSVR5IqdDRxAdZTBw9CW/hp6zPDdNWJr
eYh0C9rfMGWN/+a4vQYx3KqrkZZlsAkiK4+mk1eNOLnQcZ9xIcX4mO50TLV6YoIp
KnCYwBrkv1jDpbIuOSjn6MVqxMwu5/Wr8oC9vcId69QYFsDlNseWrAhA8kcxh0TJ
KdalR9garreXQ1ntkY90jh+pnjCD2P+e8Ix9rrQ3ESyOzwtZ9MLZMppa9zvnW6Ef
y9iGhej+O1TuMZoHQH5DxG+OweMZnDCdcAx7IrpNO0PzJw3RhsPe63S0py6yRtwU
dTBkPultQfiV1AiLkwee25qWOOryTQW5/F657Icc5fqe2+EAYqXZ63YY1z1ahlFR
sX4AY9+IBU5ewRixJzlf9QXaibmWLqDJ1ftMW/k3ZoK0HSZax/RvpJSvy4uHDLS4
5el6DWNAxBDwnmLOqSTChJ+Pysl3A6tY1j8WKqqZwyDJLsNx8bQMjXvcNoHxEhif
BF180B+PPlnmdgisxJ4USNo2wd84MBEgoQKINdB+wUHaW94H+pyFI1QwsLgkrEy8
aEsFEb0ZOPx1UGaTgjddLtRAiYrjM73eokk0Q9hHm3hxgOM9wRTF7lcWePqFBQEs
GJjIvfMaesHWUO6lFuJ771aKUVRFWrH5wvKldixZo+iLLZls+jnJog5LofpuksU1
fFApDKHXZOjgHimaWUCCs1WuqAWmLLp/ibDORwPEvDopnzJjnk5LA/fG7rRab+/N
g4URfZiGQVE47qPPmANjLHSKSbn9i7KJfasY5iii6gX3+0fKgVFDMiWkLmC5q8Ic
iGYz0Btb7XY83tjEiLvxw6oWHoftgaBFytEZH3t32g/JoSnE5AxPYLNGw+UR/Ec0
6EvRpUjly6MZTmK8j+Pixsnof+5+1UAQwtKaQnNmW86/CMo1A+XpPnyjIXcjdE5+
OBA+aFEnpDA1MnnJRTT+oDs0GMIFxZJgExl8S9nLpsiz+DDr2LBvLB/nZQlKt29L
BIiuJcIxqKZMq94OPGteJfKoZT2n/QB3o0wadQiB8O0+sl65bVnP3s4X70J+U8Y5
QR7D6fzHJSDdMqGfJQ2tIAPQHspnc1V+kOkpKCgUszmof6o1B6GVi9TCkwjjl+0o
RCC79TjIUjRqMkEvbFM5AqwzOLvwwIy3/AauTR9KEb7acqEU8mk+abP5FVm5BAIi
1LIa0r58WvUaFhB19wq2spmOt4Bs3uLbv+/UcT4w0XSy8WMVsyexYBgzw5qTkSND
g3d7xjYOrUso2rQ57PkzXA+LWlYoK1ZY6efc8oc1yo9z6+wpVUkEN2hNjR6CIaKz
7c2hAIFJqfraa/lei1yJU6S1X/FsAzjtsxn36MDGSjGlPxeFK7ll10k3YAXrUSDb
/F05Czq9lw84xx6XthCO6k9UjZ4Tv1qcB0zvk9aSQWXP5xjRb12KJukTYJbdCQIv
aYMtkckKIgs8GelgC1glESFXbGsVCKu5VzkX33i8K+QsUMnbtcJloKEINt9XAysK
TmX7ka01j12UHqvM9nkfCNi2g8TxFG/UBvqKseBuMnJg0eWiByso+VAe4EWoBSoA
jf6O33AOcicspfHrOyNuI655yRSSk7l6hZHLKanXFr3jprupGJWR4VHf8dBKf1hF
pjy79RXt6xlu+4uHgJrbqBwgkVspn2/Dqe46TVqRN6VsoPX/YnHKDJGKPu/LTDD3
nY/dQAy/CvV1P0cmHSrgJI0fYUUjlMUKnz92WPA4UJnAkXjWCL134z9IvtTS5re4
RUOoId8aZIaC9WZufQ1W1vcRZ9fVSsHf3U9Lz4ZnZuPCsCY9Je0SF120Z1ZpLMy3
p/tghvFz5wtfdPoZK/pcaMnqnfl1DhO9mXTbIlvGTLNWaFNsH4aR469pHUAIibnJ
lttTMEHEyAhdLod54sTcUWhNXWt0LzSCGsciOiajcHIo/S0M/IfBmN8SP0TADExM
wezXs8Z0D4GVD2+zxo9wsMSaBzd8xHRPlbVZGd0Qnj8VwACSMuhavidocr925ahM
Fm+v+OEKFV4yZGnIptxhGAYEEg9Z/Jdsn1/Quah01BXpOPZJamUlWUifsjyT95tZ
guKHXQrohZyBlzVpMRIZKu88OLd+IRyMBCQQ3o4QlwT/ePR79MTz4zIE2UZtAdsD
luOTMF//2+neCdeRUox9BrJEw/bqMJ4mY4MP++kkAEvu5nTWJ4+Bnd529UWVzbh2
R2vct3qEAEf7jzmB5TSvKtYnJYDefGj44WX/LPbQtZ+GlEPUAoDn9pWcIwJ4XyxX
MF44bKvfmr0H8CfQQ6cv+AX3qDDecQufUBQRMSTIOkzyN7g9DS1pBqGAV69Xw0h0
YW7Ic7luAMsQHvxe7+gd+q//kxqwpi9QbbfEctUklvc0QoKBiTJHMNxoLGuFu80v
lLs+TNzFHJgdlrfOOlOIV5LrLo3mwy/zAsa1czi/46puT0B+AN+GKhRxJmYbi6qL
Rdcfp6x9ea4nWY8/Eos4ruqJlMAAiCQB4zCzazRCRs2JvydFX0onxkq+KUH8NkVu
9iDp1FQlBNfYSYeGk6Saxm5un6kjqsP2MHCfrwx/ePrxNYdVdwmyVGDgz8tDscmv
5SRV2Z7skefpJq6uOUUE1wRU8atPkqX4s7s4wd+BkjndUIWvn8G3ztMBslhy9BkK
9H5bNaOyxJH2IvpD9Qx4GlWwgYm661T/uthOcCLPttE/z2mZ+oxrNbfz9YHlv5hN
0z2Chn7PwWWa21yOevJHFVobTX3qpTapVjIED9DciP2o1AZbvu5wkm4mt0oylCG8
F9dSJy9ZNIbgP3DqSWBmikvu/b8j/uQSKOcFjHTy3Y2tdGyH4WiXbxLS+31svqyP
2CsESPpRiGUh59MySypAhxqtvhm3saDvhtBiJkTl/C3LVKDi+FJPHaueJUueLLYq
Vv395Q11EBM0YnSjZS1HvoeeJHdcdswY3q+/qN0P8dqk5ZUXoeYFrxSm1gVg1Ker
n7mk6AIU6u/sHQHc0xDdKCno0soqbvvM8MhInqIq3fIVwNc6P8EW4xm6ovaYy3N4
XnYKV8MinZWl/7UPpqx3sv+JIQ8MtNqk4guFZdeQnOQxqQ76lyC6tL2QrAXY1EFe
CmPjWtd30Mex1Cb3pxGFayqFNEQC+FQs6coRVgj0+f/Aw4LBhrjZzdc6cHlSiM1n
TJpDMWaQHaJAcc9qPo8PdZJ8wot8FIwndOzTT6Gh0INpvPYC539e/apuHNbtBZjE
ub2gNVhUKagixoPOhPKcVxNlw+wvnNTK3LkoibRftcsfVstfZxkhvbdnRdZ7B1/i
A4RbDOxAJNTdLwasu0fmaJE4hntW6JPDKxOYvSpnLDTfpnSWxLAeh2OPJgaEA05p
4rWLA4ewuA8yID/lihHBz3oHrKcTBoUoAMCTlvfVakj1yRwU4hXKWUljAQHArg4D
0M5iIID+JFbSQi9WHAHe3nqAPdFGox3pN3MuAviRsB0DjGIK72VcWAM6OyHd/ULS
O0RQ/9vx9VuJ/Qn/swKk+6e9Ee4awyBYmZE3DKQJ8q9En4mMutlEdnShwcnBQG+k
QsXeNPHUTM48eOynJVU1vk3ZXz4lChyZFd/IiamQtnbrHX6ogRfR2r0XJreAbuzd
+/sYm9ozH1QlDlIbBHyO611Y0FunNIvJQlfAgBiaepUH3g8kFxQ3HKB/R+vICH1U
9hEIsIpVBcFYZr5hYMwwxWUtFKLOsHfCKIYRyc0Y7NiiVmCiNguG0wmf0Aq1pRjC
ukCftDxm4Zeg7Uo1804vfPlcl/NL+yXWsWMIQVVcHiUKv3rDtkCwsxP263JqJ0h7
iuXIuVScleyYinKRm+9FYWvvIvUs/er32Jn1kqBBWxpWnIbxGiNPbIdwusROqPql
2Uor/rj16NJ7km9+5T6HL5t7pYbo6lYDPUxmjAHvOm+1qbYMasHdjl74AnG7Ahls
6nQBG09Zfjmjtpx7jBCu/3DRkswmxJAbykidEUoC/h9PHeRiN3zZsDNP9JGJsNUV
Z8Ld5vt5q/Wm33rwZ6zsURPXsmr+Z/yR7ARPqX8T43tOprWV40HZ5Wc9g1/ZnJOj
h9LCh8Zi+igX5Cvrxqrp8d6q23j13aN6p9O+v6dhvUWwSD2hXrXoPf/A7WKqsx2E
Z913kvGMjjG9p3RhKSTNO78OFc/rPEURGfnDWspWd6em4jLbZKhrkU+KlzZUUK2q
PQUlH6RbtpInaZi32NeC8GgXcW7BGyVFbHTmfD2k+wVOQ1+knRwirSYjCeESur3K
JOd7+FWVfDvBkXkGUlM+3Rki91q5iYd4ry7e4R596III8NToGOaOxfCpvM/s9DHL
a6Kam1xXr6DfzR2lHCmxMmqmIabz9vfIPx9Mw3QeIkpnKabEULUV5VQUL/dhCsD0
sT8I49LWMYx3sOnbFltNPRJRjHoBkx+5FgoW7QQMJt3rNh2Z1Q2Nah8sOgRTV4WH
GjggtmsVu0RAt9X0FJdgFXHbVAigvZKZO8kK+4NC3UwVRiL7dWXc+zcsbXzjX+Sa
OR8qF9u9MiNdvxjvDTTlBX7wzARf8nEnhoSxIClgxUzV+nsnrqNCZjj/6aI9+A/M
cljrLhKpRQzwjVn8QbwCHdL1k/dTzU6OnfUGmH/BY0RylFg68/Z6MpGsAgK3DEC2
XQUyIVhbHQVWPhMsL9IIACQ8anX4F6tsbI55B4MUjt36kS2Ujaba7wnc/Y+jA0A2
00uGYmviJegKDM2vOiLX5sfX4bVZUf35HKp/qbKesa+lHZIWwyAeN1ByWXJpuefR
ZpbMgaSg3i/3dTBz75dr/BAl5HwQdB4Wgm/JUi+b+9h/fGJpOmV8/V7n6fZsBe7w
cK84fsLkvIFXNcFMMHWF8O0wMGU5XQb0PSMtYPBGYxmwFCfwuS0WuSBkJSB9LDgL
s1ZO6J+5x4B65dAQ+RhqcFa2OlPyBMzbNS/lbMYv1qhkhxpvKTJEEb32TCQYWxIu
ex6V2Te7n0dO2pIZlA/mcXIz1/LIzOj5ijH363w0s3hDU/BbUNuGXz9iRpBhCJ2m
BEhYWk9l31fix+NO/HrrddvNYglwjss/oOZhfob5kzXoewm9JQv097AFGYn2zJvA
gOyJr0IcbRQj2b2lCs8lvAceYJyb0kIN4oJSBt74WIxV9R3muXQOSwNEs9nsBsAq
jredS+8bQSeKlJQk873UmORxzLwHGwPIq8Pn1r/gKw2Y/revz/JxJjfzyh4y7Jjy
bAk0Y/tqO85/YWo6XMyxKQO3IRjBNU+Z0t0cYSmAf1oJAVWu58C9oDeNJJJaDgrO
OvtvNtJjePromg6x5HWMM0fhvHjhtVbFXuW+JsVdoqASQ8LCUnfsNOmTSy522o6y
6siyURslvPsobguJki0NUh5dWloFy3mx9heV5foMm6KRa7reqMrgzPP48n9LS82s
Q1qZ9bdN+BehdUTmODZzZ8uIu2EKDU6lJit7MK/mSmpKK3F1nieSuz/4toCpvZBB
MJe2e497U9gyBohjW3pxTkpk4jA0shwoYTwa5sa6lLxYBIT8hQiI+kOgDOde2Me3
Dyt1ZDeuegCIWDLYhfBR82LBg6Q94AvuAJZQT5lfYJHjh/Z+L22OIjgeoM59dWZD
qgErpZ0DDQi+JnFfYNwCJQ/IyoR5kloPrHjPJjyV3R4XG98R+W2lHole8c5l3lXk
lpXejg8nm33iS4xbP3ZAS0M2eY1tjsj4u9rE62A1Q7d55Q617WIi5A4sh2YQNKTd
siWH+R5180wumDRvP6nG4xG1xvNKOhfzljYTDlqNs6V0iWfb7uvIC1DXvbVlWStp
QztRCzbY/Q8xj5E/SlZmG8plxfxghOrDpcrF0WPC2kOalehlufh/s0naoQNPqO3C
FCrFbZqrrvvPQ/vcy+DfNNxKi1VwSXv3rqOQBG+22CDwAT72uFCtdhpQYpRmkLFX
x/YjJTPcWZL0avawD0lCCg/uX1X+79G83FaunzM+ebNE2tiU25bZYNCfoPKlxO4e
ShVQBJulhNdyG8vngSdCc+iaeB990lZMEfMYxlFYANC6hSvD+BzHSiQ+qN0IQdgK
1BCMrtA6RX9hRRqKQBKHizrlD6+rf/P2R3s+BoLLkEnjltolFeBnJrHZpk+2CRVb
SkCqAt9UDO8KtpV+QHigj4ceA8l1t5u+LWt/E/OF1Fa7GYUDJlX4ixTSmqpUJt4+
mO0Slv1tGuRuxFz8fNIT5MYvs1ob3DBFZYLH/hmE5hu5B5g9H7F17qtC6e2BrS7Z
xFDWyBBe003YmDLC8Zo2fQ0krpByL6DsTCQjaJ33acTGJdtZ/X4lG+tVJKQ6oHIo
I5izEY+dLa8+50/ODEOQntp6UmO01fA5VhDVnjHIfOhX8cc97llbyUcST6dxW+T8
jSmdAZO3KjWxHGajZY25J8iCS/VYK30Mzzg5xJwEnE+aoE4txWSHk/ql1A6+nJnQ
BiFkl9ENU4NH6fJXTBW+nfsRCt7JYpSjC9BCSDLzrzuePtxA2G6GQCfKckGUX367
heXiLelmCrHG/emSGidQuInKUqfiLmF3x7W2NLVzyQreZEY3f5a2321f+UoIlBsh
0VLOa0+QCrAukyrtRkOv2B34POzz0C552haOeKR5oFrnhJDs4g1ndi+GZMzxoH6e
hbubimlciOwR/Ch13VoWZXemTbgIALgOdDaEZR8/mSFz6lIGoTvGSKefhnXj4EsX
JXXEMnO0wensC+1vNrfFe7C47VgoonIMfjkw0m6k9UIuxCYJgV8fWYv9hjTqK75U
XjiX01gPl+gvMHdd1PG3vZaWHm/tX/Ywg7wHLHd+vyJm7FIJrlCHtAudMw1gYcJ2
9EEvnr2SM5fwuCQNvxcHZDn2h6eIp9z1hws0RuzzN/R8xkfre7ftse7LhCj0hPZT
3PaJyJz5355c6iNvY+639C+EYXndrKEGUrNuQVUZsmBQWKdAlOwrhy4DNo4FH/hT
MWHbQr4Po3smaJkgLMJEULCDlxFdP9gfpQwQCLom3kqYPiCK+7hzLeex69F/cYY1
IfkEKDyL24BhMkAqw36DRixcn0Oyu70RuzVULknnrbcP0QuNVzlkHwvbMCc/aqEF
SSlbEiRu5I+u1wEBjYp458Vs/x+szJ+kbHRXadOTlv/jB0j4I6EgkKvRA/cDHIkz
Ojhh5C46ujOdK1II5J+mCopzYTRW3+PXuzRW8b3e4u6YZr7+hWnvWiMRF8ioxC7b
aooKG9rlnHKcut/lXeFfzfmhAeobkPo/ioazDwsuJLT5TFduH0JgthaQ7wTMG/83
tZ30O+PEsf93C8MFcHvsGSgVZYLR4t4IDbbuC+MJTTzCbhXUe9++OWjtbM7xSedi
frydwlRJ5YzkdWUMzFJtUpaf+U4lj4eC4Du/8MF/vIIBeL7zrptY4hjopinrzmwd
zlS5KJTZqH5oUjCvXzeRT6RGUdCCKxqYK6JD+7bblrvuTcgTA1951A1p/uW9T65/
k3O947KZlURNkJxEmOSjr3p3H+2csunQCI8Cz2chrelQQuA6j72edVdRSZenaxDz
RedE4Rbi/6dz9+2fRFlJu49Uos5SO9u65SYj1GA75bth9sGZh0FEKhyqGndhw6NE
rtuS1WKOC02OEWUQxbT+GmFqcrXnZ04A8+eZGbxN+La0JisTVUS6PuMVxgHq88o1
mMVfkxEmvW7Mg3iSYqBbNGfHsYWE0rHX7wsR4a4AO+nhtJUduWZP4vdkSaRtSM3+
GEXnxYKXD8WCb2d2O+6P66/bBflvC/3EWMAAZdO3tAEgxLb2U9ohS8w9KXdd1NLR
xy4OPerWyDrpj1NJzDQFs28Ixr0B8lZ4Fy1hZMc4AyGHLnUSBNm/I337S0UswQKa
WolGTUj8M8HX4gWrN/9qKj1xrUzEAdFexLu59u+jA0ZT44qpCtqqfc0dDCjM1/5d
5zjfbVCPlVefVRh1ht7PaUG2mLwWrz2Cf0lOiFJl8fMg4oCnl9UyjisO3UHjEdUe
HV99gN1toTnrsoynspn93ani/3WqCLMhAOqHuOPb+h3GG1MNrwizb251bo/BycLC
KnUMrOeHL2ftpWM24Bo9DQJ3B4zAKbCU1A6za/ejNMdT7XL0g4ql8EkmSekybMl5
g+h0hCSclVZPsMqTlX/lH5z4i1hWDKgRJD7+GcRjapRcJ4Gi5fwfPprnUm8nA1OW
oOHdYMzAXUakJIH6x7OpPAPqJNFL1i9cfFW5PMKtoHL8XacaHlPD5NXICOmm4uXT
SksAUxkBd1cy55nVBXqU9PVbpQyfLY2V1dHhW4nBSfqsUFhyArcvamKA9IqPjTem
/AS9odmT5KHPXTiOc6wQ5Zj0Cn3zprpWws+O6SweX5iGDVBJBkoLzxZPdUq5kwue
tytneXV9NoLHHq418TWCEdWqeKNjeNAB8NMSYkU5O/PlqUK8yWHHg4IgbvFh4CUn
dSzqAqo2jtE5FtyjFIIfbaXJfC2vhNMQzElmhj/wlIp07tC4ZD0b2ld1RlQWMeXa
iU4s1Q2rVgS6whK9nZXYZoRkOtwr4G8BGL7ZYAWrX8j6s/kVKzsrTwaaSeY1YZWp
adaIUx/RkYdm8tVqJiBRQcwfImfmAqww1fbT3KtrDxmCDehSVfzKlRbf6mdxs54F
W/W304UTTAeEwo596xFhR0mV35iT2Z+0NijM5xEvC0vdJBGnt6Pjl3lbqa3BTdAL
1fAdEkqstLgJmGCWdFNtsnb85CCbiL3sFZ3454ugpPaDV3DzjGOKWrbL6gDmsDQm
82MMx+jO8mpb9UXxDqI0BgxpIADhXMjXS723rnpKq2YwxeYH5Xbyk1pInBmXpyVx
lkqzYawcWosQ7DGeCWxb4s03tCFGG7m+4b/dgDPc80ku4gvpPRuRxjyAqaBii45j
mXUvccmACZrnsAhRrHztjaflGMA953sgto3H2An5TC8864393EXIQVi5vWvD+rk/
sP49b+WjWPNfLM1F75wC65SxHrXw7GWOchx+L8B9wmRsOeND25PMrUgc2gtcqEfw
zzQMF8KH3rCGXeTuNxF5K1PLO8rb8rIXQRBWqPaKGkkDPGaMZOtEzKpLGtVwoi/P
g52+Jb798e+ck+5oHe+5rxPqMdnT+tWgUnkpnWvph5M6frBY03YqZvP2QIKfSfqp
A6k5AwFQAyDV8M09ctLjJkh6VrkAWP30Ln5S8bCBO/eP2UMo0ZU8csPUqLQnysAZ
+Lr7BNLOUr9cvYZCiw8+dpAOQCcgf5ZZ5ilmMGMuziXps6IaDTJinHtWiZzv+El6
p2u0KxJlrFcG4IrqY4kjbhR1DzXb3AlKZNY5Jey5EPpz0nec6gcqHnUR/zE2Z7fP
q02jYw+EKrEdWEtevtcXnrJqKWQOVraH60e+poFi51oClWoWqb79OPUth/nZxmrv
mqQD9dbAoLAb8M9mj63hqKBpuka14l8yLyK1tJq4ycpjBelyQaWipz15l7xuVyT3
b/0uU41gBZbrRkoXQ0LPQLBcsXQVAwvGLWhS7s+bipZ17oBtzuyExC1QBDh64ftL
nGjqnDCgo1ZvP1M6Vm5OoXRmpFEeyuy1VFKXEEhxb7wz0ipOwUuMYFBQF3YMViM+
LcGCeZitErlXA33rJ8Qp1x5IjEWv1VIhTAIWvUJiZC9rVxVdXm1ww6POE9BCBGnX
AgrJ2p5uCL1jwURUQUjl6ECyfBDMdI4by24wy8NPA5gvJrfqm3NJsZcVHsf4Jh6t
9YY/W8tLE/T2EBVddV8CV7TJGAlC05fefk/F2oRSgQHy+41mUaUhOF2YfVPx/3XK
7yim2EklXA1wB5XPRI+U0R/YGtp6pQHqNJdJcH4i060w3TKQm5QpQfNiwoGJ7ekM
Xi9a+EICl4nSBkkjRiMmKAtK6ClvXAI3et1+8t9bNj3byOq7nSaJj9AfMqNENjl4
3ZpB+Dp4Ua6czOnA/xpFLF2sovuanUAaNizh2kpXYRpBieK9EFmnAdXjAiyqspO5
k+HyhBzszPfXFrptNiicUZa8CfO/O+n0R8VZRKHAtV8p/wxSryWVrn9zHDgDa23y
LDjZY0dUAiexAlKwlZtj5OVYB7DgLM+xAkbeA09idrsSwhLrPQJ3IaZ+o3MRnB4u
c/D6h2/WTuvUPzexhQJ5vaTtDi6z9JRlTNg6BGgV+IUko/2WCr/aZT7MvkoBpvoY
pkIhxqgrhFfaAUnuEIFb1MHN8LhWMWu5pNuzSvKrS2r8XGDBot5HgB8brSaaKNJ2
iR5pCICEYc0lVMnivwDlsUB15g9eOI4gL8cgiwdpAufg9lTt+MDN/DZaPXnafRMM
KIjOqIwrjpC/HdhvCAJzwzx84Gp1Lu1bqc65tKnWgaiqaL/AdoaT9igqsEqTo572
gF+bGAAcMk8tqPzfaj66qIvlHmEoWW9z7A7FTT2wowJrU6Rc+nJ3h7K/SvTJuPVQ
DWJlNs/2bqearEjSC2Ujo/LXWPBG0jkTR3/X24WArVtoTgQQIu/0nKpjdWVopkXc
uPR9ObUMFRXUUpv6pKN32kR6ehne90DvnCQBEE3XEWpN7NoqMLdLS/B01sTdFpxB
l+qnmCOSUWMTfk/ksn/UB5KdES/u4DIHoxIPf5Ybd0hcL2JLjfY+nV7loQrnOff6
bV1lUOoEuW5XX527mAQ1RHrbRzdGPpX6R3VEaNUJXDM1OaTufgGmhoiO9mDxMS/9
ILJWDE6EcMrxiEppVAqGILIQaPiasTNJAd7hF+7wiGFuayv7aNWblrfgs0sb2DJJ
EaDQ8bUv7WHYaGV37dnrPSWjkp3PANKr8qOUi45yLA4GbniXIer/g4igvuEmPqpG
mK68Jqj+rNup8CM6Zd4ek5FqnEajkigFtKja92HJhardEV0/1C4/bU4H0neTnU/g
lia9fRSluRNMYYSWaI3K+JY0X4dMW3Z2ulHtHJOGsJsb0BcAUpQslo0g7KZGUxj/
txoFJQe3nfQvG6+qfv1/EBkRPNzaUZ8TjoKgpDDyTo2CNfjLyDtDfWen1diNBXXg
tuUxbEHyPgkF9Xycic1KLlqjYf4I1h3V3KOJH3BU0uTc+9DiLZj5GZ23vfjiqxbh
1GEruLj9I65XrqWW1ZdiMUXN6HJ68x1T2m+frtbcHrHPrgHDlWuHqq/d7/ejwRfU
MA5qLQN0nW7FbVtkvGbyRTwEf3RQu/bNF2S+wBUJ8Bn7/WvJLJNfachwQleH+g2y
5dv2YJdZTO46mByKd8UiNWuZbTBLVhRutDoFunAy0nUl4jdXtN2V3wCppPbtjihS
qgwygWzNyHnVv44GCYp0uDwCcGotTDT4ST1ullyyl+mUB+Yp+psCiOTM7Ar9555T
k+uq5lMROKN+vD/mYA6NnWWhjfdGUCIRdDlGV3hbcwa3V7lq7alzStAmcTNlX47p
LgxBuOmTT3H55q2L/6Cryiwu+D9G1QXRBEtT6WlSsDGTO2LoaSKlnBL/0OJT72uB
4JEXDQj/DybHl+ae7FgmnHTEhUNjqkzjQ/5GshDbtymOtvZdBy0zKXNeoBISAx6k
ey5m1b2TYu4QFw9qEozkspAytSmPoUfscEDkv9mDY5VwXKrmvcVWgrLla2XbitQU
p+l0GdmmkWURlnfVtwLIu76VZg+k7yb/HTEffXTGPtpm41fGCA9yLW9A3fg5unWh
M8TgovriYc58heHd6e7P7Jkmu7cQRglSwC9i5kdlLFdmHF3FEnj3Nd7Xw9jg4NH/
7nzlsSaVb+2BEhwoToh+B+0V78v7f80f5ZU7/1NZdTBMog+yMhyl/vemVH8yQ+Y+
7OOWYmdl/EckGfO41Gh3ucDpSDQXo1bYzEuH5lUkXhNzY1/4XPdwGdRgfe+/AcmX
zH/rypKyQs22leNz8cq9WBOyZG0wvWu3BY07KkCOKQT5i8sGaIAIdaPwnEJ7EdV5
QZIkT9KeryvDvthkoJs/NrF3byrH7gf00xh3MgSHxIte8+qJSKJ2udcDJgvdpTRa
hLXnKLr1KRnWHKng7OQkEV7MSVgkovu+KNtIEZHKVgTWTz7tKVFby8r1ImvD7jla
HG8iuRFlLNGWSWgJ9aCvU0de2dnIJSwKyejUMt4cWyL+oMzA0YaBqHTcl+miI7Iq
GVE4Ck7Lg7ppO9H5cFuoPcdvwQUARKw69dVZLfO2npFDc3QCRtVfSt7rOcX+wVyh
NF73gykAy2NZkFC/XWF0tr9bvF8+2hzcF5ZtBAx3Lprsu7VwJeMrQMnsn0YGDj7L
E4s+wKW/eR31Jyd1pR8ioVCc4z5HlcACc8Ilw6KBuyiLIftl3H5NSTTlrXNeYLdQ
n/LlLth4y6drIlw4vozCcCpTAbMSI8sa4pa5/3N6kK6OsAl7phIAFAVIgVs7eJYO
PU5mfN4f2/je54WuSXaUIOD89VtJZ05SrEmRUBuVxoHty9NUg+srTn3tTnBAnWgl
3lIVKxQerCMJX157hXffCW4poey+CmKX2GkVYcYOaXw1DavKSBLtNtSAUXrfhajk
DphyIpOEpSlAXiW3CvYz8dKXUK9J7lGpJ55bzSny2C8rjy0uzRW8akLTD9spu6cd
HA6Lhb6yuNn5aZNun4LETVRLrvsPU7/mEFWKjY6uRCSldwjYF70m+aHRSpcJvGAr
eYkgdP4793c+2iWo0YaCrMF4kFNKjL9yrE4GZKyJeMroVReJ56Cug0kp68wlhVFb
Zwq3/PXFTg1JmkIAQLVTXXoat93Ld7vZcwX1uSMDRE+pjxF4294KzQzBUG53qktF
xe2vtMDm4SKbPd3a7LPKW+lvzBrupMoX00QePHTJiouAZ8v44WNkRIqc9+6ego/6
GjKW3NJplP/zlgFzF55z1V5aizi4LDPcrjMpkrW962zfKYpZ7pSXlQ9w4veR016j
RibV7r9LxrJWSUMrMHqfMkSMF3mY4hHRGV2AKsYy4UmvS5uKFCNxzrUMH1Lfa6LS
rbQk9tx8KcdvRJD30P2W360voUpp5HLWPxbK06SbxCEMRhmOlu7Kt5OzLErwGn4R
IljxQ5hM2MO/jLwh1ITl4I/38DGOCIUopSgI+fWdg62dg2ox/v6/52px45icWh1T
ak/6XluygRaV6r6R9ENMNT1Oii7yqzqsn7FD01pjRRhaJPikLZl4GL7Cv95Dl03E
hA5MZn5rgZ39tf5R3gtp8jo5f2GAF/8zgWpw2lYAsd3riv3MWvSFUoU8NQ2O/38o
NQ7eMQGXTqCvLoYcdiI6enNbRr5weCagIYAsrdkFkpMvW9bPGavjkJ2hhDlAkCGv
vgafo0mIPpuKw6V14CQ1iWQXz6ADeogrS0sdCcGfWilYjN2OiuW+ee7mJolFyEDv
lKIWNOqR8V2dyJFKp999CQLEv/ZHFUipd9opEZ2vRzNAF+/q7VIxvLvG+VLJUUtG
FHObqJMgAtR8dXI8OGn2xHdCEf/tCmelxHaYUQZf9ygjozHxerjunbDdkOe2q5qn
OutHJaPE0tr95kBSejzSLRicmkkdeJbkDymlDYk1AuFxENE0wQhANs8IEteeCfNt
RUVWpT9RXkEH5LpBUHFsk+GekyQC+QZSLr6gPeaMWZLlG9h/gHgN9n0egfFcV9Q2
KGUruwbSyfitRIZi+Hwu8gEEl7OqUXcX7gOyNUTSNgUFDpXEBkGd4tKZ3JHtc55+
Jdx5IH3X5d8ZBXgfI7sFWYmZ5tbwsfmG9T238Z6ecZ/DfpQHoGK4ZtPaXy51KZxC
Fcrq0I2ww9cbIQekC2gBwYVGBx0V1FjshvzdbqjK1kpKHpeVXFH0gMR9WtMXel/h
iO2J12Y0+rHv8IrRVs69/Xbe9RbV58EhHI3bNSYqLuSsIVWa8kLo+qDVYeL+CVVJ
nfkcdSSDH8EjHLrtLiVkeUvtpIPIHu7HMwa6Mk75YrYj6JCzv5llwl/dhw24rPja
Aa0qZedTvw1nvv3YzXaMhSbRmYvzBh+3rQ4FA0TJLDAA1Y6iBJ7u979iL1XYdLaG
TooCGalSUa0Au5t17wpXM1R6RwDjWnkKMlgesQc7czJBLdrDvf/uIjB2e2VLXppa
LFFYqO2hfu+kz7sJp9s300maRgnNeIMsxkevYf2XUthAIkZRJcYT/a0F/X9ebxxo
X0beh6vp+3qQh6CrwjdfRWioVjPryWc99bmUXaFDWSA7r6IhgH7BvJSLLnZen0kP
7SGjz4wvzL+x6PBZhyVPZoS0elVKMU8vW4Cu9UkdEQ9B/OgYedEtpAwyrAel0OFw
6BXIu2QfNncPripBTwvAXhwsHCkEdeNCQDOnbxSc+iQonUL5XVnYXKxnhDBi/w4z
atrHuetmG+DkbwPPkS0f4XDaqSQEjLiLb6p7T8L7zha97oxQrr/2sArfMIUy4ie5
JzlCHLXeuThf8YGTXkC2H43AT/V6nRTBzKtcChrPGESgqaiHlcE/zBmW+glVBP2u
zA63ZOm+HN5GmoIeJhBrvUr4lW/48YSkzKJgmsBVvR/F0dyiuTdIooLXaz5yajEw
93A5tGrFVrPP9qIWBZQDRZawqALxxbI1DyYxEbnYOxZin6AxFs7ElKqUDpijT1Rg
O1kPNeJrt/uPoeb1M75Q6MGhg32a6EVMxk0Lv1+Qi+YloqINtdUI+mhnea3DrCAH
eUkhm6sRB6E0ZwLrMRF3Su0f9tGhdfkXGQuJrcSYdRBmZYvmaUZdD2Qrl4bt7b+X
1zarqVRKLYI7I3q50MRIfCM5Q7X+dRX8FmW4kfAhFp0lkZ+tAlM1DQ5HCgzNsTIx
vcQWfBYDi+Fy5zjrsJKaj2fn+Ps/zqsRrI04NBxqJckB1uEi900Zvwq6ZObtW5h0
chlHcMJC41T9c3ZF/iSUJrGwIvKB8lMWJEmhwhXmXD4D2LEjCWiazbyTSS96UfM0
au0GhWO2Lg8JwjDOIVSIhN7Uo2Fri2N5t2TT3xWR11AcCE8w0EbLyiHO1nhax+ut
vMBfExw7Ab1gWAbWHirKohPEvlpzMl4v0KdSuTgHbephRxiAiu+ZVreUUcjJOI8b
GMdxAOtuM14IN8fM2ZY0vOVost9aJ8ox3nCiRVDCn4VnJqQksSCjiIhX5WV9rXc2
nw1UjQNpS99EN/Zq8gej+A+TTfC3VapPVefeLOA0U6K0cFyjJooB3FWAcug1jFb0
tEToktvJ6jAq4kaTMsYiAqPokgcCo103tUqxAZhu9Mq67XU92CF7s5X4eB55ZQUS
I28iEs4TTCKBvgEEzdbI1XEh4vK94BlpTdcttLvewIhhkiwF/UHqtv/TiMxmcSpM
g116Z+0dcwIxcSR2BzxvNabRUYoK6KgfWQbTCvn0s5ieG23x1rjLGgJLsn6c7lx/
yWBOcwrUlz4TFksp39FW8X5K3xeZEwI2h751SFrPQTz4nehpCfepwZqxn1kkrGIC
6VCOcY6au1xYr/ETCQDfyfpSVvl798apKd23/tehUtOcVbNFPZ4gd82FrsmMfx1M
hcpy03R4PbRg6O6tVeAoaKlA0P0QE6QEF7XZpcr6f50dWQt+GDk69ubnlN9SJYlt
Q/qdw6T7NssNOkZ2IknDgPxOxaCsW0N6ho+vwbNRflRjWXx3lpyNkrla/VTbRw2v
uqDJHYdjITaJ7XyRI1zr/FJmIjvgZ2sl5XWomzSCKx5N+ITYOj7P725r8pXYMmjU
W0Ryk6HD/iHIhoEIEC0pTIrDU4HIRbPBUra+1CcUlpd1Z0Gk1oxcIYUPY0K0//GE
mtivfcSi60uEZxOeifWs4OoMActGEiNHuoCYIyE3WjSFrQN+h0aX+8zpAu9TTaBb
VTIr447b0dcZZ6XSFq2OTpvCppXMUIPtilagri/xAB43Zw0Su7ypJ+YRSR0zQoqK
ayHrAITKWzt5GDyNNDaT3seWlrC8zkfOHcIbONwhdp6R4FwMEnRNVcetpgxfQC9j
LEuxhiHaRJK9/EwKP6gJCICbqaClDU7UJafJvwy+BUQcZrZAFSbTm2R5jgX1fJGM
tSNv72setok3hyMgVVxIDgAPDwzNyYvhxjrCD85xKsZ314VoOInqAS8bIFANt+m+
yt+pg/UX7tliysogJ/7W3AS5g0zWU4ptvs5xlm4A9muTRPfF+DZgS7jZxFafmLCR
T7nqCreo/YA3q1zkCrHJJTbqgeZ4XYrRcBaD2BPGK0QoIZ3JQOn6tbYu7qAocQms
hQKrLim3LNRDArNltQ4KX56b+CwmezvYdkK7C7DA+fG194bTiNxJ5Fge4ArVDVyW
pKLRfTU8e8+ENQo3sfJ58kAqIUvdTr5ZAGuY8hM0Dv38L3N8HeSVAhICdhBXt8K9
E+z4e+UGFs+yzSQCtRgfi5HAtFaOwo4K5CHdq8b7/ACeMi5tZLwo2MdQpnwwgxrz
LJNYo6Wp1HilgK1cjWBg3liyzwFWc1NnWegS0NUfyr5zB+4yRzME4uyaWXZNrQxh
7OEeonCAIGxyVh/bQl4ljoqsi3mEPotUcdtOpPnUTpPBHOFFvuk6ljPifftdnDoN
XCHnfIpm7IO9bZzy/yjRI+Ba4qYc3czLeyJLZcMFzsQzFkXoq8MTbVNdUllzL0zh
ihGwBwLWmbisebpn0XRL7+9RFR7/mYez6TcSbc0Qe9EokPgTvXnu1NFVZImEYJxy
ANDy3+5Ztln0L7fMPWIsHZDkvBSjtI35l1WP+kmA9vrnnK7zbYPLPN8C/Mdtuw5x
mltm45T9AFU1ZvtxwE+iYySsvjEKM81HBBB033y4wDci8DMvpn9KLOlxp7ultVBw
pTL6pSxUrK6ORddui4WxtLNsz+StlNPm2w3fnxuaW9z9WsintZzZwqy3vkZi8Vlv
CX1eyAYCYxMQcVO9LN4xtkKOQn0tWpvgEfhVHKGRZonPkxC95ZupUuYPcB8IaHHd
/tSpr2PbabW4Y81pjwVCFQIPZ5mq/874fhFdUIb/nyqjvclKMMgLGYRLXVpJH39P
LaKjiNTolxecI4DoxvlOqqRgVrPmoC1cDhl/5MrSJvphO1ZGq5OdMTLeqgT9/a/B
UcjCNx7pzzEg7n/Bqm26PYd0WCbWCzU5IUo/UKSPB3bx83FM/thRMQf0MLsJpLtq
Nvnh/2awronYclBmfQj2vHS0vIsomd6mrbnFQsBFxfsWIonsOB1kQbWQG2L3QbBQ
9TeyYCEOSuxjE4ri0ZHfKdUs4l3h4tZI4/75mX9ruciOWcDs0kuBXfy8OX3JYFNy
orITilNqpTYi59u8QHQvIsIC48LkE2aPTD/7QNbiPZ53E0Bgt5ux6rZEJu4c/bYy
OgSoeYwKx50QureXDK18VdCs0/0WG7zOt3697aRKuf7JyJL26DbfFo7oYIaZn9Jp
EhlSP2MtJOc6XtRfJ9qiwNzjm+YEEkM4fmI1VmtbFhFe04MuYfUDEmTCVUC7ACft
0mV7HXtGmCWgp+ZRFdHwFtZ00lOIgAsNILu+2eTUhQUDPUxJkjfTuD9Klq2oj81B
QhC8RWnYS+qkjF4IrR8c5pTZu0F+0dX0OkSlVe0i82o5S2N6RbcPb00hN3uO0aiH
ZNYufb89aPwYLpDIjCcsePny5W2ZBNmvFMCtlCu/f31KQCGHryPWmR/4UdupQdrU
IbIbEgMkc4XJJAhInfh/A4zPC13egCrf/DSPdaL3Rb37vyBh/RBdDDfG8xDE/ARq
6+hLv9dPcTJJkdpfiNCnKFnwSWGDAfYQexbRxn2UDuE11mb1KYWUbJX21qM9mo9G
eGGJarODrxYT0z0x/dcci6U6M8+MXetyJpp2cuWIA+Iz4P+DfbcbOshxbJJLM8tu
56sJzDfe+fFCxLlKCuMsqEJ8FoBLJHr+8f7q8Cwt7MrFK2zgpVYUHyMJ04m3+mXQ
OrgIcywKYHnyjY610Gbc57VJT2ygNmWhWi3SK41SDlFvD/aXavC+hyB/FtIUkBEU
kvBKueHDYlqeKrANpGulbNB0htTde6Vivg4FEwqrKdvD/rn0xypXuGSt10XPkJWX
tc57F5FgdQezhTvMTx8YT/UmzyOMfYZyzrpvBaeX4VDL946oUWgSOM2Iy4T3ps/J
nF877xsv6cvYDs5nRrjXPwpMFra6/jrESFa2Zri9awSqrpBOP40y5oIg+ZYIXBEA
6UEJ7xjcoAQzLsqkPUlzvadduVwzDUHcsr8vfw/qfqDlC+X0wWdl72YLj2CSYH9w
YcwRTLPUoOWY1T9sWTcK+9MlazzwST+PjbFNIZkRX715zE9tLy2WaiCTzSSFd1zi
1TwZ8At3wWMxVN2QCQK0t0kWkrVxpMZTH5T/7KCZtKlR/go6CVL2To+O+gmm4uDv
rLYbzrNgmlbvnCH82W+ctwFEHU7r9jozmkEFyv5TRj0KjPZA8MfFnKC7O9WxYo01
fCgfBHn+4ew1byQOweGyQ4VgtrmTLxv2DrluYgSMXLkauuBb/KwMQjjAr8qmcUzF
kOa9wxI52xmo+sU6biGMhMHt99thoq0dGpT1xPw8FV+6aFiYl9lrYcLqpBb0QfcK
zzHufDDbiziUYvKjpTRLJQRc/mVFezBGAPr2hQAAdPjbnzGqJ5thYY5Yjq3s+jFX
uI4ikd3xq+VsqRnPyaAwNGloCYoYTHcejhR7vVfhjqzy/s8cJtipV8uHURe01/vp
ftLwOvfyzF9hciN17fKH6IBK21WcAqzEumEuyEDfBdF1lxbKac+6Ta9rM6S7z9GD
I+9klODCBxngL2XdKGuHvgxB8JGpp1dV3plAMQ9zQd+zo7GaAINXW5+VVuLCCFDm
QnbiBHlj3xONlOYx3NMftW+SD7mMnVhU4Z8roOXyL+ELIMGfRM5MIfaylP5cyFci
gUUn+eyiUTAhz7G3KxjJhjYixVFIo12pQyShBEnv6bRHD+4f2sAnrNehkQ9laan8
Dwpz8Rjl/vR7b8gJyPEAXJnY5exp6wVLygFFGpKk9Ef9CKJQcCQMDLdwSgEfqtPM
JixwQmuu6XwOWOZAfjNguHlBp2FxrzT58mQICSIImjnfhQz5HHlvmUWHJydNxz5a
unJzzIPBeos2M9L5Xd8SDeCLIYf5mIWdYbGV8OdFOlTV5KrysvXPliIqvhIRU7Eq
Sd2P9ZO2Qc+mlnt98TFKRmAFyrwCmz9x9xLUqkPIPB8ui8SspzN/Hxf6gWdOc+CR
SiRnvn5Ro5LLz4pnphIIgRhlrv2IV/OLKCAPectewRW/8ln55wLyKAks3vY/1ZlM
L/lTenR6OOsp8d2OXBkIef7rNc+d7dLC4LUJlG1brX0nrFfWvL9+lPs8uMYOk+jQ
l1hV6R1Y4MYPVg46+l0d48z/+QBzb/iLQ22z7GjA4a+YVWuYtpt6cd45wIeBmT7U
krtKOGOJ1s7RYZDncn4tlcVJgwT2RZKYSnel4pHvX9gIjn/F6Xcpu2HWdep5IgvD
lrI/jXyNgaU1dpFeuWY1krgqN4eBTRml9lv0y9IRZyqjFS4EAPEHvBkMWTJqCur0
ZfgyCtSZUoe2wquICE91QF3Z8vHZKynasUAdU7836ilsIh1ALLvnQviuguk4KNIA
57vM1DWOKPQRpu7ZkTLmGkNs3ENN/BKTun+O1myF/UYFoZbhWtuUgeyRUZz69402
uic+Vg3t5uAqPWlxjVcf0Ir4TCFimSKAqMw4G7+sjMwHqH7+cjKWh5Bz4CUZrJFv
y7Zv0+bTtDW6HdeerEq98RYaDy3HNJcgBbU7CnQ8BL0ZLSwzAwPLMS72bh6ml3Ba
Kpn08F9gqOhwfEf1cg1lkMxyWHhTxavFxoXRwn1GtyQml0wLNAgTiv1B9oKXtPDE
AgS3YDCEzre8sOuY3VLyQtnmjjBEhmp2CjawnPbWdKadgLK34ewT1SJVV4dG+FzO
mG551QTJjxWtyAGZvTejQrdSyDNo0Ls6VZz6XqoRYSxR5SFoX2VlFOIF6rfikzGM
o8lQ8P8sg43BxxUYShsN4qDoq8DvTOMuOJs3wp68bkr8il1e7345GxpSU0z3Lk1T
yvCyVWwny7SqN2u0YOF2Igb6P53d9oWpGcLL9AKXRpS9YusDwqXOSEAxia2Z3NSb
MOsUt17g81lJ4lGG9A9dHOdMG3XIcuauyvtqZZsvfx2J3XCC/G4F/0FBFOA3yiiE
a2wF22npjNYnGbqkhMunltC0QdD20GYmy/WneY8yRQ6OZyixegc1d6e7cTL09jrp
KJY0OJHKRHmBImdgPwjM1UmVPYmurpFlDIUz0Y78atYkS7DRFch7OLb+xiwAwLKC
eUSvcNnEmCAUfSW00QtQOPXc3DLY5pMvlQFkuaBkx3tibWLDza/7ubaSe2h99Iwe
kdXByhQnh02M219XDGKaKFYKdhn9tezraRRltoii6FgVXhkrqEbaD9f5ErHAHqrW
kUC1npgKe7bdiKPerWkK0HFTngYgIrae7CBK5nb4W8eQiKings8dQ/39Y9bOJx5q
pbrSYLvQZmoqGRwGD6Ft5qohwaekyJL+dOpBatveFUVvne6mwhyEWFmUv33w0Tt+
Mg4+y1dHlhEk5RkFOgYUjusSbL/rd9wts4wCbOsEKICjxVHG27aQVEeSapnXKKGb
89q1pzzkZldT7yczFvD6WW5RRLuepe4AQa8D0sjMyO+9PaYEMFYyEBPbvQW5yJCy
4o3IR1KFBxGGriM7pYgCVV2+OFvCp2F332608MWNG8jj3ZjKhGi+swC7En4FeuCk
6VkxWkU1joE/5ZoO6eA6QSENPkc/KUdbGe5A8egBKVzG/EgMowng85g/CHDUYIzf
Fp0DAYVreJAjk1IeRmgCXTSEcfTKmIAbii15fgHfaTwqVEljCcB1fK8iuK14fcd+
XunSWRkx9jSzYGb6zH+2ajXqO61FVcDYKqDsKL/xbYCHg6SAds3LclXA3Bi3RAzO
6T0MIfnBVOBXxK2aqgKd8An3MByzo9kCqzUYB/td5kEkVXbN8bcpofIYc2+3I9/Y
bL1KHN7eYKJv1WOtbWIFd06sgl6WFYaj8F+PQPQRy+u5uNO1W3GOnLIBj11Lkqaw
yMkHBAtP1mk9MvnRHya83OvZtWa8W45X/5+lFRWSKMxLbGriMfnDARZFFaur9wlk
CT0eR8RRoKDTQsl5+6TULENgyvZkZh/dBSBzya15BxhJU82mLQBQYH+ceAlSRJVj
kdDdffWCcixsKh4bJKxJDnki+gU9eICHXdq9VlJR66pYvh2qNLv/YkCUTtHGlj3H
GkrG8Jd7cq06yu4TDtv70OdsjLHRwKSYZMGXuiWdIOtvPdI2hlIBZs/UJqHX2RS4
ZMVbmgrBY+PL/sMT3Bz+U7ucNbtmJtJPNJle+vNumZY5Jci97oUrtgL6VcYwxEdd
gmynl8aa6VuSe6t8ClHupOGBlyzxKnPuOZM30AqH/U11bF6XeetuOrIYcf/Jn6Qr
lvGEcrKj1PeUGHRLhcvi3sSxJNfF6py32oXrrmHWmPjGSq+OEQkS7vV+MMRBZBRU
VOqjmErRUOBcVAImsG59yoH3UuYhcZ19ULG8RzjKWDp4lYlpAWAYBwex1gPSC3nz
gYZtVtDjTP1CPRa5R2cA6iMk/LqWFgv2jr7FyIDcG0gAtXpqeeRcK4TozNrKDBQY
NevPyZUz3qNPdVJ6qa7jPp/fDxjyJTbqVPgO/FM49kDWbueKWYHdG3KEA+IUyJ4B
rj6gZglhI7WDsT7au7Q8ufh0HuWOIi/AeLbgib+osbTfA+IwSGGgEQbTJi7UucGP
Q5fwIMV/f/6sRQKVp5zvXLAIRFoNaky22TuOEhhKqVjkYtV26bhKTMUr+6bO08A4
YL8hkdLAsNuYpYNEB1Z8dyBl42TatBzziOrePLVotORcSNFPs0+QuhIT8LZn6gtD
NJFmCqNu8UQRrFzXEJ7c4YkInMMCwSytb0lyNc/WNl0hUoY+Zav/rANSUw1cz+hn
4G8wEoM4nYUprm3n5B1NWEfjh5A3hqFx/acNP6PFWZsGoqswpIMZ7QtiFgSLUfqt
0gDWv2u3c/T5EuiLs5XcP0HdXLUy0Mn1sqDFobP1vs+GyHXbrSiQ/0Fd1dEYMLEJ
r+4IADW76PXVhA6vqsR1o5FLX0AQnWe7l1Xs70mNROPb6F4z/IpKkFK54MG0xhY2
Act+4lLEgR/WxfxM2wTMRGcUMmBwrcVvuaG/elxQ9SvUkS6BBxSjPvIBPD4nk7k7
Ix/Pz3+f3Vvh0Ch3FM3g0Y4okjx+9mBvSQL4EyW3kOcvBGeGed46sMAhdNdzmyS1
n4XFjY8PVkV1waPwSHcaBg7L6VsOKceEsnhWLjkZXGl8/ddm81R0ouKlpqiYnqaj
IkVn/EVWktYCm1DUoYO7tYC6bgNncApkw/hssuxM3U/cbnltHFvfFqrS8YE3QOZl
twOj4vI5ulpKD6tQraqlqhHgMsDVTEHgEoTlWiCs4HpkjOPaoxuTsKuSVJ9Lypaw
xDjERwrf+n+NjcKJQpgUZ/0tT91CuNAiqZeV2lGkNDiTZYF0fXoMTiWs8XKysqg5
b1zJq8R6J5EmQayTqEQnWA+DIi6QEZofPshpg4eq9Qgjr7tNcKCHPZSAfYYa2VdV
6e3ZpsjgAZamicGCGQz5KNYCkjlw1FSJWeaCY0kobN366ec5q7Kk+nJud+QjrRkL
s2V43OEbiEAEZMSnd39YTyMmxhnP9YAZohTjGV+8k0Md+lijsom7NbhGXu8Cn+mS
MNEYDOPeZ+EedUpPNhwPs0yjC+JW9LzOwY6sR+y7Su6w4hQf8GD1+nAIZHnwXFi0
s9S3p6IlT2BtTEnlHDQRLpKKNq5m7dXEl5ze7mpacsapu2sX+s250LRfmbT1m8rh
G1TDUm2erdBNXfAKVDxMCDvuBjg1+33+netP/BxDHYKfHc91OgQQLUimVi7oT40e
hrQq1VRHwEPTNS1WJwNQxJDU+Vd5DrPubJS1Bq4j1YbEBuQmoykieFWI8SWtDGD8
AY7BdkK4qmcjCC4mlrgOAxitJg4QLFO+WvS10/AkXM/iAmkUMQr24bGgzAqCWx7V
XwrlJbz0y2XHFfIkf4Dw/N5yWPPHNoM90brzs7/bkRmoz3TUzVii90AuCgZ2X2l2
iRWR83+UVEc2OHnVCUIZ7BlbtyOcAQa/EW2MWxkSOQ1qsRwesaT8E2Ixbqb+Twb4
35BqIcyvhJAapqnaJn5rZ8RVAh3IbcTHXy6TeFhVKFs74LHHOoi/3ALITJOZx9KY
a7w26/dEdULBOCP1pct+K9dE5hSaFkVUP9SGe1VYM0lyLdXyHShb+xnQioThfK2Z
TMsulbogGj/jP3qcDQvkMtccit3Im5mwHnQQWQbDI3Gcz3xaZ0E+yTZpBH5rmwX3
z1WJvx+q+MRWcNZhrt4bwVjIOAKOiiRqehZQ81WyzoMfI8kI+N4zr/gtA0Z7Q5RA
aGoPx+OmYZ0kLOkUcouByw/0jtVVRE5AKdewYCPvyxtK0aM/pLY0wkOCbE/M6cH/
9+nhKXFVMtulNl92tZH5QtqHa3V1+LRmdyTlvCX09q1qj911Fmq1vdOMKE9Hmy2t
qbu7/LIcPYUv8PyE4ja82qdj2kqADfLor8SlJo6WbvS16u0yhTmffbuXXu4E5257
WLr7WakHyPKO3ce0V/qAAe8e/FF/udDG3J6xFALh7Bm/VxFXv4xFlF1KQa+smpC+
xphLo0402uae9a1aOiBZu6q/S6x+lFA6iEbaohjY3gMEN9IvW9FEbksWophSDnk6
QLeOWX4w0ILx+7bGQsxcb0ZsPBUE5z72EsSVEIaptvu3jPJxIKebWWHQsKUFvYUC
WHtYX9UtBqUzUdiKdt21u+93o/GLMv0sJFo8zXHGnQHGWA01a2I96NiRuWHTWDeh
QPe7Zo/mcKgDOQg8kV8+6KbCvlE//mHUXnqI2M3bIHSmPYbkCdr1/o1Juiyx1jPS
FoCDnX1o85nHAFP/Y1AkvGySR0QNGk9W8Ns3D8IcI5mONdeENcQ5r3cGvEbQ6dDo
3ldVDm3XVc1l7vBUtP3vo7Io0hbORn1kCGca8YWnSEZLypJvfBp8tbHMX709IdYE
Rm9zBN0nZWtJWZ8daUaf2SwM3UfRQnDqrFtHqc25ydSmHs7DB3AUDY8u4Bewj+CZ
EHbVRnHVeUgA3lqt/8oqCusHnmPGGLEfg7ohofmPW9cyBOoXqEfh/B2lSwk72GRR
Y+59/MGWY4UK4Lb+FHJxjLVFqDfhQHLUdgsY2Z/LR4rJIqmqQP8OOeLJNyBF/oEZ
k6hTr7mcw2r+yqOp2xuK+tizVwyp0QHnndr6ET/wMp8XzMcPJElN8v1XJf4i3vWs
Ay6FhYhypAxxf6B8afeqIMnn7ThZK0Pg05W0YadOycwgbwTl/irCC/6LvOKG2zbZ
wLodE1ZvKqRXDBYAArzweg5bIZWk07YVJLtrhoHlppq8ENj/X4VNgk3yyg4DOjZG
Fnun/6hq2vOSmo9PveV+loy0U1aSVcUJR1mIrhkhFsUFAkVZ8CzefJSp7dSNF/h2
mty7CxdDkaR7rHzKBtZRQ2RC+QQoAZe2ldky8GRX8kwn2izRPLbzyvXAIOasiwuz
+T6YRgXtUWpKwH/8cZF8FrTOBnY1FRzs71rd06xK6PgCcUcA52KWHjLAW+hgmefk
6s94Hgz1q70yGxOt8HHBeaGU0qoXDhfnfQFTd7o/8YB4qgdy2QEHARGqqfAFSFEu
2x/SUMlpefXljHH3HITVZy6FYKA14AMH+Stm63HqTjb++1eFI99R66MCJfGJVo9t
Y23lJqE5NYLPLROm6ewI6SRRHElLZBBTKRjCFLNoRJVv5KFA793mQ1bQsKF+LTEy
KOG0Kj8UufBgsNKAN6UyJKVP5By4aeWNOadhpoB3El7kG+MTJEnihH7DrC4am8p2
Idf5NxM0MFkMoXxY3z7lC1IMsED45EMSEka8e6kbgd1IJ8godyrNxSlCc5Fh9F6q
wKvbL6XFuXeAqWVe9tHNOFjhbCyjfvqg61eFAgrb8v/NzyZIw/J2wqJOmeo5cN0x
2tmYSaoobCMoY3s6lnEdlvZ3la1yZxCelv5+hQruAXS+3iZ90xq2Tj8pi54HGKVd
DRINah4ucwi8FLmyC7Fl+WXSX+wceafTtICq3Rn33n/aBEdy/MqkpILi1wvaGJtp
6ie4cvlAsu1BzpJnslLYMsbLOFa7X4uMJNAmGfCefkHUkZpkFh3B42uTCKy2V0FZ
t6DMUv0c9W4LDzTc1tU6qnNrm5OvDiX0G8/b/2sPsfLKAXwVS2v4itkySRG8VNyT
hFazKZaCTs1wKyPbUMvnN49X9y5C89Q2YDEhbIfn/ZC1+SNLZ8yXuHcx7gJPEaso
baLMmHCs0A6PqiZqBOTDksMXj0vwaCyns4hZHD3056pQsnRv3T49HXklkvWyrCgb
PMnfZRXPRJDMgnzWfyDsDkMd8imAGRrBwpS+pMzoen7BQIVH+vtyJ5Xp0g9R/NOd
btTqaXhMYm0CsiG2Z+jz4jG04+FL1IW6c1cWWVjXyRIVkUTwG4cbMyoYItJ7AxlK
xBZjgngm0C3YXZapY1ZZVrH9wcpnew0sEU6ZhfFLyKv5hLNVY14Dt41gBAB7vA12
OoOPb+RdmWM8CsRIVF2zJlvKzr9mXXZW3+FLgZapW9ZEik1fRH/7YxlxKnmzJ8cD
yjIgJtcbfprvslzdGqIG6cRDmOTonkc0ma5QGe6dHEREA9a3nA7dLewKujScq0mv
jdBTPbGQt5y9WRYjQFioytxi4VvN8T8qxMoEdjeULXtuwAYBNnIqRFFdaOVu6CBT
zVdW2002DjtsG+Zwez6uLkvl6hvC4fvqQOT67KqbMn/9Cj/3wqnlMsYj5ARAj9Z2
VrY759p5K2Z9TDCDQwbU6LuplAe2JgVZT2+zXGmpr9oGEjpP2cTPWSthOFL/DyRf
GYdrrp8eTVDQw+ZDXSo6EixrSavm0Evq4lrLNT3R54E3pECTmciYHdzCAlOJtNkS
efHJ41uSQjf4K7K1XZspQe5AjV92gxJcAqGe+59dTePElOLzkMIo9f4UjRcGCNXI
Pq8ZFyufGYuVnU3SkF5bLZ+W/TyySQgPADB3MD2taDiltJuAyVeNnQhjNl0jvpfq
shV6on85oEw2G74GitTrLcayVzWmyRCRku1n7LliFCKWHqIMpOVY7nQBU5prJ7Ry
+fPe+U0iPD59XugbxhHH7CfLcmKR28IBVZhx7z1D4o1RN4K2HFysGX5WiCMhkFU6
msjc/gyyPGtF4hj51MPcxqKQA01j6QIo55+bWlNbWTTemjiN2q15YxCQW7CiAnb7
JEpVgw52Onju/15MWwwoV/7kYmEfnzr24BZvJKhnQrmpURK0eu+zj78AhVqdWQ/1
5HAM9Rr2XfryXyX2bCvmdFqC6AMppE0vZC/nMLRPt9goauZqUpyfVkn5ceDjbsEe
BuSd4ijq0eHT6Tm5O/OwAAB57rRScPrS9v4+W9dweOJrnOaDrj8zyuHmRUEaqkoE
BSGY856VKvZphuyWUpPvm10AdvrezUkrHpVcTHLWZaQ0nvTwx/qY3+TqSebhQy35
vHjKZ+QZOoXiNHZqalQVBhHhG/1RQG4U/rqaEqHUtR9FdAS2Pf9RWTpRu/HPmNpC
5FvOjmFBOZJFpxl+uvHDjcND/KkIX2tZhl7X7tnUxHj7LAi5YVr6IstpwLH2A5A1
OopCm0V96oM8JgUs2NPMlCULCk8xbx8FxAQmKnadFBdTH61Je3r5SJLS9x7i2zoc
d0/T9i4gtPP1uJmpcB4fXwLPbO8FHCHKX15A/a0qXyKLjQndb6BXm6SJjUwc0b3W
c/aGh3W5yLY56Qdxv4GZZ6Bxn6fi34tvg2o3RsjX6Fswv0UMY1wCnOe8/BMKMmmq
79zBxB6KgvNXjEG0pZBSJVexOr+DcLFh16e3rTL3GTP9Qe089xMtGR7qVpM20o8u
eZw24eNZPee++/o9+7WPjipsRwIGqXf3cqL6SkNC+/3E2WroKYVH6HDVd8fnCgto
icDggxqgrBU0vDdyKxTtFuhmza/4G2kN0CYfLeVZfpPwOjSo1fkTmj9R2qgNPdEJ
+xvvbxFVLR4ViyEAmMEkFbFoJGXHrWmC8ff4yqugfwNDsVLW3cyb1kEC4FzfzUI/
UU3y0mzvIsTJIikpgvka6UUr2sKqw13iQjXG1QiEpOGQg7903sPWCQa3Uzoruqck
XuZMIQbfHIMSVEtkv27E/Q36QakNUGNdSW468d2Lv6D6XSq/wdaYQzexMA+IxIyq
2ddgjty1QO9LxHq18Icx/tVf5kE6MhpGA6ntR0OezYlEPzdMGObkj3eGbpSR3igE
hflMf1qEGpWodLT3elOAhE/YraU2BZsE9V/P1mwqLZmnT3kY2hx/jVo02UOi63tb
rnsS82+BlM2Ge5bT48nEA+4TUpms6ND/3ZEmMXgL2nDudQU0bN3CiSZ1WLjp7UNE
RdrEYws+ezhZYNGZEjDLqDztAXj0VYuklPxBFZBO99K6qfATSim5zBkztHVdhKmf
Pn2bbV6bbQgkDP4fKw4jBY8vKaohuDn7s/B+7JYQ68SMEhKqquarcN/rS2WoKGWm
flQK7NSmzdsRup1FkYazm1pS4Z5gk6A2ejL5LOTXUe9m+kUlOEQiCN1LAjTLEIvT
+dVsFMWM3YXn/dv5eyRdHfTWuO3KM5nUymsAxmpgIADhBu2+nJF27D1SBhwvH0mQ
fi3VYPGx8tjynUJ78K0Q5b6OMHTgEuBQ1G8pO8epSeZm2Ls0LURAL5mVPHkVbN47
VUjdWWgmflBiesy02+Vt9YGqMOWY7SLuEeNgxrHzzE6laZTBTbY/B+SfG3uWq2uA
BvIR9Caennu4vrRy4ufCKXaNya4vtAD58oL991HKP5CrVF+okOdwquMloO+S3F4J
o7NGPqIaL9uY1yYbs7ACBf9bp6BQBR3IDmIb/I8fjI+wyHUffLNlzqzdQZ9Jp2i0
AY1IGzpUqyKTx7ll92TB3AjZoL+KQtQ0P6FR+BI+wPpZxfIMfvbk2JZq2XNxQ1yh
jf8EKWjtgwWay8G6lQeBdTHIGaj/UTWu7b3nwsse1zCtA+8AK9zSXy7maqPYzvBJ
bRmZ9lRvWwzFqLbrol1Waw5m74GoWaGism6M4mh/MLhMtpjUxKvETmeqTDSJbMBR
XnbgYhBBmjDuA8ZFVDjSwT5wBKFCpQOQHTBL/TzYSamjAAiJ1Ugk6IWNrluBMPWB
/YWJwmOyitvsBfserKwEYfe1bqIjQ45DVUc4lDy3fDLInXddyNm/eiYWtocnVsMi
BQoGZhtbMqNrE9sgkNJkQyPqEuKa9YAyv/m68iKZdZtllHgz+YRCq4lCAxCb87iJ
+DgBprJEgqbUUm73Nfa8EPd2kHeZWrXESmdU3AyZD9o2EAnimSnRCPw7q2uvy5iR
dAOnylFTe170rB0sIwE0iNXlSuVt7JLBeETADzMHD5Zo9z9xbjNaLcjl8pnQvkUh
FBVaOOOF4YG92/MeF0DEd8uV2puiDZEpuBL6ZGHgiFg6nXGwmsEKZOZ++U7lDUUP
v5SYAfQw/+u0hIboqQ9K5ObV6RU74zK+DMrhrM36Nxcoq/pNueOYTErTNKalKhoS
IPYdm/sQe9n4ARKKgurEZRM3Dvvf9wDsnk3MwIDmDWY3/NaL3wW2sfHXcYHS03va
mIJGk84pKMmiLGW9UnWIYCvjREDVy56UY2cm8Br35XlZbspLjZDTiB0ShI4bzs6F
Z1DDMrnJe0+mFeODgY5PhuL2D1UHjisoJtEII6hiYe34YHYm2erQ2De6EDW/n1QZ
vg8nL9Xzd8lTzvNz53HQNtDfZ9JT2aSdO9HEd/RLo4TI2DDvLjZQoJivNnUa/oqh
QqW7sIJnJvE+hiR3fhZU+uw5lLxGICpvF632nWwTgzzgFhiBhxrMzrXLb/sLY6um
urnxDORua3LbqXGyqnUXE/oriEmvXxyGHPNuu2pS2tzCCv9uE10sQP+fhjdvJ2+Y
ROWyRYGwWK5dudV4Mu6DUnA+SZ9XjyWtw008N2UujYAmaz49Q/Wkbw7sJJ7+QBs0
IuRN+LA3vf8bE/owO4sWZvzUUq5zmWY3j3LHzGZqUsiNBkRYRq5XK1tsGeVJdrMy
I+8M0DS7sxNq0QRlATk4XzJR8BNo7F5A7k1+D0TW6G0zkET9Y3jj7RAoEHkJdIPg
PICRjohf3Lptn9Lpnw+wArjAm9BrrMd3/LkBYOeShtl3DHubCz64PchKIHB59Elj
xSBdvkbKql9mFqWPDlDFDETfJCsejWfQkQNuyuIlcNbI+k9xhoRwfgAD9ejrDAo0
uBZrRNiQWQrMQkQnVbt0UIBRNVqyxBZaNzZxkracxJh4XdDIhyaMqZdxrNooPn/H
+BxKsFtOu1X00wsJElSL7rUHUP/8cJoBXohU6je9FRlAGDEaG+ludlYBh0Sog0uc
qGpx2BzdMIO6moOs9mWwsikeI5y+XwqkxwONwH/S4E24EFq6OheFs6g9sQQLZqYj
nDOSNNzAdm4gHcu6YEkqBqO9DOYG1aRoTxnYaxmpx/50zfhGppt6UQ6pJ8ZkEh1M
d/JPOnzRm91HEGlQCGwV1CtinLwe2Cz2hqgicR0fU50LzoJq/w0zYwGFZI2BD4Ro
q/841+NSpgMvE2k3IkWkkUQzMSb3TbUqekNarQH1MQhvdTvep9sAJeRXWW/I4Ha+
jEzweQHNt+1AhFOV14+S/LKGezTYdJ5D+IWpm9CdDln1Yf/byA3xlBrbjNq9r1S1
LQml3uq5CLz9UlDxHh7jkkq8c6JspZJu8dSepLhT+Ei4nR7JerYhmSlxzpMkk8nS
5rGEta5ebZ4Ghesi/Nr137lyAFhm7SKU9EC6TCj5KHC/emP79HQJluj4b4Xly+rT
Vdbrl0DtVsQ7l/nyRkjXT3B8cfQ47FIS7NiHyEN5xEY8BSlqNclglrHWzUIADJVD
znlSguQDRggHOWS9q3wq03KhX0Ywi0cXwTeh7FNjU35Q1lsBxD9zMXGTrpeh65EQ
Ww9sjQjW2lFmQAU+7WWRYuW9FAnGJzFjEIymTXM6MItw3zzqu5UmyZT6oT7ARzkE
qqMs0dkexA0lN4OZ/HHcnFEmrYC5vZESlbU9XPGsC9mWfvUwwY44YFobuBH/LiDF
ozwUb/VLRCKpu+Nc1G89Xdirjxugm4XMyEXBKr/egbQ3XuV29K9C9Oq+T1KqDdWA
6jKrurb4yMqNuGUk5tO14TDYAbTky+ETDIkwRWdfyoxoGKAHrZyPWshIcKWG6VEr
9klR4n0JCuSB3thy+U8twx9Ps7j397oCV/wvseXXzDX/3sejPtQBx+eDFwNeIO5g
c947EDXLX2/cMebzOxF0eStrVIOgw62El0p8VxAhDjYDG9/CvEd+dXPW97T2IYth
ixdEKLUylHWADZLPO7hLxzpMDkgfWaEuR0czHR46bk7RBBGgQxT1bIjXSTtSi5+4
Yag1c2mNUCcmbVsPvOrkZLvVbMUL+fYFue5ROTlawqwUtl9dZzkgUJOoW71uxNo/
Qz7WFQEXDMnBZgwnGiK8VMfx4BEnsIUSQW8EkG3AyKszVpl1YtwLu/wbsA45Jc5I
+eQ4rpFs7gEwhyK7E6HCRibmm4cAVr1AJxe0g93Zrl1+RIIb9CytN1NGcbRrSP0p
Vqob99efrtGMSTruTlq2dhDbM1Bmuh/4Jk3/ovmFBn8YXdUlEYEZ05S4NBJM1ZeD
LwRT4YO4MAfvXGwARlper/kbO6aJ1tAJ9n66c/oz3guMI/djr4vjrUzRn0uy8SV0
PHbJh2cOqzCIdg9MlPb+Y/58V+FkHYdApvYvLJue99wqaziy7HyS67UZCRpevuh5
IaBI/LPvKBGFswKsIjczm3HDTGWKGxwhXAqH9OpQmgPNifLWHNymtq7LHRL95tiA
w4FfonFP3bIJ81UHW+W+MlMvJQ2u7SjLsG6/2mI2pKHdxHk0ODZuBPTW8gDNFLNA
p19sy+FL6lmdBqeGb/3pNGAuqXOjOAU9/8UUx04XGNyvIN72Qv1vAh1K5wJQCN9c
XWyNjIvYULylCYmtao9Dv0yTc9Qo5vXn2zuzMGVv0diO1yYI7u2jzVCI5fdOzQ3s
ijODBl5OB8iQ9ao7Hgb6ANqGWPm0IhN2H7YxTy//AAvgBaK+SIWEHqffdft/QLo9
WWHoMxN7XwqjHZ6K94/khmlgqKgrVU864UmmXZlycgIFsxTSZ+gLUbw+gsGejNke
E0pAm2FNLhhBP2NHNQy27b75hSmAJbRG3BWdEkEhsZQaBrNLT0SUVXk7/idbSGv2
QEIGxaf2caEpHh6UCyHVvs/2iv9p6Waw1P1kQBVHpYbtVTuNiDYUsuPaKb5W2m0n
uAG4c0S6w4LDvLcDeiyQ6rhxhEF1eiTrqS4C3im1AAA6kSaJqA2CtZX+as9vG4g8
OFp2LTIq4pmfCvQAyWCxoRN2Ykhq2YazVVkqRRqaADWcfuTijT2zq7J0/iJQ/GaW
YhinCD1n618Ko3FHTygNzUtDWAZoVmvn9owc65TKT7d98KGR4EczPObRgfmcyCM7
y3Nujn2pPM4R9XnE1DKEuZEjfoWDK16ybNy9TBZQVy1oM/PtwXtzSh9rPagwdvwv
Om1blmDzof+B5hl1B67OCsBFQbf3PJ3a196HqdbiBvPV6Eq3XTr6ocu/Y18nMcs4
6vNvabKRDCwjrwMox6FTRpK2MscN9UkEgRQbzpKkU6Mkc+Q2Aec2mCtbl4tNYfiH
NjWCHCDWydO5nwi60aRfDgYErbvlqJQ9+dohXjpRIAuLYXxyYsnOf8qZIco5xkwG
ZmXtKLiNe9hCZl2FyJjx6kyEhqkoSQnmR7rLmg054VMk3/q181wwPdBVv17hrZzc
8/kCsLIpvJkRwbBeS2U5IVhRS4DlMc9FJ1bZY4b8FmYHwiMEbAjhN3sC60r+mehI
9ngFmiSixfODE9CmVp5Z1Et3dstnYjLOcZDtjQyzxTDMnCNW8U6Uck7UQMgmYebm
itgYc8F3W4bIPSdcE1ol54fYEN3QRayD/8ceQ2BixuBLMNg3qwivS5gFwNhbaBaB
Eo0OgrKMdwRLAQCnXiso+Anclp5lm623o8yXL+er5INCiiykZ1PWu5YG5nBdHmgy
yVo8VEO9Pa0fErnV1SzREvlKSEjXD2fg8jPRjyDEdYTdtHMIWYQfqJ25QehqW4ZN
E0fNcDNhm+JNM+gXZ+5PhKg3+Vdt7pSsMJjlPCxrSpHMFZtzrsUdnkVok7a7ajGo
kygnjvrhDPa/ENDGhj3Yv8NzXtHS9SLHTS0gm4bcJSTo8PqM4NKDhaUhc/lLOMkR
5SiTFmxuSywwhFmglYMh0OFjGIY4vp+hpqMzpdkjEDQychsiO0qWxpGh/aRmrzaE
1VVl4ba8fLCmgBqcaZGI6rVEvHbGVW5MhZ4YUCBW24IkclxKbm6eD42LwnZzkugs
1ZznaBspdSbAyHedUqDmdCqIiNeCHjfvXl8hPuys23+shF1vwWmHTnCzudrXxBXF
Af5rYfu7839LkoVw+5o1QVbuHVmg8vye/+0E23is4yKovXr7AR2BHepAu2xFe9IT
fQEwOsu1qk4oDy7bNphjf/j2VpBIG6xwvnMMXN6q16xa1hXrsdmmpr3jzzjCP5Fg
cOPTciSRLprK1vNL1OYuceEnBCH9HWZhgTNyTJJ2RiNf/dlPH4349EUUJzQl/zju
+Wjws+cgcUW+x6KEuBWQALgFJysw75gL33zbvxY7U+Rhwm+F50GNr3ebkokxzVhb
ASTLZEoXt1aljDqZpRM7Ygl0AV/9DFJRcoMD+9SIectOEPjxUfPNo2u9xml3LKKT
pAwWXj0/EPHyy9chAWDexykBlbY7vEhvq1ZqXEO86wZA1ztMoImM/52BxbhH4ZoI
EUc+oRvv3BH4BkLHhtPckqiF/p8cv8pqqmr/U1tPUidS0VagH/Qnuz6AwgPAE2Y+
ioDp1TDAR/pZL/8o4s1N80NkWrWKUVArlZsUojXtAUfA1iG7bu/dBmBh0REjrze+
epSxKHhmjeUFPVo9lirs0A0fm0/yc5TtCOuypUXKWfyRvzHLiHOrMgJCQRasl+5s
eAX6QCCzGR16Lj+ry5wNK+2a7GedSZg4vGC875KTdrgFTA6o1C5CjGDa/3sQYKuu
GZ4INIm1giXlHG4rq7YG7gT4BK6ubHH+mnzozXCRTVK3dH2SlLh6Mcy0ADDGMMyl
LJtSrwHWcpa+1/53xN+yLTp104Y7mOxDAkDcQVBShUUdISAFQutVYF4a5cgIBnl+
uVhYguVU0+0C9XExYODKxIX6h2uNFz+KPVXg/vh0Yl88sNHhVRnen5YZWebvH5nL
IBRhTmWt8PtwMxter6loCA09FGzgvV9siIXFKjZs73eLxiFdX0p2LpSNmOfLeKW5
2pUKaE5Ihsvb79yM8Doe/KWWsvdQdJZNQyxQdFGrGTtPuOLwlXHDerEsvt4TlqNZ
Hfw78iMpm46uAAmV3slVI+sbzggyFSSpHK0Qm2xr7LXzMIjx1+n/Ap4OFd4B0auM
PHvddFaKTQ+ANBtR7HHlGRn4DB4dqBEQWG9AnIch2uOM6Yn95aQuj467RJcvo7/5
3xyX9KAn/x/TzA8euXPbYaYITc0M93w18B8W+huk8//WkfYGcABf3VbtoE8JQsJh
EJE/WM2TcqlE6CzgtLzzQBDqjGa2ux3Pvg9SFnMa/BjjXzh3k3zNnaj1pwMHmWMp
Dl91JQPp7ntCk3dXYVl3hid3EQ3IVTj0R0GvmA60QpI981UncHMOhs9EIYYSCE/C
9EyvRAKztg3ajHj+ty0vAoGkqxiPQAXIjpXKfeHVrmTsaktFDyrK76yc/1pqshzv
6+Qa4JoFJ5ESvzCcha2UP0zY8lTkcgnwKk6IpWD3bW0wFYBjOGCml1Cuh32z79hm
MOcPGYgANWsG45X3+IYWV+M+4AEe+rCEs5YQhjNVzxZooIWERSGLHvi5hgPquZ/U
zQveYE4t5O+9UhXBkKwGK6ukkbYcyA3cIaQq0/BtuvEp7HFf5cVrU0gM+8X0KsbB
2ncq9Bx6nPXCz+0yRPGZLx4Jp++5xekwrYHvK2d49pLpdNm57NfJ4ktgeEi883/4
ukBx4WymZAWnLi6Wp+RTOWmabanQeAaqayvjOBkiWIk5IsvurpmHPI+yK0+duOlN
w7HChmgoMdGhLZlhxuqe1U6E8T5iAM6uQkE7u3qVJ4+x4i30y/0tFNHDkvoaGNzR
5Kdqy77gn8ajFMCe+LsEEH3D136kxDYWUBZUJBxTlMD1p4fTemY5Ez+2LgHSS7eP
h+YAxFe1WGJkBKmPmBuGOuLy6JWDnu+QgIbDZmNGekSel6pKZtTOfFcc+ioHlOXo
3iRnhJxaUmY/PqocNe2dAsIJ6EeFKKSsPvCd/OGry78TjSMs51QhEIGiKJVrkj46
sK+y8gH8K0u3MiHacpDp7LZcEcw9dOYE4xvH2q+hPepID6on92nBlAQVx7IO4YYS
Vq9L13wVfPP3Z0FslbpVMgHziyPtmTA9to1OcRMnlnM8zdddwZtODI48JCaN+tfj
8a00jpauv38vWZS0fAEMXeA6iI1LJobMPQQB0vmU2xMYf8LKryVbHly5o7T+JEdC
WorPXmVLR01jQZ8jtMm8NlLHzncP5xsobFhFeB84/WvQK/G+tFB8DKr0oExa7iY8
E6Ss5Si//X9HeKAfKGxJ79f36wdq1LIq5EwjftXLKvliYoaSclsrSLZ0eU0bPp/i
YvWiw5GaisEOuLgRB1hUMi/UvXsULqmm3IyuWsIi64HPR+8pgso7zhtlD7okyaL8
tR0e0EQp0IV29R0eYv2A0Uul8v3JQr0LkO325NOlZo0pMd1x7C3jD7h+1/XFTe9+
H6VFPt7el7A7Mi6lpU+Tr9ofGQ0/T0PNluyC8wgGIBvNryhkfULusr3wk4SPJabX
6oIpxSaKf5VMT2ZybbJX6BLjxoRFiicjj7QPcmixTM9cjA+e6YORbIog1BfQ1XJm
91lzHh4W4whg83DhVopJRMHGJI1XllMbM4aWrqeJkFhrt5Up5e48e1BMPv0dKn2C
yV5+RIceObSOw+z36dgD12MfqhITPhpBrZaW8Tj+vKvNNAo8D8ELbk3Amt4Ifvj1
E3frbRG9cGSfW7oqCPR90SrAZcM571Vp+0pOgV1kzFiyt9s7zTDOu4oiIUCkomC+
KmzscjNL3NylwayVLVEeXezCDd6Uxf2hn/XE03WTHKDihpX4Nx1gXqlrCC80OZzM
q9tfCtpk4CAOI/HARnZvbJuVXqSVNMxKNxNU3q8nDBoNzaJcLglIHIdmiaSB++NV
ri2mokzW7EhLkhofOzLRtYm+68XVkHomqeQGeGWp3dVHDkPsbYEwttxo9IKAlEes
odltC/HF1lJqnFyDlQMZ45GSGUPpD48pOvwFwyNsC70g4TdDlf0z1mJ7UAk2Vh0b
JuF1r0aNgipWc2C/GVEOo25s/yTmha4VzMuWEK1ZAsNjY+fhMrorzOPp4eqc/3TQ
wLqAoC07LXqbDfxswqT/AoT8Lex1MrJHCpUzZafQtRkwnh+Skdx/o2w77amk+hDm
uRmRXTYGsFOC+XvZrqQLS4UdUjnJ+GFSpV+9n8BXiQwKauFqtmjQy3fC/whyMfbT
6j2yhPEaHt9kz6/IiKxPmaEe7/O2DG/9w7N4C+ZY5pSfpP4x3R2zgrQoO1sLMEp/
TxLgPOa7S3icqz4Hf99Zf9kpjI2KEOQze7vNogNkeKWcw0XGHyXXcQO2OwoTj2R2
Axlw6b/CWXiUfOx5FyCpqyBPUlAWXRgHRznrUELHF4oPFZZSyGDpyPC0t5zYCDpb
XBxyH6JGScdnaP5mwo0PrqN60Y2uT+l8ECeUtlrbL/SiOX+1BYAUEACFjyNqf/7g
QAvorZjZqvY1qo8tkmO6GOq9zQzCUvEO1UGRoLv9fvIrLepY46qyPHF5ipka0RvJ
IuDz7eZa5KngqEY98I+c1YRCc0K30JCMPNirLgrkbMog23Uc3wTgPnNnLgQCEJG6
VQkqhjtLyfF4AqJUtxZcfspMNZ0XDQIRtSIy+rpw3UzWcfye90NzEn1voFPXBCqu
36rT38L+aPp+lqKimD3VuWpl9XIVYBlb39H06WRRvm8KpCGduQlz6fKZik+/jggE
LVgNKJqBSKNf+6I/ie6N8U31gV928hxT8KgjIThdSfJfqD9HnES9hV9+Q3cvDf8s
acNRPJ4D1mP38VF42cQMfWPRNZujgo/YJ1ci4Tr+PvmE0mg97db9SxFoTkKerLY7
EjifvE8na7o9Nn7NL7XpAmFOPTvL2iuYhnKW4Bo9vpjeXPjADmFP6+0QHQYdVYHs
6Euui2oZR/TCs6/xUBvJsVkLwSlfYM9zk/Br5ZzHE+dB37NP4pCXIUwBfHeaiXhg
S9MdFlIjvuR2H4HL7FoBg/h3x2Av+66y0/T3K4JIfo451eX0pSe0n5LR1Nm9GBVR
6JCZhzYw/7j1MjV50vfav/8zsJdhU50ti6riBJkBn8gpewkc99lgfWD+EkgVS+3u
ZYfGkjeOtGu/RlqAfJZenfm2EuWDi3RKmY9+GebfIugYRtHciExeiDZrQBwYfJro
8x6asah9m1uQH1PfN1IeXTGeNEPtbjp8WrMTOt4e1QewbY35Nk+7YBNU8QZ0U6e3
PJXCpDc7ZBlYB9F8gTIsAlpJr6BeFXMQ05IQeHaXCK/8sCgrBtNzLsQzifGQGWi+
MIFwhe6Us04+9AWrwEsRJILHo+IDakkww0PcjL6dyUpctuO28tUD3RPKNUXTVzGc
70c0LQY+nOPxQJFjgZrXQYUoxTUnOyE9h3XY8TboRlNV+hZrGzyI/Grcn5pDZQOh
YSYU1E16+QZ3k1TJTrecV9HoT54yIF40H/HHf5fnQU1BSfa1ChgtnHJOXZQRbbfy
LfG1aMb2rVP4hCMERLRWFmpZDOWifFKW7C/seFAoJ4pAg3RdAjevaW6auq0zcZdE
NHGBgSqalcsUB/kMTNVvtm+UYnKBY9wXgHTVaicF7EIGzUwGCnJn2vLOFnVgdk4g
yvnO/E771SBuYWgyGIeSZBi0Pc0Kkz3qcs80W3msAJdw+KTyQ0nAcZJJflAjsrUq
JaYXPfZyicp0mVtAQuLC7ilRu32k0fmccFE8Jy65a1eMu8Vutw7OU6CH/jrXY0m6
H8Bn8YyRgaUKnJDTmsLEa3tVOsYWmgRsDuBTulJF9i+U5x1vJD3ak4v9NV1SXiUf
tjEymlxgeLgDrrtQu7cY+YIf5FYqhS5DR3gWK5bKR5IuvFSQkVHpezEudLxgfama
o3/A8dpvHuY/TMLnVfksxJI/HA46qQa620kAfQ5t5B5vJysDsEFUcpn6f23p8n8Q
5CRIKCJOZYPgbTkBZ3P8nb2B1keujAX+uBQP5GY5ENQxlQIUBuzvWN24kD+2SgN0
dawWYDv/xKpboq99tnAI5RknnJUbQuxNBsWpwfZT0/3L0X7Su0SY7j7anjn3/hs3
12L8PJ2C+l+i1tM1AWI8CiC4ZDIn7f2al/oIEDCeZ+S4WjulHR5hloTTrgnXcp7I
3SsXK/rFf3gTidj5t27sDuKectEzpxjQGvI+0Ozr95OynuZ3U+5btOLyxbU8nFp+
hhmZOfTDkqiu/VloQISfO/LHEyfWj0L1hVKDqeqprxC4k2j5rEVjARxt5du7vf8c
UxO9rmwzm/A+DYlEhyRZ1WG9BcUpVrZhanNCmgICVROYbzLxdTY4qFIwoWST0l1q
TdvR0QTrdODiND18DiIBlD7fdHdDbVUBepIiBZYI/kZPnCKDBvnWYBQLWj2LdDKG
tX342QMkAkIcmBq0R67RVXmm0c5pLAXahyDEuu8dXTBP332TFj+18F+Xt5EuNdz2
+QGoD8YaTCd4i96KHGWxgG3yxEIuYUGPi4DAQKPgff+Yg/AGqSxNh7ijywd5czn1
oPWjoRLTvwN1tV17sCogBC+VbsYMuAguKArToug6koNrVWUD0r9ELMcXFvfOsVLv
F+YOT5bbguDai9tZIgnJOw1adttQiuvj2xacMSXjhglQEgsqqXSQbCQ9/L/jnl/l
x4uE2OGLaUp9ixUNtwE/dELtw5AGRlqxeXlVPwLHmRAKAnnDWDRCAHJDjGIX4cXI
Qo08OQD4pwS3QGYp5N44OfD502VOW9TdSF6ePyDkMJAY5U5xLzxW53o9pBRfFqRs
jr8X9YGeIsOkd3znO3Csy9UkhrL7iQzxj4Ob9pHNYD4tlbwSWyO7zc2tqh6YPoIT
Y5w2k0AdxEpWY81axSB1qCkjK/cMnjGNtShDOsH9tIShlGhcXAyadkDdWNrNwS5o
wSarbxWd1Cg9NaQh253yAmYTedA/pV0QS6c8a7syjcTxC/lIEXLZN5mYMB6l7o5p
5QGWBXQdkhmWRnooNv2JNbhfCQr1QsFDBK6GEis/v09dNaGE1hhpvg5079di44yo
cIMo2mFeMq3j/NYPn7Avs+lwmgMcTSaK+VzBwMaLCfcRT5ISHNMyZTg/KJc8q/6w
1JZ14W1++BGNzWt/jj3VDQdXT5CgdSHDjXlWndwy2UWpDUg058edv+v06kf+cHcb
sfZK0x0zHLuHNPxFf4Q/YMs6mXgqWc9JBIp/oHih7KrR6SOPIE8EYfU6RuglFhLm
7zuyyVF8rYjGKf50W27GEgB5aAqmITloB3B12h4kcvTUD4pzFMg6SlrhCnLM42eJ
sS8ffgHctaicepygq+nkzMFcL/QS79VZt6a2Qy8covo8yegLBShZ84+4o3Qf1cgV
Scj/O6rHdIQn3IM73CjxQROm/YgeBmM41fXPS20BUI5C4lnpy4uQHxGDBgGKTeqH
rssVGUyvV5l8L5LNRI6KQGELKsLu/qiAfPIg9dEQPyp1Ss5pbLJdq40HFeHLpCUA
dvN5b6rqhOoc8pWnfTDRr1wuj6xNdhe5Sy5DpBQDtx8d/uphy+UdpT360cfMCSW7
tLk0bFd/YMqhulWijWFhLggrK0IHs7SIouon9TAiS9iuHrb9qUEnDarv1BJJvD1q
bl4gZa7pN62VAsd+8FGbJn6B6+GmIIlEtBiQznqc7iLe/PolDm1HWYwoEUOHNnlE
7s3GlNkPo8t0nHFiWNQgOP+8U5aQ9NUtAMV5n2N8s8wX5ye3tqSqjYfKjNDVdmOg
pYSU8wLHcn5nZVy/RS2pdvo3TN4RVoIfOue+uG4SeWOWotzlINEpTpqqvD9oLC6L
bFHLgTaNtGq7GAIKxOlysQdC/sXThIDsR2cVdaBC5U8W96rUUgcVby4mQZW2A7Jg
PF7TQ8xsvimrSJuRE3LAXWRR+dPXmDz4mb3Qt0z4/tHFqmeBx0IVw8+jgUbGU94m
D9e5VEkEGbbdHKD5onDHP+PxL7jKf5SiEN8diGZni9oRdDhrAiMFnZfr+Jo1RXnY
CUltII4nPdj6fd1vBUb2fW58SBwHAULHkNCnpRtn3DfV089od94OIGzW7IJxDR+D
6Xo1ROxJRVFS3wKtuxTfvZbqMkbEx7J72WDx5WQRyXXmXgmaD8Y0HUFl4RgH2TPF
Brruz5UTVT4XbGOzPiiXLF8VUJfG3mxsg/3UXnEK/PWXRluhnFSOI+X+mOi7RXd8
OhJsCFzhHg6K5Bgh59RHma+2iaJS+WI9xBEcke+2Bk0OrllriR9+yoVtjIm5fN2H
Em/3d0t7oO1lYbLcIdxJ9i0l3gbTVVlzvWLl61dmkMd3IkOzAD/gvXvUAV5SEecP
aX3eqBT7fRooiafX2TdPFN3BLD7rnpwxKesPWzttOH+sxwHKm9QzNPmjEq3j7Luq
CTfGEyl0ESwBRtIodwn9ikMD+91ijaCzqg/QEQ4HaC9VUKqyB4GRp5Z3n0R2Zm1b
pA4sjfEy0oCzXlcuEpBZ8Em3aW4ye+vYU97mICN0v4F+zgPpVV/yEMNTkTcnSTmy
GEYTGqdmWzZCDrG29e5qfQYiXDrVKYHcrcnkMV1tRcX2Sy/Xsn61bn/GEaemQlwA
PNp/xLfGPBTsD+e4Wzdu8BpSF8AmZ8u6WJGuaVZpUhvL2FuDcepngHFvR2hObLpO
SN/+/AylkeOZ/q/yam0cyVsQh/RybleG0wO0rka5aFsW83g7Sm+ZJ0CVrLGMmaFa
GupB/hRpenOLMmAPEloLp6ruZYfNuozt//91RsTMaYv2Qf1bvqfJi4K27IPqP31N
s0F2vY0CKkxhQ1/8k+mzMu5MejXS1ai1RG8GfKjbIrdHuF1YyP0xpp5pDLhiKxUe
4csEgfb86SWWaKXzXfT8mI5yvEqPDsCbLKCGSPKHfoSjRMuIaPNqetEbZThwHWnu
E9aWwkcmnllWJcnxXPtzYXJlo39Vwzc51nia1oPgra0u8DgrNYHHcbHic10W9/g9
1o3vhcf6Rh6Q/hnQX9G6IFExHeSFXvLDRMDl6Jz8gvHMBsbrlQ3YqTMQnDqycg6B
jXfGwUqhfMlcbWyYjos6A2dNsdNP6x7Sh5U9KNjY2c7nhdBB2ot5Cqdl1bqpCTvq
W5SMM0O1zy78RUqJhcE7XhJXNULoy2Z7g6iDYMkbNxr4bqvORmkDDYUqZUE932+0
GDJuaMB9GMaz3vQsMjuXncG5hv3bZsjbAlGhg+uGUqLOBG528nId+YPuCcWn379g
0lVc+DS0soZtkTEtfwO7LVN+nkGlQigxHFoGpcuuEUXh193FPn2FMiuZ6ED0L/QG
+6K0EEC/wnOGmH2kr+Q99ysl6B5KpsmLrZcbv9EFPKN3Z8S+VWmj8em0QJBrR7l5
9fpfabJOGgh0ggTbgLfL8s0dH5atE2d93qA1VCDDKVSBB/jDAMD8fWImqcC6gIVc
OJc50OsgV/dAh4JCpvdCZcX5LkC6x3bBJsWIfXQn0xcA9ZSgC/4AM2cd0OVSmQzf
QkpLJtAA8CkGwVKeyBp/crAQ/Y6Mw+Iv6i0qs4KO5TFbMSsCMIdBmmkkGh9c9u3x
M276WgQMCTsOrbV/ILD5BVNw2aauLb3BatnHZfOkBRwROfF/azjj9YZWURUQU19f
aM2btCLyC1x1UVUsLN7d1ndoFhCwprPOAONrvCbDirZYjmoDLtpIajH+itCFDb5/
d2RzAy/c7BmQujjxkULp8VljFGvFTcVGYmYTosxJ94/tv4KJyD7Q3z8Cv+EUhYwk
c5r2akwKEqznHrkvzPJJkZ9ODtq1n0xyCxoqFIsL9M7E8NH3G3MK2YRHZiuTvykE
MhKYFlVzS4eo7LsuC+GJ5viA6SRL+6SfcfdSkNeIxOi6+HbfcGKdCYWbrUfD5KMe
0X7PSAaHaq5HEUDAzVPA8Rx6KHPgbL7YiK6zzg2JURMoP/a80QPNXyBib25MLEY6
GgtYawbpwnfoS/P2Wc+BxGHxnxyWvYTdOQV2fC4vDDI0LIQWvptx5Hq7WvJtWDhU
vevRdvFbZywWVmF7f6WVJpWi4Y7oX1U9ViF2mcNN3R0gPpUBQL76/b2dOVF52flN
KpIgrUygUB6WsdR8lkeYLylH3Gr5+FQiW/xKGP1WxOj1ca9bfvr7sN951ScRbGf3
WJ6s7+o9I3Rngw1b9JkR2b7sdO9Pw8WyUxYK0RkOrhcnnVTeBXqWOxJsZWht8nlD
cOZXyi+vcrypT2YjlCn7BrpGL3flDhynPVII0t7RLOYrPIsXmqYUK83m645p90fw
Drjq5DD4N3CZV/jfhHxcAqwJ1La1Dk+eO+ClmxEIvkhBZBkuESYZso92PW7kDPk4
1IYMYvfqfTuGdb2zKEUo5ZXVA27B7TzExTD7aJsoBBb9UlLyLsg7gywOLfOf+s7u
rJ6acgLKckntlW72zTy/llt4aAo/r9/OXL9xMoPKJ3TVIHQzkXnbR6uDm6UsrzQG
5jqf0D5abS7nF2p+C8hI3WvhF398SqAoyqJ4UNi3hb1rU+8DUTRbTNk1C96WoEba
ubPwXj9E70ne4ndO6jMT6r7YWYFjRJcPrgTTlt+SzQfVj81aEkNZFgELpuie1gj8
OqrG+EbE1iNu9QjCpxXtiHmPqlnjC1oDHxJ9R5XiaXqxVOFQXvcqLSBUm+0M42f1
jJB1NOG/3brXr6YEWJdpMpRyqrMlZw8iKecAmdaroKQpnD+00Dom/MtvC5Socgzq
b7XHIyg/WNzapBQhWirQu4fOwbZM9PiIAX89KQCFB+BCzpQ8w0wLCvmBPyY6LHuy
agFoB28g8kFDKSs3sTLT/PGkpRAQsLezQVgDVjSsjz2d8cueeLXZNbDHGNu9IfQA
ikKz6XaRnDR7Jj/2ous+oUxjjhpZhL1ckEeRtD/uY1X7Udwqj6AwiIhO197QHUvE
Tg0s0itNn2vxam8V3Pvx0YrxotBjTmr1cak3kdtdxuPNKUeGaiD1MJQK8J05mjQj
qbtY7ZnnXYdhAkjxxQf0V5qhkOG8bV+eTIjBLFV0KlejIENu3h4hlAXvscNTbj8w
alg627mS+cg62tsNjWhgPcaj/ddkil2M62OyE1PsTC3gSfI+dadHTs0kvofBYj2a
L0Ma5mbdryx02d75wiTLIVzL4kzlNa4ee8a2sn7pmBYe4LR3XLZhdT3lBgN9BpZ/
itmxufP9YuXMuimRw9dPIQ3rz2DH1qEN6A3ozJKGgi5Ny9eoy/ukIDLsnGBKTCOl
7/LTK0KP8mL7gVmcGJ6bpnUPsKGhu9LB8sPzVsuVWsKi63gxV+/AMk58s8aplLTO
xktU3Vrkv+U8Po/U9PRIbUL/YUDQSgoabRM90LzLMxk2kML5lmDczqtVCVL1YZoC
+QoRxsvrt1+SDrxdeq9Dz4gmJ55tJL6ghgLZ+feYWWBG2bXQvBdO+MFx8lJmiD9r
toovU9fGGwsNSu6D0I0DsqSjbdDQFZo7/56D7hdEZ94Cfe3njFjWlEOteAscgiNe
8oz9odRDNNaloL9gs+KiD4zHbOSpaOoyZTumsNt4UYNLqpPWPsk8vlCcn+blA2ZE
y6hASwepuNin5T5JAN7xW+4tZ6qAqxHK7onG+gv0cnHc95OSfpFIfPYZhK3eQuVk
dgxBKn4CI48HZhlTwnyZIdbk6Ydl3YddMZAR81WvUQlrMWqZ5TmvySPjJkZw5OfS
78C7U+5PGiQOOQcnWXELtgctjSuXvO+SztOWEWU83KQKSPoesTFPVp7/lb4TffH/
Y1gLY4XcEOc4Mv18JFO4Z9gLjBEYhk49bWoVEu7NsnCtIox/6Oy1R2OrVPcdSqau
P0Ac4rD5jBomwhv25Mh5bSc86lm0V35yTs/4YtS0z5kZQggTt/kvI7sSrFurdydk
slYMnOP2H8sQZPG+jaXSEFI16s1SeI+HsSg5gZ+yhkGTnmzaj6z3+mxycJfE9oJC
PqROtaT/kdAL16PUrSCGBTBWL/zTppk4BYn2m0V4OtAPSm6FHb65DiI86IasFe07
FQIsy2lfpMdh+Zyadi3Tbbid0oXmEwH8RUAqUPU0QUHltIcQNBZlrZH+fQVcNmeK
zCcEh/t6rg/0BexB1fO0yOnC9FtcRQmYvVgd+uWsq9zPSOrBirCEqTYTuiu9aGeY
90xhs2bRk0i528wfUTtDzUtcQcvTNiRHE8jG89i6Mg5+5ySaoplHgHhX6T0l05D7
7a3eY8E/EOk94fZoRbgGsjRJqUQ6Ep2T3E5hlRcgFhxSEM2HflDuM5P0S+mkd5jq
LgNtFNDWVLq22lTHCLEnl8kTNK+2zPxi5P9DUGQ7h2UGiDtvDJPNc83TDNjxrhkb
4GjLCa3QwDqE3+1CE0yGWJ1+RIET1hm2KRdHEJ21Rv7kXMmVaHFfZ18RNvjqS0Zm
7kvfo6BLznYGf0Dtxgl02h3Nz6OwSZEex9bMkIdfpG+43r7GGPP+k5mC9sTW/Cp3
jUpSp8jtXTZbN+HivEkzdupb0PQxHUPsyxyqfHp9KYGtSVWCBAFtrmi4ZMLcLo72
uVL0iO86rMWdEwo4RD21wlmKYgbo5UQUywM5eMENSw9jZZK09B/rosslxxLDaF6z
2nPEn+jykcrj4154JIg0FAOvGjTJJ9LNMAYlAM5fe0PW+wOn8EF3cX9yEGVqH6Hs
iVTTGAbsce9VlcCCwsf4tXSfjd3HEzCgvxu7PTkJoRK/colnRelVOQx2y+Ltncwk
qrtRm7m6gdkOGYsd3orjMlxVcurHVLl0gpl2R/Z1jS4Nknjmrep+PrS43zZd1Vs8
C4NrPDUKmfF/OZVvfRedNM1aiX5sIqZwLzVf8+4ZbL/gSYBGRxQEhF95IcQ7lud5
oZpCozus2sogbr40xZsMpJOpJM41P0mAJQ5iB//lhLAt1fuizPNUEmS9ctjuXA4i
8lRtU5UYiaCZQqqWlZezmYgALodNf/7/mMGAqCeugR3DwoPeBKw02J9NTgieKlOw
O6gMJlHgvFceS5lforZww1d8q5PBsXJMEVDPP5G/Ho4HbGr6/vf1Y7L8fEAxfXLq
BTtUj8kH0ertLyULgwYSnTIHVVzG4XCSROSAT8faIwXelxvxx3gN3qjrR8v7oIzZ
+edB1KJCFvogRDyZ9rr3+WQtqTvZPRZ0tWQ/ShrAs3Q3xce3BtfhFSrFoyFunNtq
zdyf64YGntgh32hWc8XKzQsrBJwmE7KQ3d3uzpQ1ZHYPp0uJ6wKEikEXdqos9gCZ
wqWnhP3FsTxTWaBpASNSX3w+Rvti4t4tES6ff1dQ+r88l9ieda6miHbY2ABXPJ3/
IbGL+h0MHMm+O+jHRT8uCcKMA9ci1XSCrDS2QA5GEjE1lhVEpNbCl2cWNhwgJbG+
T2nWZgbP4oWgbcidwcYPxSfcOgl3/Z3gInwzw6ZeCk/XvFQLKHvVxLyldstwlsVi
giHcsZ+teNZMmjcC3WKMinkCM1NiAry4Wn4TpANyanLDu06NLTZvj7fWBel6iUFt
fGg5peadj4g4o+u1AI/0pmKgcHVsn44l2YDSy9kg2vdhfceB18zhYt4lDZQIUACa
TAfjBcPymBlOSNDrdVb5YMu40+AV/M2l48rc+5s0hKnk2VKoaPGiqMC3uF+3Nkuj
+/PYQt7p7z99GlWfj6Igncp2GvxGLJ5mzYrAX6Jn+CfT4MW/i07C8fVgCMWJRxb7
7qIspFh/HxiS1e1Hu/MVGiWChYOfGGmPumoujbRaFdbXc5UqWrNRPyUAh6tWRY6k
n4BxC4xUILkE0zzX6mYcDpUYSyjj4X45sJsdA56fCy0Ez4S7Dy3cNJ/rHOd7GTDt
GuAANn0QvBeAr1SaaJyEMND9c7VX98i9ZMV4kFxFq2EJ0aj2QvGslfUd6nAWU+ME
oekUu6+TWqq0s264/Pt/g4Wi9Xb0p8DtXrgtv9SGxo5xMVkg/b7T/Kik9H3ZAmlR
LElysvJoN4gupRxrp57oL5bPoaSE5RJ5nfStdkfBBNQ0ywhY2wnlnnE8XJWCMUM9
PofEkBJtY1q9aoc3AyuBROpjkkwRkyuoiDBOB//wTKqIZqtN7rvp1FhCh6MC4EEI
ySs+w93+S2Oq68jss9a7o1g/4o2JCABL2bbKcsy2slKUvRkv5vI0lG/LTmO2myMh
MkRmrGPUpoaL+KPeGD4qAX68Hz0ncMrU4Mn+b8IUht3pKd6r3DdBf4rODA7P22Fw
wGRLHl4gYdCZIIR/gcG83PJ8oXQVqGAyt9czD4o0lfbr5tTlKXRRE6qGX1EWA1QV
K3X6TkC+55WelxlPY7aTqHxDuhUukBiP8qBEJU/fW91DNsidcRL6OPZbSo/rnBDQ
Zx/gIuQKrCjh1C0boKc5E0YnkZzexgZ/kQydZ7g2p52xo+hFoq8MGvGWNEm7iNHt
0PC3lhC3CyIk+mx2Fu+tSYpfMxGyzSkPWM80tdKjf5ebIddDOQyldBe3SOW9FS6L
t4fzo8ceUW0vVSgvCkbpJ1jchSOVR8pl4p6Y9F5cmmwjQteRqyaWY/h7ix1gcjRi
gWlN9v+g/LGE2FyNRmrkijKF9IT2u6dcBqPdKENbjW3KQ30RMC4JDXLYUhoeX3VW
SvdPmLME/DRzLHnQCZCbcLSuufB2pJ3mRL5MRkxU2jrC0y+n/33O4LO1JzqWkG/v
LkTU7OkRi8oJ+EXVj+JGc5L0yDAbIY/cauaKrWhN8X0xk9QCv/5cYTGB60nty2TK
fO+yQSW8dxICFxAcOX1dTe1ZJDZ6wW9gnu8XH2sbJvkQlGhKdyJZFTMijKrhU6Vh
FlzTHl0+DAA9ITXg0nFH5/OkwnDVDc8mOJz/hPUW+g/vNAkVBzGR40ZhUurj5og4
+RsQOxs3jXNpTCC4x23QGUru9Zm67QWJ9AMtAde88SCFnzsTQbh6ZSFfvh0BeqKm
byo1m0cFoLJW2T3mTQ9+GxjRNWG2wq/qT5fMkdywlGLlJ0r+msUDXKyE+SmdhOyd
GH2vvCb+nRfirg+wdR5sn/0k3E2hj37bfVFfGnCMEuiELvGL516taB/N/G8gusRa
z6Tcx/47ChidSiiz0r7AnftAdfGrKmYJzBm1HDhYAREqXEW14wO1FIbhRi3VB8YU
pXnnxKTCoCMR+5eyGLJyKk36NAGF+xpXGHMLbpHGvU7kdZpt5CpkAvsgyTCk0haI
CnKftNvZX+TXWH1k01jBZzdNhTHwx3KAoCdPGhoBkwISiG9mR1iuTYnsRVK3hBII
V2Vtqg/UsDTwhQe4000IXBOJgnoAy291A5tkx5AQUPK5b+u/mNza/ZpEGKcHzrFL
iXzysMlTKAOqrDHisQoKwwoqhFZswrX+jer0t8BhoMhUezbtjPcg0CIA11e/VGL/
eXEAmniGHL/m4FRPDYcItzaXnby8tPG2n9DG3MZHDisgoBJTsMYcYX6o/YRtlo4B
Nq5D7e2DNFVUpt0ljY6RAXqVyC4gtW0dia99MgaAI8ei8NxrZ+dnoqkeLBr1kN1n
XJvEalwZFwIhkOiTzDuLQqBfwcR4Oppg2w6rYE1Y98AbAoJ6kkbwGivrjePLdeM3
4x7BUcpGsQDL9/GNCg9exuV97Yj1Bgu3+fDQmwQluBs8KwC2W0pqGSj+xPuLxXFX
4yrqHlDzrP70WbkiYXHgibwqql9fJx6f3dO7TlUMVtWAYTCZioKcyOZ1NcpCW8mA
Iu75Mw2i3/ajl3XOsBgsapWuY9uPSBAg3p9Xw0L7WZPheYO2W6to/3+cIBgk11jn
s6D3H4ovib4vND3qJ1yQjzpN4KxcUMXpV49k7v8WlWOKMYw9IxIKb+fNv+biPI7f
awWFnAdSMdTgfaxIs2h9ssZSQLxCRqCGa7HpvVae4rAP+RuxmQm4UeU6UM9G+XFs
g1uPCxd21yx39srzDVbYglLguncqUIwvAT5ekiQ9o+KpHhrpQGKFIrWhWt6N7lEU
e3ZhLK3mn00dfRlhwbAaY1S4Yw983U5T0+fipyUMA06J8XcJ7yFC/2nw9rEmgwtJ
VVwM868Woyd6VSnn5Q5uz+VL0gxPM4FtTyA33E/hdNaf6Q8/2sjtwL1OrIL8JznQ
jnhYaEoP0EiYUw84sF5ZjzxxprXJmtUXsW2FqDDCQFOBlcNsZmExrTvPOl1meeD1
/4sCgBLSclMR9aBAXlu9tQ4LX/O9DEeC9tsefmx0uUZ3ZH5OZR8V953G9FtDPh/q
jbw1fCf20tNZBpJerNhoD5hW3ovSYcHz5H2bJvGMbnlJMWgHLXA6kW79EU8VfJ0t
3VITjpGWiVv2N5o0jpQIEsf+pUTOhKIq0TIpJBft4atkfDABWVRi4MYxvKpAScCX
oLiVKDHxPVCL8dwbIBbGa5Qfk2HzOEVFyFj87u8tdx9w9kx30rTLb3c9wg7nTmBT
KiM6b6xcGwDvrzDYufRXXTjatjHBTg1Ixz7rjEGDT/JEzvQJAdFti3ylIUUKUwTJ
xpd4PPQLQokmmZ8Y4eH3Ziud1F9U5PwSI/IiNFbe7RO9gFeNzub7zazm5tS0bK+8
8fdmHMhYBhBRQibLdMFpKpdYM8xo0WVj5O5J1CBh4bZXgwsE19FUmeZ4Qq52WLZ4
7q83atUcVE41NQd8L21mELSNqfo+CZsN0CnDdWdT1+bM/9JfMM3vvxE2igCCO1hq
bzE6ZJ3B/w/rZjgYf3biyD2+q0He3c7zZAxIvjCkpcmdHjPr2AIohEGxaSc5n1u3
gYmUiWIDjnnaQSMPtipbgcj/32Eme/u2nqnY4k9FDHbMzDLJo0purHuFmKXQvanU
Y4GI4JZsfiTYxFtN7ahVLpZtCjXNV+cN0AoqaBwjPWSki637Fio9Vd1lBOgoWAMt
Cd2NN9YzLx+VajtyjBV2dQMVU+JoQ/pBHEkMp5ZrkrNnbjP3/CQmX8nDgT2zBr1O
z/BCk+pn7SkTsiwRYEv817JciZmzt3H/6GI1GVB0V/kHfptcwP6yXkc6oQTGj4oL
8h6TOAEdvvrb/tc1kQzfhQ4JelttQYhyEhxt6ksUhIvn2YOJe6oJL32VEa3W+xCv
yMlfl6+zkaiLMLSjjv8dFhmFa0MXAR2U2B8aIbR/jL5zdhfN0U6GUrN71nD131IV
xweVeBquh4rENviRttM8rOO3FBFvmHmdd1Bb1Ozd6nsFavQGDnvGIAx7nmDj3wOU
W3iN4CSKtAYdMJlU6iFzeq3D187TOoQHuYtDWuc9A5KsWlS5FUSrTVRF8gYVCzDq
8d0Xw391gq6kE7+zsk0hMldYXUDXZ8owOSYvOJvjF8oogZEADTUgdQJjkm2qrwuU
SvpkhLt1XjNKvP3GFiC+A1Ux3LW9B7Qf22uncQXXke7fY0rWuw5okXCdlaio01Ek
YEU1dHmsAtvZLQkYJFgJyxp2TbQ0NoA4yXdIUi9X8EiYxO81XDUAonW6ojaBGaYn
BLXLI3RKiSawew14QYHSHPQzxHtofWzxD19uKtBQ86RyN/vh1X5Bh4sjKCkllC+F
PNyixEdnOLV1vnhSLPQEbNIVQw6uzF3Jb7+6EYGqjRVACiIE2I8FgfzMFXlfJNpr
+X3r3OtL7vnKmhcOtBT3xRe/wxU4V8RXfyv0whkaSfOom60eKoaU56jit9IyrFlN
Nq4/bWJRj8H048u2MCExzIAAOC/9vw+QDyBzafu70zYVnrWi0EEGu42z4HBslIYN
hjh5ByyTdQofxH8q/2Ekri7XFl94b9YngY0d4jXv/yRq6yYnS5DNE6bD/r9Lsmj6
kFPMtdjmAkAWTdePCT5ZyQ9OSBpHfswlKE+JzVZ4cbiMNwIO8HaOA5TtJwViZPkA
8IEicqnoH86JYVwkVhyVFCnCkNA7/B63Eo5MhLcnl4CgxAVseoHNepEeN+MDycSI
LsTqwmK/bL5VMmCitLTkrqsb4+KPMvrAa/pvc7e673IcMLk5m6+LuvbSnpuNcKd8
nFVBNcj3KRDaG6GzXTakzMDd/2KahvLlurbgPbhYvQN0BEThwhzmPM5fMz78IDvT
1PzlG/1bv5FRWaMv70K3A78vqg0kjCyk2eP1GemOBZsTd7vdKVuRMso3iDeB6LF6
JqAhjPvzZlVJT3H4Xc4gffB6BMWCkLvYs9qf8KU+u0pmDD2M1veSrN0iFef3Pk9k
J6naUwPNZ5azu7h6JBJSQuG4wW5EY0pINApkje7+1AUPRcq+Wg0oku7CgiE8hdMf
5MFHsNIhz0jdWTRjCvtm6fXouZ/AwwC+s7+wDLuyc/iKhQVmJiVL3qPZJCM2lm7m
ao7rNlJX5D7aagf5JCjyF2aRJGZNGx83FfuY32KcZ8AAOXDdCHMSDzjWlFfc9c22
8jWbrD3j4dZDZVT3PFNLcS80qZTMMHcqATjeiXVfSfyBuze+zXsiRizj/vPe78/8
wWCBXuFZz4tc4WWCacvCQfGaOnIvS7PcPCy+J2GAk/VumXWGR2IHcJ90vvxdcliw
vpWfMRwRz2urpY/N0RGN+KTCCw1gOlp9rr4muzL/v7wbynZ+DD5qZbyS8cWKLKZP
/2PSwAyk0C820Z+x52GarUGMRH+D+wl6ILRg6BjzgL2guqeDiTNJHalWzKCZrNLP
oeeFFd2YWyWNoWDCpDHyhbIfCJmiHp155gZsJKb+S7yTjcrtAOXlSoC63MDEV+JX
/2VkqXmH/dAoNf1sfWKEikYflBQLVhF5nlNlfGRDR5YMtt2kBIqyTsO629tGQYqN
LjmWzpIXaoZeykgIjN/qhMfbqv8nxwq7a3vQw0vB68rY3xf2S9JofzAbqB89b92i
fXO9f7IatV6VigKNYBneaiaTTW79f/D4mdFotZoMYd36o3qzWT6sfu+9qn17U/m7
sNpCtqwSlwB3WYFd1FNXdQs7TEuuHbNA2WTeYTb4+9qF7TGZKNzugirjrQrrcAB7
MwXijKWRu9UQIBm6tISbF8Cu9/Mta/q3xr221xR6fMSDRCyx7hlySLJ8Wm4Q6BFl
tbyDTUm8sKzRmWzhEgNG46Z/oYisUDovCKnK3eKhIQV/M/1sJ8Ag1Y2wZgZpG8fw
nZsXX5t0adGCfu2KsDE4PH3vKHsr0NEZPBYicFG7LUSgKJV+jfpcb91dmGhpg+tl
ezbjX86XzQktJMbIpet8Komz+g7ELvoejXOvPXCDDkidLJyKjJpCulo7TNClNp1c
we2TNm/t7NoFZTgiEIUmjlpM8vYthqkSbdTMSsFcQwoqBmkUuvAgDt7IT7bRO7UV
rCeVFyRXQSRLeuaXutOY9WJksOARp8IzdP/V67RPt7pN+R2yipAE1FoyKlh7nzJU
GRTDZVmTDlXR2RwfVarULkzhrEUO9br+JFoK3G7WyrC7nM37OI21M8wRtHKgf22k
Xb/UW98lc37mmbxqENKHodWa3ttgRF+Mshij1z9UZqP13rgTGRO/YN+rWBOGZcUF
Pj1cJhKcCxWs7jv8MR5mhRKUsX4AMSXI707ZprfhZx75zSimqWMbDwr+sC5kBQlN
51FQcvvhVD2Un4xvBBCET6KgPN12mgEjueyylT5ILQmhFlIi4ConDXaRD8T/ViwA
VVJdUBgWxFqQgYSaUR+iBqEpoNo9y0qDvUukXrIxge7wU2H1MyUlQ+KmJGFf1J3B
uOECLSXBa/6HkuIg5wM9WupGcEIrwPK40UurnPm5WPTFy+x2lG9LMHGHZz8VcDVz
E+7x1O90YaJUZWgtfQDe2XyA12kMGic2vI1wL/eOgUCoS1TCksJzW8o8d/5mI7uC
JbCeeDz0axM/9CAlcqEQfrVnCRNysyG1AM8jzar+UwTWPavoQqMmjd8spR8e0sd3
YplPqHOJeRRpLOl7WYHtpJ0rDfNE5aL2Zp+cQuEgRXm2qjBosDgvQmL/ikIGOBuv
a8Hi2cvQffpE67/hfhFlIiabb8FmtileBsbxEQd6Fm7+lkh9TfaOttRoMfBQkXHc
JTI5LYowL/MT79W18ZWeB2tVFYMmP7mgKQvYJFhPGbsRKfn3q9n/xcZBGjztQ0Hy
kkvz2u9UCb80SWCIqmTlo7qDbiwvegQ2OkQkCWS/JZ2Jh45rqJoSP1/jQOEjnO9Q
jCHfITM9c5b6F6QUO/yjDOHPxPiCQCOs4Br3J+5z9fMFJMbl0bfImgQ3gKAdZ58j
jcT4gnqYvxfNWP63tnjtAKlUcChGDHz2i1o9E/92UQw1BasY96psAcE7LanhbJ36
c90F9BYYsYbhZalXReZ7lJtpfUavN2vQmb+ilRaViq4TrbFpSAwJdkmCgoPdEgQ3
fMiEdr8o6spFYcBCys1/XGdl63jpDMk9UYqcTl6272vURZUxdqoB6ZHQ0ZryHLXr
3J72RQhj+uHpQq1/IZ0O+h0kjHND/j5BBfRcXgvT6JBXw3WMzKsHDLKb7wW8QB+1
ui+gahH6FWPH9l5T9GwcKUis34p7Qgz9nPb2tT0SefJbHImo0zM93yxbA8YjFKqP
5gxKMMRDYjmx2Q0QZeO4ozhRi7S5lW9dvMFb6g7xvsgwxU8JnCc9k0X2RCJs66/r
mtehIpHgc2gnu0I00jiTE2Rc6iGC2j6aWfTxoKvP7i8SbdHDwXOgrvHep36jVdp3
kiDouB+bubh24oK9rgwSYAIR/pQxc7fhYmp+TxRZ9zG6u2HYD6apEkDRbBVGGmp8
7aiEz/ZPO/EhpkVdZ3a2AwHgEIlI7ZO5oKQIyNhWRYWip6e4nn5Oop+oTP/U11vo
L3sL6gEcuwSYMdGP2Kf5Qul8xkiVFavG32KwpgwOh/dz6J7ehx3hQMnLA7eMfc+H
GXf82aDl+4xv7tUWJsvjGejxe2xY+LMvIliUkMia9EM/nhY2C0lKaB6ms/zs6ZiI
k4YjDMqtUPTtA0J88n76ks2wl0ymCR5Kv4AD3m0ON/0Ffanc8vr5Eh+dHv+NaAXs
WJCVHEBZCH0sFJVULQz39OT8HOIWm30C3DYsLe/aVmGahsiRAHetNeERHVLdJjj4
CkZwvOXgXHhImY7un7seEjaiQ0ixwvTVndIznNEibyCDC9CA+UnCA83xhDCzMQ2N
d1ZKfbgsL25IPeR/50RUtJOCvG9vnyWHiLok1qV21s0wfRf3KVGYp4Gxa83cglSI
lNS0tsAUTfJhDkPGCycsum9bJpDdhQxVcK8WiCAvXU24QYSkIZZ80mwmNhoeK/f3
twOCk66JFQIPq3lb28Xjz9lBzesL8UtU0SvbQADU3sRAJX+5sGgaM26+3/4H1wgm
yYTByG52BvXx4MwunxywWq9QNbLspZ3ytrr8FE6RVmphRL/nDqXBEex4oP/bnw+m
vppcHaZtRZCFkjA9y608d8r3yJVpPXeTXAnHBAoeFOi1P08gy7N1qjkqUauoYmrd
Qw9b0tz4Md8bCONOJueEZ0ZevfTHCR1vqioQi91gnnr0rWEbjoZJakQ5ySjorjiC
/c1eRe0LvM62YCAbmFRkKPWEeeU7jGdtmEkVAfxQKlMAfqlhoNVqLU0WGraiRyB6
jd6RXtosp8B+g2UrpVaakSS0R2dXU8HVToctawtgQ67krQTAL1FyXi4PywWrURYj
WHQnNFWImSxuaEe4uNlAuBx8gQbNyw/SmvKbhPDP9+XRCMoPxNitn/faYTn5A0Oc
6XzPqU442ZoS43OBrzGPtIx2IkzB+ni6XY6RZCtuPblZtKwDZkjNQPzQ7RXW62Wc
3acvua+LjGBdL2JFICib+QYeV+Z2eCqSzehxqjmqzaVVp25YAcgvD9anGpkLaORz
l80jeQVTMCf9rKbI0Kp4Sg0Kxbyws0h+aIp6CJUnx1DDLD6r1A6WVXSyASkx5AyW
U1MIQ7Xh0550COSnfTdSqwRbMZPMwYCsmpa2fWCUykISjYyt/UG78iQShfg91kKw
vrqIAbOtPm7Jxnj4eGRmEQZMC2uHmphNceIohrGu8ltOmDXSyBRSt7GWbg3buE9h
7iQ2LTfr41ntEPfnQgzrzQrUd2tQMbGvR5ovCXuVG4GHPEEVbo/pkN/s3m9ThI97
EsN2ag7rwA/hxLb9Ub0QaP1oXinIQuhPVfHGD28zWJrr2sAV/30XvcBZnuo5MYSg
7lAV+ePZAZnLTlxvnCryHzm0rgtYvQM/4DAwEvVrotVTuQ4fKrwIJGxMHvHrbsfs
571pwoqzO6PEqz24xnKC3vYbx6yx3c6oBLMkyAl+JBhVISIdyXtBJW7raQGVqq5T
jGRwyqJ5DwOsVo0feOPxPWx6iXVLwv0YagJUd5GPAmaip2hVmIbijlI9m9lGp5pp
kYSxUN8cI96hdXPLmkpiw9XFGtqvZ1nKNt4T0X1/ALk6dZZuaseQkJUUlJp80TGT
mE106fv8EAfom+NAvW7LzfTAquihCPjUdeD5mu2KQW1CEOGZOeP9oqKFX4uyiVzH
+rVM7D7qCo5LyfATX9VDjy+SrhKcIpoAS41w9TlCvSbwdhckKn7VSHJMqxCFNW04
IxXK7gTTpT/6UcqDLuJwgZ3ZqLP/lHYWvkZqhkO7s5qiNqiwa/MwucwjCYFibCaM
otbY7rLTKaS4us4Rte2zzpTfiMKj9MKrRm2b3wzUW9OHei/+rsrAx3ryoxFlwV7/
N8cjasmYKwMCdOtTonXWf+B8LrkHNk4V2S/LfhSvQCO+m7mSYTGP593zcXQVwlsz
fwyP2BPzb2HICwYyMxKLnVJEYLaGF0wyLvTcRMsJUWDxr6mSGFvUqeeo4qIGzuQ0
XgbVIEcv37WW+gYY/jdB4jWuOXhyOAcbEM9lwomlHsc7Pq/5GK0neXXC8iy/tFNn
PaRCXGwWMaLJL7f22k/MyyKtRedUnTTQLAkJeZt+DHLYKzsy9e3nwj+4WFZmoLRI
Nbyc2G6S+4iGGhENTnr5FylS3y04C0ApKCVM3wb/QObIOfnshvJ0aEta8oT3To4M
nt1q+HW2Y+scjmDa0G41ZWMv2pDgxvbvzNoPre9H3cqvyaQ/Rj37jYUXWPQ7ASpL
d3ARcA9m4fn02R2M7uQQm9/oaKAoNgCmY/RBpKokFq1SQ9CQ0Z+JAO4zEtfIJGWC
pR68j95UNeYmZuoAz5X6HqIMMosMWCXh3QKBjp9Jmd68bJs0BT5yOnWudbNjSyCL
zyQNDUhdPq9qiyihfq5zi3EojpXseK0lSJLPQOpdPhG+37Zfs//eUEzn9EYL6V4r
eXaErOESt+XKobCAw6GPCFaRGVt3B6+kTl4sAMoJuHT9efwSdw+5ctkNJTerAau/
oPob9ZLK1JVjqAEgLCkJJ1VXmYMXnvubE7DqhD0d1eJ/YSBjG3p7FlsOroh5HuLx
ZIjRmHgnu6Qw1RpZG9tnCx2DzL4+JV89A+dbR0sglm8QeJdVjCPro9z4SP4r1pQW
CW/GYOFBoX6CeMoRmZiQgAOs/vujL4imnsJbQUKq4XB5iAYpF0HREhcxX+Lqh1Q8
msBxEGsby5m5ZjCK/mp8+5zIiW+KsT+/5O+ujpzupgJL3xbDowunufrSN+WX3dsA
rPBh0iXs9tdLINraKa78KRWYzn8bFnNnZufGJUzZHB2Xdny/xoSi9RXN/szklLZ8
my1z+WdGYzo5LwMzZ3uT02FJa7+5d40bhmyVcj7arpBHGgRSQKdkwkWbS91SHRGc
YJ4+w3cv8ESUFirczJfTWHxOMekxH994M7GulKsuxd5nrPE2u63pgzqcobB4xYsc
1Y/mAmFLhjtR6ylb81pu+2m+gpU5Vxgm0n/zQ0enzefce0Vo4U/bsBPYQJsDgv0t
GsFcUo/sk7gpCPokEjwFcmevvAWYYGqfCIzENEfUltWFQe4fUNKJb86lBMvz9sWj
gJRuTPne2zNSZqRil33FpMOu0RgkTFT2chLJnrfJDDs0yDSLzByd/ebmvP/xBkiL
cVs2RS/uisxBRZlUtjSxLGWeCU8rlQxgj1mtbVfO65/mv59irVLN5B/ND4WnbMLQ
Km3a8vTbN6lm175puJKZ0yR3YFbw3cl/rwSd5guXTtE+HC2ulSo1nRyFC+WUv65P
J2T/Zzis+o/OeXszYmB0X2IqHVkJUdk425rrphGZ3tU66vQueWprJeHTIwC2SrH8
HFAUBZkWMhc6q33T7HkO9ppe+E1WbCUMJwWVEymXd+UXPCZkRaT/CfFWomRsAXxb
Q5398Mv8+8qUCzexHZiwfsvoB8Sdodgas6mWg6ZPhHezwAsYS6m4vY4QaSTOliYx
D8XEPw6ql80uavrB4voOVco2pL3VfNINtE3D7DYPDID/56izpkICfs+r7jCQsoxs
lVRKr7cAL6IcqBwyIquOHltd8LJSnuTCUxTLlY6PuS+CCyYeJ3FEYI7kTcuyzh46
rERL1UPLgHYKls8LQQyG618rUAKcahSTF5E1AX4BOg7sEgx099kd1hLTYQxnvFto
sQiVZnHfcvqPQSUWGhlymXX4w7rKSjYtkw5FYCaGPQixLwp7Z10/WdfEo3cYOdSy
qP/ZWWRLVKlLErNifov/yJqgYuX+wfiYgKW7iZPr9s1ksDCvTtvxNIVkyiF9sNIY
sdiQ3ly3ccQvxAic2awtcAtu+Klai5iN8Uzqxft2NsBpE0eOG795oS0bb1ouJfB0
COCk+kmCMWblmzE5h3sWeK1NCnGdUSrXo5AHHBQL+fGddWyzXkqYVW4wvBStalop
LqtI4Y8fniMu+0SdzJQeFqHfnfesK8r1fHkyxpRBRA4bp6uRQe6lL3GRqlIB2rKl
gBG/hAjo47i8GJqVVLJ3hyNenB8NaXtrO964SVsfPl85BSCuDsEnm9duGD0wfus4
XKny2e7sgS+Ao3eNU1b7dgaXegcscX8mGNTdYPXNrgxwo4KXMP2+0MlPOFtj/T/Q
FvaGIN+XI0KWt5MMc7RiVvAeKw5u2cG1K3z9m/2yPnDy0TrgxUYWbPLqpzv+9enU
OlVBzA/bPE29v9/MJCQTQRwE/6bNr8Ldyx4KEqv8LZy1YXfNIZPAftl3Vf3U3NkS
j3Ll0BpbIko5hQhB8FTqDui0ilG/zAGGh6dQFSwcoKpE3TElkp2Ts1cSvlOo42P8
0yZ7XdnMTer+7Lfql37SqwBAJDQGGUPqDNZ1KrH0SB6p5lC/R5EdJEpR4QrbtpcB
2a1zHFuSGwlwSpmXBTj6ilHpTHGMm1H+xjKfUBKwqFldUpuUQcqwNESTzeJNYsle
X7+3uHZdvSU1Qr3/GrHyvRMoW6CC6v9MmBtbhNLCAC16DxbZ2Ztqyg48dBiWutdc
7u1KyJpKeuiO9mSCqs7eiemnV/B9965tKyCB686HgYUqswjfs+Gq2Yl1uRjBu90n
4cE/pMdgxlVHBTZxAWiUjvslDe2eqf6VHZ5bGmwTVsOf8xVhQhxKXtZ4gN3Y9V9g
evZgDDNskqwhIn0fEcTga4Fp85+UnQHUEYIJVulPCuyJW70sO57y/7zwaSuOZBxi
FDZZfa9+10m5dNSmAVmTGf2z9k3Fgj5uOLMp6pqLt3Y0xhTIepcPT1oYKgS3VeL5
r4xjuqROOlliZ7Uq+62wOo9MjmPGcRxPWEc6u9YmM5zzEthG5jk0WzdHaL0rNnbn
lquJQdZE38qOpE+TM50YXEmbt/+aYuKFYy2jK67tOpM+yXl3YG1cKHyQGMe7Q/sF
2cTFXtu/TWBUx8T+ajQS7OSBGNaQ9n31hQBcb2/uebwMx04QLa/EjlFR/scSf+0t
nmRAQPlDSXVwIuyt05uR7bk7TAPlwikpF6Oxccjgnaq7iojF2potimL4qOXwJqOH
QNzHpT8R+f/Tr9n+/MkzdBwVFi8QwB+k3MujSPVf8jTOXEDe9zfq0VlxKLGxKh+H
w3lmEGNkQsq2SbUkQXw7gMpnTqxP518OZWSfVZUwpViFWB6hg8CGJBAdaORkzw7F
wJB2GMOPYKsCcFsCur7gtgd2Pa81rh5CCQ9mpdufkZbH+f6lXUdPYPTIEhYyUgNr
sbdVzePmBqOYHDH2vmcyiY4NhF7wTynQ47XgD0BZgZhhnOMNnl6HoJdKQ39DB8NV
jeQLxWsWCAcnR+HUBmdtLIhnsNGqFL+KZmqC8uvI9BuZv7oNW9lG8x5BO3XpRRvF
876Fzxs/na3MovuR9g7srEH3kUhyNBuc9OsF2AZAvb4ILrivPAcjqC8GInPuM8mz
z5PbUikEvGFvdkGFqvqTBOIzqHLg/UCu1eVhwmOSvPOm2Bwi2En1aGMi6umv9Gfl
cd1W5oEuuCUcIzWdtCkXazo0D3cD/Q55cJDvBTm6k3Lb5Uj3eSjuCoxODcfoKuTJ
CF1McmHKWcICE5uYH8UV7Amr3vz4gEyrW55WjZ5zjVIP97AmdISWFD2zyrHx/QWP
mViHsWO5Vn1iOLeYxwuFVyj9EM8aAT12MTKbPhIBhhAML8ZIpxwEpATjCg1agrtf
YqbSnbLejn/9oeTK8gXGthY4ZurEgECw/RNOIze3kxPWlCYy0ICNC61B6yCCEAMf
ypkMS1Scpa5CNcLBHS9SX8IWwd0nBdevBzwcROociWeNAGodVQsjwqMBiln8afBv
yLiXgMkhtf6T6lmJEefekgdd4cyEioFk8vVORO6Jz2kaJ4ijJp5dF6urU6L99ryK
nZVVXr6kGjGowYzfc4if94NcqNgopyrSssqrYQwqvOM6ujKFb8Iq4MGkG7jFhV6V
xLTicRPNphwJBaLjkSawkpSTWuR86rSfuNPOaMQGvqedcB44hru398EbmjJJrNv4
SaOx4htwH/q2yrRXJB4XSYYnIgHU5UQnB7vwPk0gBdWa8/8LxDbhDCj/gWfQZIBp
tFpeEsVJCKWhUBZ6dEZ3Dz60PhqpTXuEHi60rM3gU3mGKbIrlFhAoSKMf0jcQEEy
mkR0hNnmcf8sjir5Ixg0DkUd/dlGQTlfnU/QuyKcfXvxPxQyqbRkXrAyjRa8UK4y
7V3l5mlAXXefzCyHLAtjM+ypXbABMV4PY/dueuxvs0iTkhsGZSVCJIyJ162pXnuH
3zeFmJMK0w3g0Prm/U9EzSf5Eke1INSVyzsJN2y2eG/qwBK8SICxFAnIGkMJvIg8
7SHq3pGWnCBpjH94m4kxVm9GcQgjquah2K9LB977hsgP/WVPefa7zkY/e51heIVR
Sxyei7FR2Ch2I3+vOOLJZThtU8HorUbl8QEhFMYMU7NTNGcP//TKJLcLLqcP0+dg
yyrgB1OSsbVXz85rjWnOc0IZOSbXdYJfHyTzMV33rLC7NCU0avaqK7RgA4cha5Ks
+0DQi+cUIUW/sGLCsTOHAEEKCmYWDj3wVhn9oB2IVBybe0mrJbMyHQPkDgwabHSR
uG3d4EGJgXlylWeC1WatB1BuvGMaNP+IJ5SQxKBxZ4GgLZrqBXH5/lyLzX/lEmJ1
l+gVvRkaVx28vBuLuJNB+IQzKn6D/VCx0Lb5K7iNX+J5+ZHjX+m3rc6dlrN+hZ7q
beErVLexQFPPx3r/yTxvHjlay87PwNaFytFGSwSuV48EOSnUnqRbwksSt55qtIYi
i3nKHk0cpsBDFTx0oGBWeW2nRTPGCjxowBgT03zfLO+LHWtv68+dT87ul6wKZus7
uIO13fNW+lEYytjikVJsqfm6dkIYVMKDHhYcbMF8XfFE321gsepBCD5masE1ACeD
imXq2gmpUVupmUnID/sYZ5ls6lhndt1wqXh9l77h6ZczJmQLADpE39F4mYVGSo9L
iyGgwUGIYsMUDDOVPljinwNQlN7iQpldZHtHPOJCZ7cuJ7tVgDNV8t8ALGt1ygQc
Wp8YWlseIOYhC4nypnvyyuWU5Pg6diiM/7ugBRIMZuh5xyB43gkrJbkfmnNxtRbW
YtEcLKKFMX2+4L5vNF+K/Ci7xqJapenYG2T+HlJgixKOpmrDs5c54xfn+bYLnBpv
4hh8zeFpNAkyP4CBYpceBKXLCdDnvOl250yTHTRbAX4tNlXxZJltz8yFjTmm0alP
YeAABxXs94IqP/I9YK0P0rY/TY6/qVsP/VoFbRAQNaUdZE5PDQ58VrC3ssjHnOPT
mHINbtsFPiJ0/2Th4JQm4HYP0a7Eix9UJwPfhzQ78z7p/l/ZNYvLh7Lmw56fw5dd
2nvOWjE1hcMpKJcX7gK01l2SkiNlazsPAmj7eAkYq6k3fjZz6nQTnowitg/Tmj5a
CveUqenf5JC4awAfhbCNrqlj0wBPv+JUu2bUoAo7joZWigcUuDt4iM3U5W2QnXwT
mB3fDOKAaslUT5QISQ3oL0ylGfinmsdeaHYwxhtFadKvwCJWxtDVzQkHebESYfSo
7a6F+SwPaT3yRUDXmTxh6NY/deqnE00zENqGmnPEP1ukfVz/fNt7SBzme58sGv7b
te4qrzeNcF7WlmuL1IsZ0flF/pa1PBlM8R5L28tgWDXETMhhACOV7vUQb9Dutd/8
S4Dd1JuYceJhf1M6YLtWai2vOo4QBLz5Q4HC95gvrZ0PFQG4NPaD8YpoEcO5Ip6a
lCb2ECIhyv8IXScBaqohzqWLFJGUCCd6GBw5oF3bFak6bLNjs+Q8TNSy/tgtL1Rm
GYs4iV94yLvpX185FdcyIhWQ5bPhvyoh6+d+peH1+M9YiU7dw1lipkYyDWbJ8g+O
mHKY5N4qZ5KQFNhuclwbv2EEM9x+3T13S3C2BsG8CKBc2SuwGeiyneVZQK8PSGSy
bBCBAPIjhdUppfzWv0si6WosC0pI2ucwn4nHcwbo96LNGjGGlbpdOS5bQo2vj2IX
efqvj17yK540jRBJ8YIxeOUEuX/XrcuA9aDhQy+FYdHavIoCc+HQwP4qWNJboDqj
JCdp++KZQ5//6V83dhnwTjUV6ErtCII92zdaB/pOzwZ/dikZEFQ6T+DdFzp1YqOs
XUkGOouilSKcENxZ70e5dZOp7DUGa3553qvCcTe3RCfIlRl+7CEMKXogYRutMfJH
kA9J9QK97Zh3PDoiuA2CJ1RDFCP2vjZPQAX0bk/RGtO2S274fxhpP1JXG++YWeU9
WQMgEzCMdpHeKWneJ8Z/zVJwfIXdt/A0VYfh4boCWTh0bSPL273X2fkCvfOCrxr9
lrsZMit0k9/YwpfBtn2uR2CmrmegYGw9nFxdqedtfySwINIe9NP1WFW7IcPPTeTK
z7zlH/y72PfT3L3N8hiWXctfD4RekVw0ac6mpu2U9SuSgSS9CAm33pTO4O0CbuvY
2gfKqis9V8VG1wZa+goEuoipO5SpTvx2UTy3SLwydtIj17z90OpfMXZihi6RrAN6
FSiPf96urJR98cvlNA6EfSKQZVFefDVrbc16jyf86BRaJoXoBJV1xb6VWzDiVqKp
KnZDqkrE7nkukGURpRHtDQmfBA389zGfgaMmpNqup8ernx0+LtFp9uyc0Qyc8SzX
jq2WiA1QM23WitglsZLm7XucnvNFcT8rz98VAWFKWU10ZGvI038JkS9yTPGnJ+3t
oH45u6ijWZho3QIfnoWRSDOiY7xhPdFmLkPFjNAEFKzmKfFdrjHyWI/i6InmiHOL
DcmndPHTjdyfXVAzb2bAwiyT1wN61E5+2cumIYjgjdKQa+S3P+yruUVfTXKuoQ4h
6G5qVtJJ5VwZGdWaesvPymtGNwsWoVVRhLXimlJbIuVP9tKhwZqua6rkv0Cekj+s
mmYzjiliarPHbwK/6Xhihclc+7UAccOc06faVC0RPRUe/B9LGHpk8pKAhA/+zkhX
H0+xRhqFNn3hn9JqIsBvV3YfK/wt+xtPIz4cFaqaYZ3s4FgBjGZx+7v5ELRW56mg
veNms4rHXcCpSwEgD7Zr/YZTRvaY8DL4UiaDGpQWRvqXMEHz3LSy2ex+nvrKyo83
n+52SH17Dy++KiQM1yHMctGcaxGV30/waQWPRuvRAFUWCC1BGYIsDTWg4qt+lnU8
CWb0X7azWCwoYOd00O4eqDqW6saRnU8UyQcpJmNocl5N8PUER+t7rg1ZafRxv4fi
lgyCzLqQPwc1jnPhCd1/tNA3xFYwmXTkbW+1/LIwGzJIFaokist0HIxqVpfB8Y9B
ve9X11xfyAInQ8Lmrvr3hYtoksYqpkxZYLBkDibsAmyjwntl+40gdiKrDKMDTCqF
mLVx+tILV+Itvbn68Mtnewkwy78S3YNuWlg1laSaW4fUeM3TW8cuyb//EJF/Mzbp
Pg3AmN1315i1OxEInGol9qbg7tPgeUwjfG8wO3dpJf4q0oRjt5ucHviqifikxtaa
2mTK+t9sMR6fglv/KU91kMYjRwe4Sttav1fZLOQnerDm6OgCkrgp3Jun7kZohTbu
waIkpRiwXnAu9dyE1z1+Vp/vzBvsvLTCZR3vFWV/ZJylBdHNMqxIJG6Xw/m4R+4F
DdK33+0XT+wB0BQEXjhkiY9k8X8LZDUe9psSN7tHs9FEze1yC6usiY/ly1TM+O9/
mStn+wuH4j9YFdQe93pEE5/h3iCAp1QoJE0sR+F0TTDo+kUU/Hhx0OJTzHx5YPK7
8wBN4eaqKwsbu95R4Ggm1J/Vvw4ZcIsoMO5fLjTa60T6D8uNMzwMFW0JzeMXOckS
p8CGHvVEapxDt4tNIZBJ9BGHnlBSGo8biMjCOhcdmUs8FiEiwCsE+vgxijikiwXn
20Lsk4V6IGUQ7OJVNWo9bW6BTWoGHOUWs3FtjXWQ0g/3n5fzgMhdTZnLDVD9cFBG
EIwYHB1HINPRR7E1cCZaPwpcnA3RFzlMa0ITuZTV85UUO3VQbvHt6No1ouqCPTbm
R+y5mOfAECIG6GsX0LYK2thK06EEY+9YpA+bbnyQJ6stunkJ0YI8Y7kpvRsZJGI2
CTEijD7yZCJvVL3Vz5PgtMjj02B5lteWYZnI/hFA9p9EDDpFXUopC77bOfRdR7Ne
mWKbfMEUp5VCubx5+2oAwfumOw3zQ1CrYythgBvV+obUW3y6fM1Y2tFaMshLl5t1
HUDT3SQSeugKVkJQE5QS5NfSJRE3IBaYnNiHt05hwSQJNyvOTQxPJcIzuqoaCaSw
85VRqEYRXPnory+dPgCOp52GXFjhGkNSlE9RZyWX8GHGhHHhRhLxyCw0Vl2L6McH
xpMqjyyfC/hN3DBdB9E44RWQrMksSNwOjiPEi4DtDDYSMGqQRfh8lAu4AOaIkfXz
1QqhoyMO41k1FKE/D9uCm4spKY3Va0y1F6wnXStHCVUClsAZ7fAGiVohsluKE+mL
0v+T8exa1hxsBrjM5kjSQCQ0mLf/tUSl504CxjnHmTQy6Quo01bihrbnlfFnByak
yW2amhNnoFvYNTNbwnVZUzqgf1GTtti7R5AjpspKNVJeXY/74FSn08yV2JzppVIL
Qy8lhn6M/VcD/5DOTcu012atFToJ/JHh4IOsVOtNXJI2XtEY+RDetS5oFrdFfwdT
m20CTdQ4DJtZ3LL9juDigVGLGwjC87mquGL8TjM3H0hCnhY1j6f69STCDwia1Y/h
ZxDF0Q4tpE53DVzegiply9oaVSPjIR2anzCHEw5e1LkUXR+Le6fYZWLktgL3hc/B
FY9Pxdiq0GPFxMSZzxlDVG+ygaunLhHIaBbhPp/pWL6VDKpPzOet2FGwDNDVr7E8
RDajql7QeY04oL0SHYRh65HYMS2ncsqonRXrdylJa3tKoYI3xDPPaheqiIqgYBuR
Is3IOE9EagH8fWM5AUZxGqtrfioBVF09EpcSNvp4JDEL3Zr/16q8gtGtw6qdPWuV
f4OJNMSMAx2WLhGeb4Q4VqgTvw+t4U8W5Qp/x4Lg+J5HHbcPQtXX5HWDXNombOC8
c51qxQz6fHOApKAaguIaM5L0iqWRvkqjJubrwD76PaNUyj95cCr1limYXrNr7Ijc
wssLZesnrC2UXCk4rlGVcUGI9ECHcddzxWdcu8t9taAR3nF4kCr71ShtJfeLzCuR
YMzDfrDNk1gHL1Ksynz+MeCK34ukK0Ly2ucNPB2BwGjTmuRJ1YPCBpS+jNJlBccM
swkdCNWHzig4pV3azWSXGijEqrLNwaOkiZ/117j3E4eEYncOGXtXCtAAwto6QOE/
82l1mXaMB5Xntfd8dyvjWmToSHNd9cxunwdFevZy3u4loL9TCM/RT3WGVgC+QCNl
wMzIAw3Jz+0euzwLKu+g0NbrELXsljsz4icPPjEFnYR+O/FEJ+bsJSDb7Me0HEhF
5SbY58FLB+mw+fpjRr3o/+5hkalWeEm+i2gRIoezQxD3943juBDfXDLc6Aj1H0Rz
bfBid9sjnDTIRFpjNvBBQBRwVLE5ILzD4cHbkyaWLaNvQwqDGPXkNXwMeX4qZz1o
7x6kf3SGo8/MjMhbyAVM56vt5VehoYmK0ou/mKEIWEiA7WJ01JYrfYMifuaa5lUG
gztPrdIVB4q/hSMPPTyyEanEy//HWElAT/p7oFPA1O0wp1howRlIKKnCpcdb2g/2
NPJ7E6k3cYEcc/aaFlN/SjMx9Ox+lkH62uxi1xVGhjt4bRPzMWCi2F/h/1gXqzzK
9j4Z+s/Bw8pNbZOLDph/lYGypeYlpXEpjyGW8ldc4BD310yLV9Mw4WXrE4dACcYQ
ofPMlU+/lqAvoxkcv1ZBADAzGSaR8gKSDaKdjiJVwA4dWfwbegJ1ChHGcXT8Dkpu
+kNKIV9f4pCE3Sh1kIWPmFhMsv9ZSVDy7C1cc8knIOouAEq9jWlfFB+aSZLBrHPA
awDlOI0cdHp26ZT983sv8OP8VjbiVs+ncFo/zxSKI3+vD53PnIBxPpye4EkFmuki
GkP/pXghsQLpOGHxtHkPDh5wtkYefx6Uw/PPxH+V5IQocvjVAubP2zdJD/BAypEe
Tt79BSIQohHAO9yqyL2nyQBKLtaVdm2n6Foc9SXBiTPRvZTwzmTpt5fekv7w0h4E
ApfTMvq537Qy7d0wV0g6+mbWE5Oc+elegBxugH4QuvQKw91Yv2Z7/skm7FDXShuY
MIB7bwzCRKUk2LAdUa1jj42Lh9CTVY65abUogxdggcmvpAEwt9Qu8eEqyHAALCXO
TtmwwrvE7UYP58ee00922GoxwSCi5wGzhKocyZcFREL6MLYDqUrVZ6jh+aDbudja
Bp+2G/9VlhcUNz9irT3O6gHRT+vWcy1dNzzQ9EbOoM1jsGuLlSURJi511KP/oSpr
8WT2S9gv1HHb3mYhXVwcyLkwU/Q3Fa86TEukRsZ/o4LBx8Vany5RyHAEz1wgsvkT
ezgF2cmjtUoU4NPdrb3YJwbCimS1HX+TDm0+eeMnYLmSZFFnKXKoYYX+2Dxtu0zh
CVg87NoWMGexDG6z8orhfn+jWOnqoz/CUBp488L1NunthRiwTb2clWevm0FKikwx
RC+477uinFaWRLofZknRuS55tJ2R5pOHyHetL1wb+R8Kd8jIzzRsLbl+d6BCBcYu
BMxYUnfeSvtdlLalK4wHRPGBEHeYMBvNkhCzdb2AWQtwNa6iAbLNmzaedsACPjrl
JTiXoozycn8BbDj9HL7GbFg0PRNeqIsWbiq3ucYjp4hFsMgjYGuc6NCsLv4QrR0W
NnMJp9UzD/7TlGzuuoC5XxPvZesXF2byiJnGHi0Kq56hvvPJ4499Plx8PvB3cJyD
+91a7fhRZdMxhFiZnxVHEAYnPEutlIPsWpxld/fdZpArdJykLdXEC64Azr+0BkSv
oGJLAuVA6L/Hp6rEGXnOWZqanv8t3korccZPHHpZkihRX8aVG2mGlyDeuODe2hfu
g3kp85M6bQ4JOlrXy29uorgtZxWKF9J/7aq4fWUoOwYiC9JWbMXVcOn6wvoLOH6c
3EE2KcKFGxFVK7Dxl15ntpEmWkhRnRftgQU1I6n4bV8aIYV7Pi8/3NHsyT2l8EiT
qARAxfWXpdLIFt24jswJiEYCkHd9zIqTmBfDb6rgf2grV1tLOB2bFgFYUo2QQLgD
vUEvOkRIH+it5WD0dejcmRj8FJlhav+VAWfN27RRnxU04gvuVV7maP8PdjYe0G+9
XmuRBGM6Z5IyZFCia3p0PmE4gnt/I9t9+EFz2J23IuYopOe/Dm2K3U/GMhP9OEtg
PuJbibduvWDlMpWlCbI/zjqGTNib1vLK0RnEAe+Hd8+xyrOH53wQmerz3TH4ptjC
mAqWlzfBi8Vq7oxh+ZY7HEDJ09JVQuajQtnx/QxhzfqhpJnEQDLANfYMTL+J69oK
HqZ+wzzIQFpj84qTd4gHRerZvHHw9HkbReEf0J1/yqJ+PPfc7lvWmY3GVuyCjD2N
//Pjb1aRQZ1bWDvgTQ6jWI9MzknUzy79e/sNcqd5tfr2fo6482WlIxOS5k9rjmHE
ohVy9TEYc8/wgL/VLpLKGRUP8llT0r7u8aBSE4s2R3jOgk+yQ2VlcSp+cpQ42R53
p+PxtuP462lHGHjzQHMqbNRL2m7jFHSOAJiFO0Wt1d9XP6JDnPD12RrejZQlv81A
t66/A/pBc4A6E2FKqsJYWLg7W9wr1VzNLuKm6hgHOeZcJkQ2TfC/DIP6AkLCmrWt
fZiTuIB7kz0MOVg/ailCHOKf1nsmIoHzjSpu8Y5gQi9+yhk9u6LdVLmeBtAR5z+H
U8sTcvd465KN7INQxa+XxTdIUYoeIiNKcXcNUvCjKQo15oimsg4Xw4efPHWDH/Vw
nGhdEkqssVjvW5Fz37t8UPtyYgYLIVZmVZIyvJJQHsSE1xZQmNeyG1Ivp3SWQ0mT
isUze+nnp7dPOoeoyxzgMQZLuZIXehG4fCI386z8tdC86VXIJ6eLcQUrUP/gq5CO
tOu+b80qJF58tfqFpUFz2COS2QnR5+ze/WWqpEXuUHtJ4n/GiP3BdRbVOLGVNFX3
Ow+kpFDKUM2BHb8RPxQlWFhmCAMgShMPhh1c/O4CKPLJiC6apXs2vFqYbDDK5tOh
f/QqCV8ZtQOgvqGjB5IgN3TEayWOHwKm6eauzEvP496pspNKoCv7bGZswFYdPgnt
JK1w6dZ06xRTjmkiuXN9wzxslEshKudMqLD6AXhlb8KrSWbpwtVvmsEJRtRux/xf
VIEiaqKkC24yeNEcPk5kxAoMAF0MMi4uaSuxAvdv1waC2kpya0cnvy21EUMs+d/w
fz6ShXyMCxZ2R0FdoX60QxR0RoeCCk9oSiXB761+55EB02WQ/ked4QCgtGImMF1C
siSzNu/bpLofBqp4yV8AIcUpq4ODWrusxXuT40wAyc2QtBDAeo4u8G8i6n/BWbhf
cuqFJ9jDudYHXbj6Du4c2l9UKPkfMWLNYfJ754m7nPfgYm0xtB27PMqL57Jpb4e2
Hyuneyg/Mvr1yAS5hYTXye8Q6r6i1qgxAflflfuLToJEoXGl+jD9K+mt7dMoBeT+
FGmQaxBDxnhTy6zgjX+eFOrny9UO8fXm/xHYJo07EqvSHOBZfd9eYUeodl2kJo7P
kTOwDNwovBjqQpVkY9VaIBQf5Fob1J5pAjYUvkTRD9bcC4bFPGtWf88YzTKqK9Te
eeA5W/2e7hCdA2luhulh333zlWfEZJyEWkLhlDpptnRrhjfq/KUYxztBjw/oF3A/
jekd+EZcEYguoywg2rEmXjW0lkrFI2MeQ6U15XSiv17eqg/OBXK957kr5yb3WurI
QGRmKpOwvOZRLQePFchS7bHFzV+3m9hVsApBz0enI34ekMan6rvNrwCjVPLeO8q5
oLrMiCAAUlbMHNebsKcHcsAP2YanRu6DWSPsHbpIu/Kgbd/NflBoTd/3OzMkgwGX
8Cc9d6ccrm6usVtQO52bGdufxSAff+hc2+Ljid6BAbe81wA0gSe3yK+/YAPP5TpL
u9P7scdEEd8LEZtFxolQHncN4cVw0U28cCSRcbWG2LxiF+N+avAB/TFdFCcVeTFE
cdS5bkZ6MNVJyhbnk9T9sMjXfPDzhidkgdm8bxRUe/vAzH5LS+hwV5Hom3HOXZw8
UPIiO/6EbtwRA7I2H0OIFh8CAbmpPfr6HE2R2pDr0eCN92r7zPP9gZwZQMF8YulM
E6ZOhGHRKOpeDhxxKvJAbLgvPU/QASBp10lOXdcYijrhn7/uaFeGoIz1+OnxqUbq
h9p9On8spIbcCCj4OtREsyq2dYWAKZOkjd8gbzKAi/6b/2cDVwzTyzxNUwXvPrS/
LRhWzciG7qDoxremAZeW4Kg9nZetUpWWJr66tTlmedK4ag7QCTyj4MLzqlAneykO
VYvJSfeQd/gnvQ83W3+D68lAWZEjN+YtIsBx3pc6Ses27ATYXYGHJNQ4Iwl2ii6n
M0tjmHJgv0REhR3HBlrm3dUSLzd93uzloJrLVk26x0lPfK8PPYffuNeKINRfMVfO
yNJBweqpHpcmdGMeq1TVaqRkUr7aVPHGoFGdeiKydk41hNwCMZ2aEWu8Q+Uw6zff
V1wmTysqj9iFbXWTPUm5YYinKeaJgD0rUTLc9iucEVfXJSUHpTQB4TRGnrd0g7Ge
DyC/Nq7TKWEzYVsJ7zGE2IwKdJ2Vc9X7QvV0Hpk7rGyCaLc7M6yGrDpJF/j9wVTn
AmAUruW6w/2HqjXA4XlzFIqRH8NFEa/PyqDk58isT6yglSH1jioQbgSmqXDr+jFC
kABVFbLvbtzyXUeM1B7skUwS+qSN1y44TFw3dcwdHvVqTiPDT62lwkoku5BiBb13
XWeG4Jh2jptIF99ghfgcUb/+fWKMF67HqTUln1fic9huqaTOWpPaUYWQmd6unhOK
DPGfigiUsBckvVqFM3ZQKUC/+7bExjgem0c2GDOfBdnzLYGcLqWnxqU+BZj8xyWC
Iapytv3cIfT5BwqLcEAHRreNJOtDN6hgBmsDUeJ9+0m2xZGNt9OR3F6zqxJ7WF9f
BxOb6JqlPvaQtGXoCeDVU0ysLZ9N4uZf658kYNKp4P8oDzS87LmV11zob5GZMFgs
eyLknhI4YF0QuZ9VS97NXe6Y/RQ+IFwg/VAfbsVWXVnBm2csp1yg3rDyMMJo55j6
+Ck1GkaSK4cWNNBlwiC27hb4ZPyVB9L1nJ5EtodqjnZqAA4fb2bv+X883djxzFy+
AaiKqVOSppjfTN58Af/ApKi84fa0aa32JSunOFKAKWIvKGNCWIT71JwEU3Zo6J5p
G2Kxt5fvRuz59XtDZd5TaqiFqrYhzKZCp98jjqN6P31Sr0L4xD7tq2JkFNwTRuGH
f9Kj3rrjldWqUgx14E97EKy4Ke/NEn/AsNn2qIsuRHTRYGowOINyMdEFIB3ecAzF
2F3TtOnDGO5nmdJ7IrYGZXbzm1h0YRyYZ/uP+p2ujDHJjAwdUjcBc9dKC3WiRTF2
kYQKd1xVIi4r9T5fCJQlQLQOW7W72ihrVVtS4sZ7ZTZBsfoGHIKSvCB9NULn283r
kTjb5u/ko++1708aGCgfs5FlvqIbtiZqvLoG7/aFF9wjFOU5lYVA5tOxb6fHMCfX
YcNczz5wRVJpHgKou7amjeFKHXg3fIN8Q7mj44L0QSO7naC8zrXPJgfkS+iFkaRl
Q2MX8CT03KmYGolbe1p/A2UVXHwgdDgKE9Bf2LmrCiQRs2rJOAq6CTEIGfWZb0nk
ay6rMlF/Eixoe/rffU4skdN1j7ueKgjEJTDqNUBq6edBWaMwt01wO0gnCVgmpi1t
TSK8aN/D54gNks9tZIslD3iZnWp6590GGXLHmooOH9ipssV2/2koSNevUliqwUYH
XfGXscU5Op16jitQwMeB8HwEk2KkmVd2DOhFN+yy6fvatpZroJn11M3QS4+BRc68
meLEKkQlhZ4hhSNesv6SvxMxdF0aBfxUG8W77kClBWDKUO5ACiQCx5tlZUdoj1sP
rrSpOBow5YazdLLrQAI+W4ut4InkQ4AgqXMcdsuBBD9oIi9AYuOAlajX5s0Z/kH1
Urrw2gHzab9t1y4hH1aOeTU49FYQUAeQXklBxuVDH5ZPaStIb259IkjVIKRenYY4
AiXTxeHGiRINFJFIzEXREK9iqljwYaRE9FNWFgrMjPq2QNdCNZcdWCqPDug7gLxz
VvPh3lr4RPIJre0QWgtC5pPmsPFjYgURikt14J9FGx2AWrrOiE5LgSc63XZVTtRI
nyL0NoqVEgxRMA+7XvRrakk5tp5S20lIXpRTR7UPsjEqBDMGYl2r67mKPnaNrev1
8iwPck8kc6K0bd3+gm845/VKvyUY5lDUBtkdY1UaP5Hzj3Iuj96LMSZHhJifz+5r
gWyHFKkVnQEeBlgooIswEwGreC97egplcE2d4RRw11ZprXMC6Hg557HBCLiAngui
+ZwiLAvAZIfcNPOgBEqN0QpeMIHwQOaWBJDz10Z1aSHDinxXkwM+dB1ylTe3KV20
oCH6qlppOxo9rUbBnuXt2LdB3Kc9Q/lNa4IK1xcIYU759vMiewkXh43daD1EmUHU
iDp9iFnHz6FC8NtoNNU4uKlhlyaTIMwkV+S5Th8bhcI3p2hmOO4tZFnjX7EeKzkL
+4wTvITG4pNLhS4KZmfnukBnnsbEGDZvgNXZ2JQkDoe5ylP9UdP8Qia9f+Cdbp8H
gr1e325nN3kZ7NVMjKUOLUZMsvPzzHEMirCAtZb6cpb81lA7U5BvcuJUCE13L0sI
FAI4YLPgqdd2HmmBh8lON28zfZK4z1zv3C5X0sNQiarITyEdekl0c1H7BiGlHwua
AgR0DBiMLdjKwtn/f1muo99JeeIPogbLA8Or2J/x0GRwAsyDzKFkWHieVpBWmvBn
WzCoN9tH+DPRpDTOcaZx+S4gjmMqK9RKqQQBxjifivQjLOWcbafN+Xw15uG9AGzx
p2XYJOljvVniVmFa3qvktN9f2nclu6BIZ+UcT7Xx66d5kWcRfW0LWSpuhxFF+nO7
CKBfaw2hE2p+qUjUd4ImBty+ojxFHRN5bIJTuJI9Zdz7ytAy11ojNupdzlSd3Z34
jHg4991aK5L8ypntNtcabh3e+y5RqLpbeIAMNua2GwRrW1ZrSF/BBudDGD3FTRZA
CYvX59JCIFlot2040oNpKsghtu03FTOS/as/YIrfBDOQa7hJvIIpAROkt/r4rS6W
kKL7cIo9MleDAkiOenbdxI/G4X6OE7o6l+qofMwqgehUFH53n5to7H0TC59VBqV8
uVUKkcFWnOzxwemNjpaGP44PCMmZ/a0C9LKdO5vZGJS9WwhYQmTORWa+y8x9vxKv
W3u8DOdCFZhEaHtuUcxwyP1RpyUJ7bc2nylq30TzMubyKiTWKKd5DXPPzeEgad3+
UNTQiPV4xsxUZhcy1kQfZorfvZjjJtje3S1CJArkoiDTfhCBlXOiy1I8KGn6g7sB
s+oq6pr3z8KjCCMQzRERdejx89y90juzMBIRvcr8RbVJ2QT3iwMXGSIU60jkcGdu
KUPtnKckO2z240Qr52Nm4R6Ss1+d7vxUXITpYMKvOtfvVlX2WfRkA1938+2UuVV3
WWKORuu/dDQaiAVuhEX+qxDiELNTb+SkTLgoctx1iWS8Tx9Ppnvse9OAcuyzc5FX
noZ1QlTYgzTihZq0vr7/oINCWCc5tPgcHAhiFaZ1k2ItTKXBipijbUZh2m2etj3o
nLxx4TG2fxw+0+PjzaejdGIm66ZrcdZ3/jW0tVDsm/1O1rX/M896ZJAjNM9l61aO
QXnDLvDgPwjicfwUMK8NsrodQWD+byIHE6XPk8ifEX83MwU5sejKfQnrvgQOOz+H
1oCkxOg22CYofDiv4FkAA9MEnd1IxgVSZ3dc35+3VoBzugCE5PQYweB2l62D2SGo
mUIbclAiNvqoreVQYdSpy/seY9bAq4eDHPOHOMKhYuHfWmaVj8EFcIN9ro708Cxi
vBftbRGvFv/tT3zQGeMIaK2O8tv3YI90mwoAllovMR8duSG/hXVz6zVngkAk3hU2
5GYhoE6HviS2GrKcibIgCvpwrvSTtgyO0Hfhem6x6PVkKr2HaTTRk6lgsrBSjp8j
O2/0ybmQbh0zSAGdxul5qCSsC0mFOlrI1lWhzTtN/gB30kwVCwPwdzuG98h2PxQZ
prMelQT//TlTKlVath7aWFKW67t/QQBvCPOvbWXem5Z+yhrWTT/w7NjGhItPoOqU
ttXi3Kam+n00+9AS8Oy+5E68B2RQ4Lhkp7XK8wShjTeqakJzoZkADbsNVmHc7/mC
RIqmdyGKSYoKBqzh/OAJkqqm4VfZG6Qq7pOG3NtqvO88G2SvLObn9YgPgzKtsbkJ
gXbKbNiH1ZYQ9Q/lej1NY1wfk5ChidkK47o3uSBYqbtgpb68wC+cc7yQtt27GfJd
66V5YFzPP7EzNvEhXPQO/x+0fqL0XuMMsCVRr5h1j1c6ZrXu7BvxZxvC8puNe5GR
Rw6J4MBXnGI93yvqAfyr96DbfspahypYcnK41//+LofQzJYnxuv04hQpPUo8jOGy
AnW3eTBumAQTuoQHDrpV0Dtdng6eiZgZZDi9KFeATgdDsbz5gdLb78fn9ms0K+Zm
Pew11SdbEfzAJatwDQwuWALeMSL1OWoBAIa7Cv9/bBaJg1yBTMpLQ0uPuj6Sj1c2
AplyQCr1Sl4OWw5ecnUZi4vq3UdTNlu4zySrWSeQ6nCeP16mPQFptTSUmgftNKQX
TFrBVy5nNkySbSAg/h4I6ZrKqiTbATZ1+VvpviIG9hRBaCrdlpnM8Oe56Ne5bfM7
AYsLI2IPR8spLN/pqShqJ1bMzHfm99md9SBzfEd7U8/zolwCCoUX86CqSZLtyCU9
AWFkypszwL4gWEWGFiYYYR8QIlQ2Mg+6rb0pT/Vk0QRoRp0J7zR/RmxJ73Q5LW5a
yPyu9SOo6ixguigFddPgMuOPm0FrXwF5StRFq+A8OdwVnW0uj8JUt9w9vFeTZBxH
/4Ys/snwVZ43akucTRcEPwC1A11tTJQFi0kEpy/FjDNbp5Ui41oeI4uDZHBOP5qh
7IqDxfkNKGqzvujfCEAl5RkbxoUPGl1lvBaOy0UKNsn5YIs4hHcezkQ2GRrdlpgZ
IrlQZnp3QBWaxAot6/kaQ8hC/RS90myqwsgPl0qin2CaCkW+bu2IaeIbGTQJhKOX
+kUztLsUvGrAODl58od0QYEu39kGD1LewBzyA3fuM0weHhvhiRN0sHwlGLsGKyhV
V2ZGKhQWwtkisjQ21uw6gH7SD4MQw+orYpo914oGPhmalFB8Mohy/zuD0DJqoB6h
+VBB/w4xgmxBCpnS/fzPoNmbZU4peErmrya61s88bbHQLLe8wXEF2L4XhSl3/bJ2
yxhZKYSwaxcpo3FBargP+FgMD2/7J/G+Viw50GXkHLPkPilfJrGKRmmAiG0G8CvU
YH4RH/hSBCYHM2MVL8vY3sJnUtkFt3ezDypLg1Tn+/snsLadOH9h8oCqlcKevSMN
DS3qzYbZTmTM2+rEutUasLXWBGcj3v/VX6oBjx+chCLKeJGFgChmk7gDfL+5PMpa
aREAHM4dTizG38z2y+bZ3CGImDAq2IlHKmzYVvkQTS04hFB2NPo6gIvepRh/SNpd
9XUAh1rIlXccCqX4i9Wi7VknJ8S4/ak1nAeTMvQ8gse8kUFeMTMYS5juPQ4aABn5
j0ZMsN1GuzNMuSsol4D0TU0tNnIQjz5083ygggAAzm/Bzo8C5t5QzYICTtOM8JN0
5OoTzcEc7UwhbaRqcP1gEwPZDV87XfHz/zgRKuP1fQr/wE9o8TRrMBgTA9sI0F1m
m1TxiolYHB0bBbSUe5aD9RBOvY9WkyCQwyMkuK2cUrKG84G8xFolm6yNZ2r5VfIf
SZRjayAF1oEXLG+BbHlvzeaj+PgYWptxqGmazZb7dgE7ytCU5J+OU92znFeeILff
31cwHzgUx3olXNwvCM3vWiQklVPP4f9jbs+E4BW7FxkIng98xWsTDcT8+QMrHEiJ
a/iwzycSE2TzSE64E1ZDEr5/S4h/hPVC4mtfEEdfnCQtFJotKkVveQ41cScNLAa/
IxPo9IpGrshBF7EpdRBDatfeeFBy3GBM4GBMreKCBouvRB1MZbpOjdlBUKWWOGbO
juwMPYI/Qf8n1O1rT6sz9ClnRSY/GXG+LAou/zF6mX/EbuGBBgzSGSmdACdl3eEh
jUbQKDwLP1we5+hPS9lnKZbkORVdHyU5D+dPnZZ1jRbjckfIdcFUPiItUZn3JMye
6k2P3PYDKtIH3vimERgR3U8hh6qZ2mvaM1t14s8DDMUS8jtXw05MyY4UYxiYig95
gvRx8Xxk4D4vc4WEn2LaIO+Ki2Q/dXjesCV11110n4I+WnGGZ1NaLs1pU3pct7Dp
BD+rrDF079XLgk8sawZjC5Pk1ddZ+sv87rQZ0ULA1DWQfs0rio9iXH9X6eF8zHS6
fnw/IO6e4EIlZDtj0a5eUehtS6woAWzzwSy2dEYxo3BumkU24mLmx+VjtPL37ERT
vwr1jWhZvhn1Wx//02S5bXxPefqXeLeLXsxxUfm/HJSrmwKyrM5UTND0u+k/y6vR
gnEdO9fU5C0M7O9un8kUEOxnSoJtSzsyLE7Elrf6u8+Qy+XzCjwdLlgG7C+NgvJD
1XbRoQCUzH3xyFi7SK2wlPsZGDgQiQIu7nVL2kX7zVd+NPAbwaVL0KjwAWu+I4RN
LplvAXDrJur2HV3Mw6Tbt+RSw+E8ntsyxkZyymnQMX5LCUfN1HxRSldNtX3XRux8
qKkb8FErWpkAxggSuiN1ZktLOMiRfHIS9VLeA8JN2aL8UxA55HBrzZ6kZV4yy4AB
Gb2oKzLq/YnHW5k0CJ+ElQJ2fwdgjH+TqFPkZWfwihn3WrvHF1yiCVxJCLr0iWoG
C5EOFQY4nyJdCroPIleoMZ7Z2y7ubgCnCZZzx9Ek9wPRnKQyJIkIs2CX2RN/wvVA
eLJtCD536Cp+66gz4nkkXh7CFW4iC6MRYhenBE4Wxcjr3IhufAopAgWGJfloE5la
ZWvDRFjwUPjyXvyC50zwYhyjZoY5wC1QIdVVQkzkjb4BWksqFoS86ReYJoH9GyZj
LJT4GdnwO6TOIn/EGIF02X50oFI3YvuRbOHdBJW1IN2aTuHDV8zWJqpeCIOzHVGU
j9XXhuOk4H5LzL7JQ2qIVvfsvLPoRBWe4Di931oiuY9jZXsnt7xkS72l1OPZcyLi
bVIOoOVY9vUyaESerjn2sBS3s1ODmbX3up5Rs4QoEg1/cuqWR0d9yJtvkBzh7rSL
esoy/CN4HNZRQNrTBc24IRkWIli7p54Of0jYCmdqmu8RAKDanuaLc8H5tizqDFum
B4sk1TuXyIie+xujBrhlrcj3bii1GGDihf3rVmpfF+8h/69dNYy17BVDKBjgDE2u
3+akiP+Rmc13elljmPWbXfCjnb1gNGWLJhouZSzEmkZDnKeHpHdTOOU2B1IKiRsX
St6snxG80YMa9YFMkQDeLP8nGihwCrJJUaKzMFdzrdG/frfFlNLsxP9jRcSGwaPl
83wIj9Aut4BABfHRPuFjTfiBcYettTx0Iif6aHwZLTF3f855wPXc3tIVuevvUeO6
RAqewrE6wBurXc1tMYOKPc5ewERh7k6vITc254c+SeVu6WEMaC2wZMV3/dIOPG2y
mxqNVg+GBU1ChgmrdmrOaNAuwmezRqPlelCv8pOn2QcdplSTx+q94bxqgFAD1qj3
18/v+OCfJD3muETjhvPLrLuvj8uaurumVIdIIod6HcO0f06wAavXRm+DR+LU+z1h
3dQSbMAS81WMGPHOF4JhBFbq5FG375wg+IM4AlZ5G/xQc9I4rLw6psksgfDGKy6/
jlu8LrlnG/S6Q7mni6oi3VgRCs4NTepBjB334VrcYvsr6SrpIIc0WvkU5hANofJa
2Lw4dvfcmkiRifW18423iZxBqYrDupzI6HGSF1aKh88AyzuXDuzir4KPUTl9Yhaz
NgTGyzylP8MJWQCmgIhcSWMJyNFhPHEb8OjlXNNGciNcunrWy3uhZv8jAIzAxP0c
AoCxh3Bn7pvTKLSZ3CjhsSiaj0BGoKTzGHL8ARfdohvAhbQv8XcOodDqgDs3H8iz
3Lognl3FG+kCqJLrJbZXsBC/6dlgs5zbY4leP5Ghoml58QXB1mG8zMwExZ5huzsp
31I+k9dJyOkmgh4k/Jnvv3wDWfqTF1BPR4vihSpm7Tzy0wectofyHHNuM1zYLRCo
xBA4r6pEbNGHlPb/yDO9InFfasnTrbfGoAk5EfXXM8yfk68kXGbpmAp9ApJcvUaV
0Z6hiRVPxPbj2hQYmGR/yk6h98rqcqEMpmNzNqx4V9P5K+57IkRNaOMM0T44sRq5
+ARPeDzNOjrhlREqW4Gslrd2Y4lfJ04szlivxnY3FF5Q6vreHaa2X/6Wzr2YBPDb
puWaFgXfLn5UOaZKt4xRmNaTx3p6o6U6KY0+3mc1typ6U0f/HUSgY/f8/UAWyoqa
6/pmAA7lpLCqPv7m0w72W/i/INgR2hfJLFu3xEeXGHEr5Saf47q3GWLGZMfMJTTp
TGQmEyvJoAkwhaJ1aC2Oxf5UOQrjgBVwE4Yv4Q0CSuEOLbsUCuiqYbl2fdHwnGhg
VnUfwqKK59at4GGvR7S+iV09rw0Tft/JCM87vKwgXtVog4/s0SBtCi2FpdFFsOSx
+R+uBKF+xumIwzFPYLemq6XxsxVt7abLpEEvDIPU0Fbj3yu/EPfODbluKhq7peJ4
JkjfUD6V48JUNKcrRUleUMGAiLs3fz7h5RMiUWM0hKAyXlut2nFEioskgziD+j3d
FCjVcLhOd8ivEiTN42N+OTfJuYZ+518haEl0HUSSQTTnX2U/RMfeRmBLtoPtrW2T
lLxUOe/cs6jGS16EHzABkLs7A4jDmM2SfoFpJOGFa1koM5GUcqpsF7cu9r74d2zE
R4OJpseznj9OBEGJANfT/qn3BkIkQEWJEp4kaV7EfFunvHkQBFHI3iWB8qcxIQjE
ObF2xCyo4I+mf5H3U+foO1u620cFqNQHaqX7cs6idysHNGWq3gkQinX7fGCC5QRe
n6zQ80ia5eohXnatt8wxGDx72DcbpDj+zXoGzl1caL2+/bCkNfwXr4kJbYaXa9KG
UMBeLEuJnqsXYIjhQd+RO6MofOvb7iMvxGnMTYm62yZqhMqwBLWFpe7WjLHak1zN
N/LpdAzjRoi0raWC5o96X0rO+7IOxkhe7dN+1JS25LvkCvVFEJnOj/qKEqE9g/JO
JI3rfc8E+1yCTcII1gvrqro2J0XlcMZCh78SsHbNnuXm8fTND+ewANIx2lbR9MDA
dvvMc6EmkS3GcaNgPZsbtuF+20BfoNck4GWgRlr68Li/LlA10GV/pfb6BvH7GoZM
k6GR7neWsvH5zpEr/OstcCTNDb3Y+cMy+JnN/pSoKVxylzAZGnbg6kYkrdvWfkRP
4SIwp2Gy0hvTjLH+FnveIWvBFvnlObF/RTVlsLN8Y+4UcI4SoGX8GRJfmrHBqGjt
NJi2fB3I9axiNmNOZmJ6ioOVwrmsO36jDzAtJSrZ7YdrHZatdB4OWzjo57oimJYF
+E2k6QockUkM5zjF2JdlQkhOLulWlxJFoBmSW8BnSzEvd1pfAxZv8oZ6CGugOjt9
GtCnZOKIBeXuyiCi6KRSx2VJQBeLjLq5EGQJXGellB9WDCtsDgN42XCNI9xECSqv
kX6hYCbDOhbPQFWrvZqZ5jYknEjFF0RzUO8nO8VQHWqSyi1f8rZ/3y8HqtGBNSIR
gS1rCRH1E8ca5MGd+LX5tumT6aPMGhkLYXns2PAHSWmIoiGkg35kz0Nu76XtZ5km
KKecbBhIJ3Xns2aLcMkMBo/dWpXIVlUHspyA/+w5vGSwoteF6gKU+eiVDxzXlo0N
mb613EsSV5s6QKBlUZZSQjXEZ0htlq0YYPxZRotpYhz4INbHz2esOYxsoN8zdCoV
AepK6rlp5DN3+m2Apx717g0mQSj/EsxrZKyY5i31RDyI7VOYWVGeLEtdyuoVAJNx
QjtaGIpa7IZ7nVpu+p/WgpVj6MnmHzM7lD8KqQ3NO9LAuamXllEqiz5lSgtdf0nK
zxBenUACTEZUpnTzTuPLt9Q6vgt2u54iEWTUhxCj22D6lvr1zHyuqgjYos5S/CKE
ANqGFVnn1srPioywKvVWrwtmn6JvJkfOYI4MYShwslEQTqMVXUcEfkUrftD64RDF
V0Np52V9BX0NTF50tQCGiehFpbol413EV7mGo/qEdIwDqZZjbQR/MMmqVop7Bp33
+tAhDyzgLyEHH8ECTVakNQ/memXpsoMJ/zTgw7lekjFO+HYYdozfSyRXkv7CPBRQ
AIYfiOW2hrXO2I+FTJuLu9daP6YKkPJvE/ME4muqiE0Dc0bTMD624eNEymipz0S8
J47uACsMad/JzhNTEYAllBWJNyyc9lTwXRMtv+LHItNF2qCCP/EmbDtagXr69Dkl
UeZIJcar3v39yAsgzptwMH2bjd8n89cxdtfZzF9R951BH/IC3mYBAXOe7ztuVnUd
UZTEDoZTwUKHMm9B2CJoTxghahPbvqAUry5O/vV3vlruRk34fI8sgsEPULq2YAh/
asW/il2PJu+7/Jn0R/txTID1JjVxlOaieBwLc/ev9SYoZVrzkP4Y6AsPJ+zGFrWH
NjiK/8vPoD6ekgPIppIgj2IzYkEsZa9qX+jSHheYoyVN1QCA+19IPzdvdxbAvvzp
NlR6pcjRT3N8oNqvEllVizkIvPLNVpEkOukRiKWhekPOFCFrNWqZHXtnjdh679Sm
uqSQrv8njao9cYWW+eT6jX7+X/H/UFwnLCPqW/HnV38Oq2tHtX8qPZx+GJDcBTbr
Quk2Q1odPtW91xxk+xEa9JlFTqiHnmWh9bdHbGvUILOKHhqg5OQZ9JmnKTqrGFWv
vYf/bzJMlJ+hhqsusCqWp6AC5XchGhns9m81nTUNHWdOHyJeKwTnhMpwAG+Hh+pG
JvV4L+JIS1wEqkEA8dn10ScOonjY3j2q/K7Ddow7iLh1r8iUBCojv2e4x+RpFQKi
HwNwOf2KcKQRG+2hFDB3/yiIHOh6Oq3Fa/z9r7Nje6B6VqDnXEbppy+tzUlxfogp
mh7AqoaAn3MTDXNlwApLkJINkylJsiSyKI6WP3CH3335xr/DI2D50s/SVzH0Uxg0
9FE1kmYhJpURDg84RiLjJ7BkBMT7STzA3jM2p82OOY0GoM/Hd7flsxM0qosFZWYf
+pnSd8rth5qgaTFcfNLstLyxCDn0TYSGLOQMQlrBsnTevgTkFbRDOcBqtxjLyDrg
kadJiZRINT50YJeOI4s+uqK5/A/wPcQdNXVIjMdHE6xofrM01Ugidno3IhrM6CpW
+fVUihLEW+eZB0rpNyJpUQXk7dlI4ycq2CwhYR7QZWO24hSsa25T622+EkbilZEo
WHj4J1wbuyTbCO8xPqzW2n6tWTDi1JyDpwTsYVGC1NgR2a5ZqF0LmcVL/M1F58En
aSZnjZk2T/TZ44dHM325+YUfSvagYaVM3TosmHZzuwTqkBnJtYeHltQvk2Di7Uft
NjpqEs36C011Pb4ZrAZZNICzRDr7lReukZ3HI9wGuRVz9Kz9tJKQ5txl1xLpNJJC
MYwrF9aEkU7fv9f1gQGGbxTGaIixQXtPZtCdhFjOUgJ49Zm6U945Kc13AibhpwSV
s1proVYI67JUKy+k/0UM9vGTpFRQ2zXt/OW6aIU5/QUT1MKwRXeKI57NaXsxP4h1
YZyBgGmKSaGKaBzujAHEyl8VjqoX6b4uS+wONxX/NrVuvAJXnel0LIn0axEVCDTO
5sNgRTPxm326CtNYlwtEb0BhZvs7LPZIRcynK9niOXhNTmSg6zNzb6Di7B9DMQpN
u5yKdRw3uw55qgHEyQ71D4Cs+FJWqjy+Ki8vRYNbN7USOzAmLJHb6jw9bZ2CBq3i
RQ4lBgQsEdnwZXIClZJ+OdfhO+S+3YPIru5MlTL0ot/7Kdr+gtpxBoyWWHST/Sho
WR0pfR5rAKqHV69pOBgdWUPm9yACEE7kflClKAeTphlxzxWQez6T+fRQyq4s4vmA
vmC+u6a7wgwAJABjTv8RUIUkqKGFXKAsBPVTO2oH8JCPvxlNQBGqnMjFh7hjVcbJ
jExGafJtNMvDXc+SpFdyutIrhK9d9eu2R/TfNDzsuxBBn2cNtv6gm2VPV/ObiAHz
rG7Fsg43TK/ZoBshxjEdic+FRySSgvK6JMiGrGFpvACsqr3ucYhzHEoR3MDm+uuL
WYemEmgljF6w0t+VzHEc1W5oG+wus/ZTXcBknw2Pi7/5UrnsClfaW3G4OvetTPML
0F2ja+YXtgOhWAEkY/TChwoGIMdk/oIsCsgyrbfM1f3dE06nOiIRbhQ9VyLl7byd
cBwaiCQmnXDEto1Q8ohyiJvtnFRqUJHZNj8B0vCAhfgLItLQa1VK247bu79ZQYo4
WetrHkbOBAkZmVVzHIZqRicM4yjPyfEPuHrfBo+A/QjQ3DItkNy2ONQkYzRCbX5D
LxKUQwOlyywJj03N5NiflqkJVaGYvWNOZK/94H72fzV3rciJzkz1SJYRdtxcgOd7
q0gZ8wNoHyvKD1j9uJz2H2a3ygGcSkkdBC+skhItK94o5gfkXC0+D7Tth8Us2LIY
AbYBud00jhufcfADXgRWtodngED18LwAeXHX5ElUwaGj3XWOmPUE6SrHzTSp9RuY
TPDXpzJgwdh8gcCTkiwXaHht7vJRIcv9rbHWzC0bwSmLwQyRr2k06sgXxa7KH7DV
FpoV4jHwGY31/aZ6RwLoqfOly2h5Ij3EUTX71PmEv83X4KoMcQxM2CXQhekP/30b
w4JVix3mW9dPguseCJiC7RASOoFxbGrdis3TLS+rQiABNw5bVfKC0AZOPo7i7fNn
HAYeE/v2nW5lUUbbYb4N1RBQgZ61dNf0Z+1bhTnCDsXXVnfuQkB5ZJT47fFSrAa+
h1Vq/jNx0eQ45CzhkFYdOtoE85pRUrMjiUWcoMCaAITy33ARyFw0vUX7QxigS7RV
XtCDQLK3yAjUK6U5nm62l3g+WmyVoQPOwaNhwAAXPIBa2SWXXY4SHfmLJ2/HHlN6
byA9HaKFnDeK/euHoaAZFhjEUbuxmE2Kzl3FA8OqESoqhaWf/+zB4QbqCMI/T0ax
KbMMMBz1Zj6ryugmMuRE/8OYncYxnhYzEHS9EcmPkWkTly/0ngBJc7wKXbS7DiMh
iR1pUXTGxW/QB5iBGvx73Gd8yKa9Q1lk0j7JYldmSs2S+y7cSOelb+/2UbONZmJQ
KGs9WG33zPjOUff1ZmLxN+vnApcyF6Ze74SwL4fXfcrZdtJcZit/KGuOZk/Z7RDQ
1LY+JdjnIoXKosRdVGxkVgGF0XQj/B7BqSuvLbSUfqSgfohksdObyw8qBAp1C8zD
zRDyPnDpb3QjnXFXiY3LgHeyqiniLkNgmCkdK4TmidDdwYq47u0H85Rx4ZbRWdqb
SR9ehaQ8QzwrkAIeDdTfqSUqtjtPLEfT7CaXdaTtzl7IyVtG6NZ6m5GeQHy96zvT
stuS+SOwTWK2bot8NOO4ysW5p3a4XtqrB973uWTVh/jZdKhewRSfkZ3sOe7qkU+n
WuEipIQH45lG20sSxM8UZBjo/Zjv6RvP9mcTl6RZJi2OWkFGVYCjHABkA42dvjqI
pLxIrAG/vYi7UIZTEiUlIyqyzn6aiOJUt7SfON9qDUZaGXEPqAUTnqphI0ynkRHs
T7BJSQZn6SMTw3aBhVyHUrm7cT1rXTArllZ4XNRkm920dvTopsD2P1W4JR41N8SH
ZuKTfxSEGAgSMtJl2ic17zGZ/pbkkcCydsSW3RvMLtIxrqefbp21bPXf8+GjAgU5
/sxO2ZMzfbJcOMpAyb9d/4NRiF+mLwUiapLZy6+70fwTS9jdLdaLm0WhJ/7Xf3zl
jZR6SuKiwpTgLfNhK2vX20RM86FCCnmuNrPh5ypLGWdB9pTh0LIWgKAD0/p7RpAZ
/1qKPh2F558NZ+/ia62QHGx3hlKuxxAmmDM69Fg47npbDYoekLPRJHzdESEktXiv
CDatm3dMGi4737aG+6j1gz0eiUObT7OIc99gcVtsHl5oCwSqdf4hEAt6IpURwfS1
Tf+8VkWdmGlSp0N9lCb6rUpa+7qpSEKpNZSmUlsJ4/KO3K0wbjR/26m8e+2Pod3u
50DNA0mDpg2BT28ZfAn9wj/eKPR/lo+sGVJk7pLwoggPPH6qpcLyNpJTscweYmrp
8DJZu2EBsgcNoGvX2PvBYebMx6FcpSX/8wKff2yTM+3wrvXq7dBEguFYQxSTJgT4
ly2SgW9+ZF3eDF6dAJ5ywQzQPAgM5RHcQu8thunpyM4FiAPLU7rgPfgKFZ9rPHF6
rpEhvC4sLONR3Ry2rsS/fXDXJrI78mYb1sN+bP3uk/BnwG01vOjoBMMvxWIcpiRl
lqY5ARGUwyU/d2dpUYBissI7DMDU7Z//LC2GvECRWPTkdd946/9tA00vddqo3RRd
FSfgQJieWKVO6DtXJDfMEuVSlAJhIxvvWht9CDf3XtIa74d/X8yl/25PNi0pbupY
sqh+G4ObLgMuVvkH/fgQ3BGLBr3l7rBxVVKLO3yI6brG7CqxlHAHIoC7ZOt8vOLm
ud8/+sJfd2p1qTLED3aPScp9Jnw1meOoTKnESWbXPP+SDvtULN1P0RbaTPw7QfAB
6OBZaQ5Y9OvV7uWjU0iVnginz4TtT4xuYy9rIDKVwXBDNBW7eu13j9zmQG4DCAYQ
jtDAWjrmkUiM5ZrtrehdFad4i+JhAj6ESRMLKdVNvBksUVwkRzqbdionfg3MD5AP
sxP7LQHbHGW5JkQB1BSr7mE9R3nw4rvi67rUcGmUHTSZfD7gPTudizu2QHvgJkJX
dWSmprN4QD7XyCc/9lNkC/xd6ZZ2lC2+vVplgBB3TgaMSrAgxA64PHZZsOdLccnE
wtfbDzfpiNPrP4XU8rGqhVH1Z0HrJl7/1sw0fWAJ1MCvttYt4EV8BYR5VuxCWZjz
cONtCMEfKQIRfASWV++gXRBwn6nrgO1ytSDyj5l7YvJYx3o4ySQZ8ozdjbLfxh2L
pL6xQ5AzKiF47R82FQt+aNuIJsWfXiFgIdIllTiWZ3jVANBPqdgRAtx/eVB6fL7a
JAUuroThk0/gPT2ncLtqtfbgISmgiZ8N+seZMxnfVG0F7o+rQYXEqDWY1M5YTa3f
RdRh02Lwj9oMC2D77WeuZayKlynDfA/CHqUXKHVmFUFGWKD7J5GCZk1cWtSaVu5U
ZjQk3IRpYJjMcbpXA5j3AL4LvbuqVSKVwre6jkzLmivPJrrD3Zzya9sUqVixSu04
05rOzA9ZsIf40zhHISInMQmQURYT7mqjgMX1iWgBH0amDO8bxUh/mEB1ArLIvvTX
B1A0TTLCa6rsv+glAhmlIospvclZgCqdhTm5uoSwiwZ+ZxRbMC5JDCgd+a8ng8tS
3YlVqJ1aSI+05X5MhAKcWMQT0VaiyO9GVcrVRDdYE2vJhdgdPZWvgbYkRkzA77b6
vd7qL3RWdM9lXjlMKrwu4RH7bUKoCP72uP4zLeCmQyoKX6Im0L7PIgm0aRRjQ6cI
fRiaHuuAdAAL8Ekhbrmowm0hSHDP0NRnb2h83VemF3ftTzB47PhCv9/TWkC+2R0b
YI8TiAKlnK8zI/fLe79xpoPBpXoGHrDj9/h/9m9L36bYzs29TQZx1dEdBqHNfx95
R++GmXKGMnbuUbon7B8na3VjelmYF8TaWT+hYemTqu7u3N60DpgBVlVdjFggmq7R
ukpceL0eB30+QABvSig1Hc7RSp8iM/AHj+GITjLcyg4ap+DM2KhEFZ2EyF7vCBWa
zIuqx9AMjh7Yv+w7jDzxgzj/LbFaBDgU110q/X3LuH/1ZacoSTGDRUvlLrzyQmEJ
ELVRq3QZEX1LWZR3lTR3Ihr7YUP8Le6PD4cqGSI7fYscaQwNKXtlBAbrDTdJd7QL
tYtXI50KCbTe0fpuaLTF62ZZ9ahH1MobFSrVxZoY2f/CmY8utav0Igym5XDivF6f
H3RRznEAet4dQFyF8ewLBFx08LuHeHtwrvFeZX3fIAgvNwZFQAOgBIwErKrf/kNo
r/TuoYaZT70HVRdgK4UIc8Wday5xw4YymjIMzuTInzYMLqRwAo2PU9lZj6YM9ukE
0E+BRzBBbbNG/sLdO4NqbqJn1K2Nulz6RD4fwYa/lIaGzR+2u1d/h3Jy64o4Z0WX
ERMUiI5crqPOVIZMgORrapzUT4X2Kp3XsVjkNBaWNfZ95z3qPO4WSFiaLpxpaihG
1ls85HUjxX2zAT+5tAxALSYKZIQnAM+tgO4YEnxT+wGq8PRHp26RJ9egLOiCfaUl
l4KsDc8/v/KMZvKKtxjANvDOH6dmroVlRMqgJbTZ7EMpJB2g8pvUe7ghArgvcfoN
dLSmszU4U+XvHl1oq9j2VjoCB0jAlqlz05KCT3olJYjGspGTWmPMXGkRXxaYy9Pl
OvxTcQnTUVyU3zGPc92rf4jq0MFiU7kMp57JYfna299qxFtClijVR3Lip30ujGCT
Dlh7cgwb6jUPP91UBxj0Q8Xf7DlMpqGCA9j2WZcIYBWdG5MagYstFrf2Dr0QG1BD
l+2aMZ2ZufOVwfTOXnCM2py6AhOKOLmFF+wizkA2MpS1lGgP3DaSSmnWn7n8sybi
X6k20S0ze7MLyTmrtIWEapwdxVwSLqhx9ruxXppr0T1SejVblV64low4mYPckAos
ufbIaB/cRYBlIxmWadKZCOtJf2vq9/cmc/NLVFrnpdpHdgxtBDDmY57V1cs0tZ7+
fm1telhUbfrj5oVDy7/dHVbs9Kh5RV07x2DRr3LCEPBXcH6ArtYXGG6YIWZMlZEa
tR8uUdV47XtGO8P1rLMAhFBKaSeOcFi9llCRWXnx5LQEDPxopxQ1lLEbl2GRXs7K
T0hfVSjh293e8umirSRGgsFb9xhMq0fZXX2BRcnXdUJbhsDPzXAHfdAWoADxwRwM
iteussRCilztIXIEAtrafWrsEnfk9uF5xm5jH2QT5yvh6ToYy3gySm1hhi0u58Gt
vSpxPPEMyIo5uXagfIlwHdNwYSD0ieG/YcGA5UANaXNaALjn2A5nY7KjIIRO433c
hfbPZqY7MUBIw5J8wjIBLJOe30u7GIp3MwsHOd1GBN8yfCkvMytmErcWANW1Q80J
I7v5tCxKkbDNg4gT4zlXIwpojjrnkzIYXQCNgHx6dn0vzOTxLm4qPPK04jo+vJkX
7/LsSTCIogTJUhdkbQ9GrCLz4RVPOy4YbFtr0xhXhrbxFOrR5rJslHr/yGX6RcLH
lGo8owwLw63U2nA6dIyynMVfcWD7Jd3omq5qY7u3/NhvvZc1qXmS55S2RZ7es2Ww
xlWYeUzWzLeMzV7pC+FQo172cGK2/u5watkXoRv0XbqcuBQ3CLMk80wPUVEm7weY
jp7N+S8BSJ/hLdiv/xjQZY365c7f/R4WyrR21OHtUSwlhC9tlx7201FdXdaN4Co0
SUHZQyAJZi2pYrmD/moOjX52BrxRDFow3IBqcrRJSR0tP3iOAmAlurpvDapdGR7c
ig1keyqqsovQnJWAgfAnrHyHSjAiWHLafTqvULwbLZTb8/KaXuG+QLLqeq9gejAk
/uQMN3NMe+pVyYSCSPfGAfyxz0p1SWt4yvrpdy4oJLEpQssFr8zMdFL/2klj0UMl
nEFi7hosjBJmINmnZHGAESo0LX/Vq5UbeP6akAf2ba+4W9/Zr8zVLyk/WCC1NJpq
kfl3CwSW0twtjJuJvNKivWg2892US7T4pXGUEVGVO6T/tLVQBtIbiAGzZRjDpqT3
tqoMBkvYWJPcQZhl6xXVHFTfjFctxpvOGPGd/AweBEBPW5xsFXGKRNbJMv3PZLHg
fUSbM21K4oIu/YPiX5JyZ6N9wrjCrEyHdEo+SJBSuweL+3FcKEWxarGiXDXcOYgP
B//x6qM2VongV6hrAfwSWPLgXrNQGMTN8Np99vFA3cq8dVw/9ijR1+Lpw7lKQsEz
2+UTvrRCFZQSQjy5e3TABfApjj95an0VmEu67k7+6WK3W0pLxLCVJbJ91DpgTC7o
ONBj+mvyanhZggg1YprfoLroP7kk6+s4ll+SbSu1Mx/Lh69V0mc1rt45UjhIai/A
4f2vflp96YzcZdZApZHD9V8NlrPpGgbit/Y3rcV9fGu57KUIPkd76Oxr8CEI16O0
ZXDsLyrrhc0hAEKq0xq9ne8Nuvfp7jOcBQp9Ua7Ed48qAkUdsll3lh6BzetgEej+
sPtBX3fQtpi+FHUN9qMXuWZ4ZhhScUez6LZ2xq9lNstte2rCBbTI+mdCrp1Ex7mc
1lXqiJInksOI+0MylGPIchpIJcVDKVrP96aMUoBeuhhdPfu6YkXeksEG9n1Acw6e
msrbtHs9mslJQcvYpja9cWlAzEVxRJB4trM2p8LqqT1TIaDK5FxZNdsrPrLOMHNV
QNGTcNJHj6vA81j+KRyOAEgrZnaiUSQtGBe+Xk0FI6pH2Wyg5itw3b1/KNdrT/s/
GzgXgh2QmcfjwNrQS7003W5Vb4Mub71uws+gVvi6iHmS3shpUu9IKJFNEAhb7EHJ
rAwFOVVh44xb3AtiqE81TJKZNciCVuxWzLObEuZGDkYfZTy3LddW9N3WQoekzQDd
6Lmpr3/dF4Zu3fNqqUvV5cEUF61lrdIKw5TxJ2tzz1KTiwRmLdw/7XEQa6jfPUCd
Uek9KRsJizfPy0rANKmLyaPr1vH7QJCg0PahD9iq4086sXcjx6V7h2hxIWNK2E0U
Y7mLu0Pd4yJhezWBUyc0k7brl9xp8uF6LDyJRH0EaOoXrjAkX044icHxDLO8gDAF
CsnDqZi17MmEwUO7QAhvs5teSdo6/2XTyrUjmR41zkoD7Zb9h/VH5HXLIg7gVxy4
2XbABaBQhpkdShuuYfsaO2Jy1cIjg8XPxzxhZspHmRXM1m5rzhTmNmxkT5qOBsAY
hU1QUK1H2jwNXLpvhowV8v8X7DjG/brTbjiW0cFn7xky1qf5Y9hva7swvXvSh+pS
xSv18dYhLRpSR5Bki5wXgrcpLfaG/yFuuEWrMD7kuF5OA1Bdmnsy4jlx+kyVOdWP
ot6UOZRsPQKH6NayqRImWsFmaZsWfXIdHULNOonm+zEGTvP5XLWNyi4cdpJCRuEs
ycdi8UwFx6RPHg2povTuxDlauOF4suSQDlgu76VDJT1fEQhImDYNJy0gzK8Kw2nR
JvEN2ILNk51fcoR0z8mqqv6Qx8GQV5Oe/dDwIOqm5WyObu3LoDwWR+RyG8QXdj0W
VsZGj8PZsfRnfNbyccMfYLj2oYkLGA/TV0CgGtf0zTeMNR0RA1SCQHGgsqubWAhJ
w8OB99HG3nsTEJ5P0pEeZ8vYc/42/ONwe6yQz/4YJtp/HQSheU7HEMxBmJCSrLgF
jvbnRZAhGqETOqnzcCJt9kU/hwnw9xp7szOZsYboubokstTDuHrYYhn4xheyJum/
TvffZrqVH3Cc073UJLZyfb1IWfkIKsJZUM/g//GBCMgvQGUe35haCs3HZ4c3s7kF
N3GgCdTdzFDwRy7hEnq4c96uJJwsAHY5/pLaHXGt1Jifxoh8Fo5TBF7tOWRvdPs8
kTiwuNiu0EJbBsTB5KkHFYsdkb3dEPJIN/2r1UCU0lqRZbuEK+t2GX9OVLy2Zg7N
vsXu0bXO/aqRYfFGpvKjEpXACT1dFo+kgPwMhf5q7Ij1QxiBLMKeX2ZwH3xAZCBG
1S3QBWBLa2NjZDf3aZn7bPykwohFWgz+FVoW+g6Z9nq/HuHpz/I4XZSulvJImLDy
rly4tRB6HzqsaYxwVLHQPQWgStLCgJ5i5ZWZTepQlXAizJUK3CLN0UMi1vxsvHOG
3eMtbTZUZRluxgu5hAObzgmdOclfuZH9VuTpIdr15g5fCLB4MY5fFlWnEIAmUnQO
anvC1q3C3uMqPDNOAXUplj/DaOktthlHrwvG8Iqg6iV/51Of0PgbJbv4p4F57xip
aEY4XA1PsGaRR+WqZaF5/4c+BuCB/hckhRMryNsnIdtcvNeZi60DrW8Doji9NAdp
aivAky7ywBL+81uIIYsQ/Leyd4rIq/+jdnGV69DMA7yVVYoMLLF2gDwOccWEXmIP
sc/ZX0t1LSmoYBHBr0f62v3qX+ABp/ePU+RwODQ70W94JHHjdVXycpq1nYIQjYdy
Vrl+ZB4GyCjwEMNPKCBzu42bGqaBBLy4t8ea9QV0iMyn0lGOoljVoMhZMgZS7E1s
9+/0PIkUvhlp0XDFC1et3Lg+bbjiuZ9qtxbX2vUxPI3sGTfF0IusOX0lXOY1w7LK
FNqq1QxrcQsNQ/kYew+5fKSSXC0XOWKhnGoIvizJWa+buOzNZ/O20BtmsUPaQows
0LFCqY6gtDOmkjz/gXL01dbkBH+D1S9g3LcpuZ/rK+xS25SeqAFqHpCkAUpbv1Eh
DXkzmpN/6aztJLq0YNj9o6+pZaVd0ChE26fiZWKJYRfKsmhVyWSRId7FjkxRPZUs
SfrKkXU7NAOU+GHyAePz3gClG3D+ET2NO5s/dxMNiCScAB0ONPk4DaCht0a2CQnZ
bAiWwp9ynEhvhXsz5FfW0tYJpNYhK+Yy/cnQ/QcU0aLls3F1xItMfBaeSfTJSIkP
vX5bRg0M4Y8xrU618VF+whflC3BMpoMKK0IFP08tlGnH+Dj+w6ZlVOrR8BqBv9QD
yRSBMLTP2gNuijepGe2WgKdSm0PVrbK22q996+3mszS2M4gLEZqiqcDkYgRv2e0/
8gu+9fJrXTWEWQl8GYvgO5YIimZUpPmbMk0g6g7FAgqSwRIdDcPZMwRqdgLDHl9n
cE3pAI4T92oS93+Hct3AKdT5V/jsNws19h+m5VbpLoQOZok8Qg6UaGjH54i8QWzC
6LKMk+rPzWCA3wtftQGeRMwS+YeKQFz2kDrno8bdH2pomctid6pyB7RDb6W26hde
at0DwVMJWI4O2Cm+po2We3gQIIBtHG6SP6fgiDLtEK/kevpH48bFUTCHvuRVRCCo
z4gO0i9A9SRifJhUlCL2hIS2rYsjcmTaD0/WfsAfa1nXGsvI3Q46JYIVuU1rjyDg
u76yl77SdTVJkc5ezsLQ0aqJrHV5X1HxtdMmdyz8r/TPgrpHD6X4XEY1xCuFH2IF
Y2c6xOukxS74P3sqjYzcLuohZeHWd2we5YM+PRd+0K4vmvFRpnJu0yAsg+qlwkRF
M2oJDB4LJ1JqWyGyRN2x6VVCnb63m7LIHzm7HIpNWRFz8zslUa84yXyuugJxre4g
L4uEQHwYJada7oz3vzpWQom3jv5J1syzc8xRWm0WgcYo5f7PEc0py7lHeBm14VRv
HzgM5keoOV0d/9mMhLEjfbT2b1LQgyECt1Owr4DxkGeQouLVyplKdL+TQBBJSKhz
QY0Fv4mn9VUIR6dJ6HHSqTuJiV0rX30TH71zidjz7fDXRKo5UrrRWT+hObTsbPJS
zcjK7CxNYXNDxFCT7LEajNgRSUWCNagTSp3SnVAuaZMrynEDedvIihbz/KcPV47B
eaxxO0dsrIeoZiQOa0Le/f0nh18Jv0sR2sGMSdIkgNK/cAM/OWWFAWksM6WAEQYB
r5VLdDNPGEkYhfsq8350oc53RbCEmH0Ykavu+kFkc5vUiisOKIJi6vQKdY1h3kqh
SuaiNV7z6n4xwqiAhSO63NdpsBhScOrQSAxl+Ih4LjvdchVz+OD08tze4gxfnQNE
T60cYJA44fIrfAnYNbg88lRXa6uMfnSq7Z4xJCyq/HfkFJeyTVcVwQPseU46Utcq
7aMqCnW4Gnuwt1R4Va3ix8RNiDL91pVHxnQvzONqZIiPc6nRKYSZHLCGtiCQ85eK
1e48DhNZn4CV8gQDKuL06LlwPmYsB6+J0xASo4nMOB5Gvd2eRuiAor2Gxiu8nm1a
R/oRDtD5+I9JznEOI0RJD7sLT8QFlBzPd4ABBHTPjWfNnTHeKmI9T7v1gBXQfv2p
hAZ+qd5zoAUl9rzyvI1ohM662o5Nrzqgi4OskMffXJOGvoMQ3C+QHKGhXBN23yAM
iBKgSlRSiPs0XuNpgkSPzUyrOOS2pqHSIJySCURiLNmpS6xw18S8IG5w9xSEO+TO
5uDyGtpq/yUdlTEsTIlhA07FCh5LxOZ0prGHMl+tw8L28s1x9RBwERERGLTSJ5zx
8sRZBxK1EK3yZGdrCVgyIkY4uvyWnzjBUoBvz2K7+yy4z+c1/iRHw5D3JEIjW2Wd
3CvKX5EtMM8eAWXY76PDK7hhD6h+xOfvfdegtyqUcLR4oN16gC6hjq/mu38w6xqD
ZQQ0p0ErbDZeOdGI2+2fy3ApbHl6bJRJa9AWHKOJLxlQple9HPw95nMnBzRtwHbT
GwLonggk+PAXk3DUpL4+8SP0XET6AhqRSISSf+isXWqmoIAzBYO1XivKkxbyirbV
1Ug88neXozAaPuLmA9mZ7gyKds0XFYfT47RHkdGvC2+h1ecnbwyjoBxvWUrvJq/b
Ps8YAZhN0MaEBZPDYKwYIEhpW2hd+t3HmsxlsWY2n++KUqOuzdHsceZclleKHM4Q
EOYQH6bet5mjaVd6lXEXEUyt1CNzzZqpCMObzBpLBzFXQQawx7U95QbdoZDMWtsQ
6rnxTXqYowRF867EwQDcGkZMTlsmSNCJ96zdP3JFdhW1ZcdPHhwhMoXjI3mTC33z
+OFown7wwUr22IqZTsfenmHv0lDQQUtsSTiUlwCeoVM9Ss5YN29Ar2W52Sg5sb2a
az37sqCzWrPZpqDbokMj200+jOQxgV+CKcdSp8r/b6VYG+LJVQuvEO5ecWILn5Sz
09o0oB3ujlBiFjdAnDtPLEizOqz1kPMiiwVUEAo0LshUdwaGqugKFqQqapjvJORj
QYmkgHVINLGJQQa372/qMI3KxcCuF27wuIUOlp26hbGQk1oxhsWA2gv2iNxDC/1m
P4kUM39oiq+GENUQJbDkyH29M0GFUx/GUWzaC9rrFjM12dYQPtU8XHhiRGwHsx3T
oEMJvKzSZrVwcN+PFP6Mq66jgkgbOCYFvGqSEtuNvozudYXNYccvnswLGfbB1BE/
065NIYWP5/GwdmvLYG7/XpqiaQVT7fNhmPx4lhzmBArNjl3PCZFT6Ay8hx/xpCLz
9hx29tvQbzmKtRWwXKQQb3I7SRryEebT1hM0d+PzlledDejM8lGv+230K+jKUfoe
8pfdup1YSVKIRrmSCwUwE/vYqrYgxS0i4hVTS7UvsYdaaL/aKumvq7A8/XPOohyv
l3bQmzRAoQesn2HajszLTLPVUuRRTAeaa9WuRDFO1ebr1ffqs4Vc+ZccsS2MaP+I
NE5OcCF9k0P2SSUd1xnTJzGpL2UOzclpH4GJgehupNyJW4103Qe9Mdam38aGpMDH
745e7JARh89CJ/8aM2qR0HzcwGeHnxe7Yv2hKUSteTPQwu3UJDJPuR3+OVgaZnE8
Jc/2W7dz/mb7P+93TShXw0FLDaz/EORH49SGZP2paRUYAX3/lloAKkoxIYCLG/MN
Bzp+tvaMKDzjrwvH/CJVf8GZb8/6kKcZfRQ023O5isHsG1koI6ItSQqwpNSrOKNL
LcMcmgYVvzGcPFpcHDp3FTEqw3/blprmJGxcKC51Esk7VFzsySR+/fnJFCIOU3Mf
oxB9mUc9isLYFCtYoUcHfjij35iAHCdv5RBXODsBkh2IGnSBqr3tMLF38U5Zp4G9
K+Ts4Btof0/luNekTQnWE+0n4Dwe4iRfLpbcAgqxEWPbrFNYpXsXQOzxaRhrbPFD
MBIxYgCmOGflecTYlQCUvqEdHAFEI+rSCJml1Jpmx2iPcexqjNTH39Q8YmUdZlV0
gtJjaOHEZZ3JiFWxYOoRS+2nXV8veDeb6X6I3n6VVJ6A/PS1JLk1eSZ1b9SOlGd1
LQQkA5V4S5gAut6HpfX8lYLW2j7248Vudz9Ps5V/fdF1e9icStwcxGSgjSumA0vB
h2wKie2W/mSD19jwj2Inn+XhhYCoRClJIcf+TDP6p0zBCsW/1mGetxi0I5vMbBlY
6a21YcpGH8twrelObqfndCAzbKSdiR9VGOSKWW9E8FWbEaoN3YxjTJdioYuWMKB0
51SMk0Cd5X8/1uets0CzQSEjxCYqFFjR0MZb4sQoyMSp2IUaALaf+4Np2jC47X7I
UIKJ4Y7IUbXpquAN5uZ91dlRmra9o9Y6FfFc16rvV2OKY5sT/zlIhrR/jBijHmaI
7uVxk3TD+tZOrmPX3cWCgivp7/Cq8MnyekQgaUSLrySvmIFYsyv6M0D21E/55LJK
6PMabf73zND8hb3PrvfNh9UhnKWwbJ08z2ZE7nIPmfuvzMhpEqkja79UD8xnt4Ob
TqpE6ODEhlgbmhgeuUeIljeKFoTBvz74p9E815Xi8QznehhbyyDwIbKDodhHlumK
oFlYwoaWRDiDARQzFDUifVnwuwiat013RCpmiOG1EEcvDhHqZbMulLrcToeES/gW
odJw+z39GtDvdboTEBTqhaOnQkh2EbyRzRgaCL3PS/8QHPXkpfHLs+zBtJ2kRhxx
sKpx9aEP8FjpKORaU52U6b+wPgFFC3J66o5RDCF2oAfbF7bgD0uec1yzgOOuHrnz
qbivaXmC03EOYQxJ6s4yJVlMgPCiUJ+G71L5L9+uuNuKVEfBC2f8xuvbSepGa7gd
USXMcrD/W62b4WjusmjpJ+ACi20sdBdmJLUV+JfTHVAs/Kkwwxm3BylL8stRYi47
YuWr5593YxxxVdWBtgCrwzafsmnhiIgwH4kYaY41K7DNqGJUQfex8CzBAEbVESv2
/sBQsPH5oz69Gmob+MJxVnrjY1JUkqVqncZM/BN3n8dZDHp5vHD0XjNabjOVa8Ov
g7gzcbaqAFV1kXQDL4+vedocwYj3Qj9mahq6lBrJlvUWDVmX8dGd5TsQXJe+mX6i
k2Este2xhypbXQB+G+xU26eRXWVLLmOXYpTYxR273CBsN9W0yPmRV//Gt+SIZsCN
pSwq30DvDTgeUUFzWGiUBInyDVucrB2/DgeAqAPmSfy/oXlrZHcEDlrvzqYK/rb0
6yPXKAYglCtiTEDusIHkpLt/ZNaJN+TV0iTlYxWHtGZ4i88HRDhKqE+v6kRkz7DS
6XcEdlsM8JwlIi0xBc8tUmgXUEVrAs+eO3wYKStd1WGfJxrGGNunUr7Uu1yy6b6R
tuZw1zAqgxJXOMAovSmribEqDmd/JryS+OiBE0OuuQ9zw9jz+Wu/24DRhXrUnsnd
ZtDjBDC/h650w+24WrNfBDCZdMAuqtJwz+5u0fbttQur4pSuLpCEnKQVVGAK4eyb
AfesklBInRu85FIrL/aKKh3dBGDCuxKQF4cofFKwIQvSDRI/25pX42xDlTsPwbVn
5RIz/GxDWL6Zq9Dyt1S5TWG7l+qo3I8R86uiPd6zBRahJ5owF/YNPIktoTzsU5Hh
pe3PX5sO21zZcNvfr8jmZbri1yuFMhqa2mfVtUR8TbL0HvDvqUg9cOGt/MJCYwPl
M+Fkf/KAptNf7HsYp6YfeX8GaRZoBoOFmdtcrW6lPhQejiKsnDBzNfo/WJV9yFAK
VNMgnjXWOTvuxR1l24zYtxuaAWRfDKcqojixAER1HrsAp9vgL8IJZuJf45uDkaYT
IOKyFmscOnZt1dfY9dcwAI5asfoPa194mn7rfQEoxB87fNzDOzLRxpApDUH8DjDL
kr0aRoXW5IjJv1XEe/TnBkAuxBeN48ERIdVxDVcOr/tvrOBBmHgfGCFQgmoPiYEU
ng85nBpkKmxrWTgmKJKUGGwuqcVEJSACeuTQ68n1IVfQ3anRYQwEIFizySPTvyYH
S40PA5UTPihpjUBzNTm2yl+EyxlWe/i636Hs5X6NfyLTQyuvxP/DMBVsdn3XGNe4
5g77AACCAN46V3Urrf6kLX8f7d/YXUBz6B3iuz3u0D5PUJQpxaq8cOv1Q5007DPZ
Bd9yH3peEKjHdj04+y+d7z3IgWc2LSkyJtGtjYezAMNMdESsYU+ZwTkkT5rYqeYD
x4YQqhGTl343dMCqLuIN8TJ7MG+ZrDyXWpR71W6mv7o1kIL4cknOEk2+KGOvqd6P
LTt6hUrfg6kqYpzAutyk+iX7ybR6YkIbtC12yMhbhswNnZYtIFo0rffw9brz0LLL
wZ/5pYoROnkuFC3DdgUthHMeoDeCZwxQWVOkl54cdETQkni8OiJjCea5yAA23Kyq
1qXU9WXcz9LxltQo0rX1aylhCJvWKzysLsAQ3hCYSxsTDS4V8Rha9C6F5yYJL4r8
jM2YAGX32NMqmvNenEXiyMx9v4uuX4kbF7E+fmzQSI91F7P4ehbUjjFT5S0wKi64
QfBiAG54frSxkpPUdvgrL5zSX1Ox+JP2wXqA4fiIe+qxM4fpEvc2CzRYbUxi/28m
0oXak0o8PwoxNgj5Q/bO2L9sFF8W0OF8gstzj71ExY/KmRI7TGNe7A6+Kox08DOO
nP7svWreLGm7YJc+xIu8PD369ul4WqZqTcczZQ/qupxhxiorfKjK7Rdx8lco0b+J
PZ0+w1YD+ntFtX66jD6Bk8nfw48Qqp4ifKMSmuANvKpyMHFQ5JdWGwOU42zweRPn
QAGpcLe09a5mbAIyEvudnDso2r1udm4YNsn+Rql3Jzu9YUbGPHaiVsq1ha6XSvvM
6/n2MZ8zbjUR6IrsmzKb7q/CzOOvcFdSitDYkzWXgF90fo8D8jf0Sq7RbbDO8jgV
y1VjiNIVWOlgLNqq5C4QoUD7TaCUJxjRsYh1XDXMm1Smry+GAHU+17q79h2iSstI
/Xsfy/5pQiVGZZzFt0UAHvlNDEfQDPRDFAp2HCpINUYx/MIVSwyJlJqKiAKEssGe
ZRxCahTwI2dfLXyIf7N5Ia8hG2VfJbaETv+NuRSzLN2q6Dw9hWDrSBQivX0qO+DT
D4cyKaHIccvQSGV3X1tlFTRZMyeIjeYBCsVdNv5L2byTlhYl0iiwNx4kKlapwMBU
u4E7IwqeET0bFAFgWqVTSYxkQqpj0yk3xQxO5OSWl8imHdt1BJZqcb7LHC36lwl8
mrK/kULBdH4o6sNM33rKT496mkTG9M8nQQaSfjJIgXBoIW2+W2jxqvhkQPMBSBZC
QkxIIopvrwhdf2aJmIHt0ox9bCkcwCKLvnkhhurxVUcdlGqFXU2A8CfoxGS5r0Lt
7JF43d6EMJzXOnsC0vnBCw3ydE1RO5iZs0oYinfLgmEIb0OJwvTze/RN06SPGhpp
eHmWJ5TuefoCKwNyE0kNAFBC/ZO2hYgiXL+dR41Zna6SHxTb0mgNPRwDhwa1iB7x
y57A82ga18uB6mvWcNPSCtGCc86QLUBmEnFoEm5Sp6ZGewn+r3Z2K/Yya/YXkwi3
t6Fu/vTOYlsN8eZAt6tiZSRFlSptugQKVerTJYfDhznYZkzW0Qpaf/tl+gVmDcpk
JqsMKg8VAGQBvModh0YFIrBv8vLmVCIp2uMK7VUyTdtVD/72CN2gvdSBUCjzQQCo
4LT5gDAourhOJ0/RQ6ZvQxfP7TOO7oMMbL8VR85P5J/SAEl2IbVK2EQCN2Y0JUmU
9cE4xrIYuXiFAqfBdD0XMODEgQl3XxzXKJP/sV1fPQxd0uIpc2/toVr4ov8HKeAA
swMiYT875QwKrUP/Gpp9ld5o8QgcpCe4vcSHf3ybcl3VV3ToMYkRjpLrIX3iKuoI
T1kn4qZTtPpqauyTqB6+D0EiYjuIQWciA7umCl+1OZv/3ImI85Ntdtv/laaPwWho
NvBuDU++mplTfrMwvkvoe324GVfZIakLuqmymX48Z2kEC5mJMGuYwVWNnLGxJKYI
7YiYZ7h8AOUCplS6OaJWZ6Vx4EJNavl5hr7y3abcFd48JAifrLlAUGKXPDyterI3
HIJDi55UmRiHqfsTTEaB0cJsk21xZrFMzkUM2dgNIhYGqvzXIbvNCzTYmQVCJxBd
85MNRRM/ULDsEU9/o47zbe3E/G7G6q9jyOrDwS1Hl+avpQT0kijElwjOBO9CSTpX
nmmorvt7xF+GpMyL67irbVy3Iip+XsLfLvIOMHsUgFF8/Z7DgGeJl7TKFp1TqoXs
yYGRvLcs2Um3xGc/GlYQm+fTs7jW7o3jdwie9LYJwjPTvakccszyyQG1LOZYLkZs
GIhKhgXgYdixEXI79rzOuPWMqlTW+IlxbnETkO0/TXnmcRjjJewaM82ab7vY2MG4
B+blWfI0Y5r3xmzUvCpT5TYwZNZ4I/eFcIMhFglU2UIkvHVgIatq8qTvnMzpz4jW
7vi7qlZJldXddkQpsuRM9DII7Hnn8R6z5NOXB8yZnol2t8RjQcblIUrEwNGln2il
id/WBXEVdL0Jl9Uf2OEXrgoZm/rv47+oTJCa2Zf8J1H69hdD/t5teBZ2ykM9UJ0o
1jbkjwmUYfnJU/AaHXAua1+5f29K5QNZ4oqZ7NxEQvqpFjUa87WnRF6jMLy0J2pA
mZMnU5CEg/uDWHYreSA9fNkuKaAwyP6YAhjfHpTz0Xkmq+yxX7h5Cg6REadE3yM5
pCw2NwptzqdyjtCzVWbaNU1SXvgBS/uD4arq0VovxDjAfWrBr2kH2ajyTxUE/vhM
/g1V8vQX+rBSyaM5n1XvUJ4LlaiStUrdVIjgD+fw+iyfwN7lksPnI1Wf42qKp+4J
8HlwhMCLXfPplAQMNVtDUXbvkUZWo4VFmk5o0NNZiKkNAdcKxoux466b3nkBSgvW
NijRtMHt8JXMfhRcRGuOouu6L15a/qcqysHCmvEBc+iM8XskTyH425vXl8KFXJzD
vgoFDTrEJ0u/oXuCUttM6XiOTwvYHl/2t+EtkR1UJKkm1OWeVc1IuSkUW2fMNKrD
OL6mlcwE2wfMvO79L8A53NHKUPEWmrBjKogZOBVJEsHVXtgdtSEu31wxz5JRU9Za
ZZq+uMqvdp5/49/FsPbE+/J8wDK/y5fp/WY2hP1w+73fT+vppaIPl+WrgzzN0Whe
+/lXjbHHKHYk496AFbv+AvNV4Hpzl0SFQ9Iry+c9kRcgRz3iYzL3f5V3la4dYWtq
GQ+ZEXhMd8fD+1w6vGGvhNqDp+67e9+SNzuc2t9DdK9cGnxpAU7sCWbF4Pq1aaJ5
pvSKiYp2WaruXL6pMtuKQryzd6UefoDVti9dbiS9VySkP/T2x3qpS+qe1s2hXXaZ
jmUAua0l+iT522fCfOU2dfEP8+gR/oIZLXGRq+4VJ208/YD/bVrd/QHlStGxQz9w
gbBJ+9Lm6Oykgov+4wKHWdgv200GkqkssqyPb11cpJWcHmBKfWMiTp/HrbHhfWQu
GjE76w77UUni9TcUgzHGNxuZFtNtrTQsCk7TVsDAso4N7nC1EBWStnAYGi19Hyf5
cF0nvah94OMMwRkzOWsqOCshtnxH8+lof/hL1OBUL/2DCL0FXExpy7JJOuHX+EMf
gkWJPJR2ta/ciLxVPsKNjJp5q4FK6fNKeTbZieo+h+E1k0DmGyPnEC6S3zr9miyF
Ldb7YVk/2uswg9FKISyMAq9b5qprmXKJcVXW4EBUo5HeDk9h6z8Wj/SCM+ethcMx
sQZdRrkDh2EBghJSOHX3dzJZyIg9YlL6U8Wht5j/153k97gYrvRkDcBCGqmKQvLi
ESTrb5VVyUIJjonbx/uhA4CYIln/oCNzeuO5vYrBVVwJMLxb9javuq0TXKBo/g+k
Xx2J+jOkb43e1RfP1CTRwJlm+5R25A/5DnOv3RaXGmR2ElldJ/5hZyXLbEDhh/Br
maJ9/FhDy/vJ2j9Lxf+WbXZ7XdxqZW98gETW7tZGBCa4ecAB74b71XCLD4198Bn6
ZwtX1EUxd25gW90rJSeNXOWj4k9JAmqLb/L0y7UAp7SoXEeKnmq1TWniwWR5WuS6
/dAL0w43wznJ/VyqF0IWyxKlGpD0bqHqXT+q99kC4hcYlzPTTxquzo0NZSngdJSp
yECUNFOVkupjABBWlYG8B8fwhMuIyEC4eZx8+GeLMLbe49cA/fRtfViufQbnPsrk
1XhbLKKKgz6p4pq2RADtNcdbS9dgru4hXKeKqE+1c4/XrE4J75zDClq6bjybSrKb
rLCnn5MoC6tFwA3WaHFXEn9wLikkfxw1aznOKFKH7sOn6tFXY98tuc45J1f4KUUe
K3GEaCZUEjfrmNtcSbIET/08WeB2ysn8qL76kAYf2tQh3dkXA92jF9pDVDR2Odsm
sQnjvfS4ri49TRZs33ogrUg1/BSILd5iiw9UoUw0ncALcueemdLQIEoFfmx2dpfb
GdTDVo0cvXJbaKgVgQmW7uG+piEjeG5pI0gbTVu3Twbe644U/YdgQ/IYuai+9ERs
LuffnpTWKSF2Hfxc9ae5Eh2mH5pIcFj288ucmerUfVSXyx+nTHCraAnpeAAQVEoB
5wpnb7Ipcur1JXxlqj0jjkDbltWLxY0EX/C877uuGWdZMi8BmcmPfYrq4c4LfzWw
mrHxO4DbePbokuZWigvkbFUpEYw20urhATuNu/7FxY4CO4QAgcS5WF0nih3PHjTK
Gox+JrgsZvZ6dFYX6l8x9jvRH3QCApjzb/7pHUq/e+kV3H34d8msaKJyaDBU2fGP
5E6TjtEoA3O1vJdGyvJUx/r0jIh8C7s56dZ7/pgb+kXoJq6ESlYf6kXBT7OWdI20
aB23LJpROENQXNBE05l1oi3+dVIIJq2dyEb4mU8Ygf5ceXR/xaf8ndecti45aR11
FEbOMZMBF5Za6Y8502E+yaZrMTDdIAVlFRxwRE4p6Ga3tewxDx7uH5FDa/0oYicj
hgTZamv/JniTl6ee9OsChSdhM4KrOtnK3iNnKHna5qRPGCnOQMTY/I3MXnlUGJPp
NqvpTAg0TyFRdUamEc3YL21D9DiZGL0IX6QLum/Ow2VrI77gw+LfnuZ+4JKEqtFn
UGxyS1jzSKsWzy3m2A51vDHvJCbLIoYl2NrF9clVJ3RmoQwwU2rPY/EOhVzbMKMq
V9l1PR2LPOQTeCj8rreAhhakfFpCnSwTIc6FkbgyYVOBaaQcM35Fo+VlgZDd6gfa
pbFQHdDxIuTovmQeGxjUQLlafPVw0KYswopaYLrFn3Y6rion8WK3zMoCgek+GpQV
CP1DktUYUjcJ9k0sQ6FdYlkt30lDWkV/MU5XwnzVFjTXAw/bgpF8wlkzfIZBZlFL
0at//2/LHtZNHh4Q3tZOU1aJZFwOBg0OOGvYUwj4JhZEzo8mOvJXD61IsnxmilnK
81pfeJz6bqMCLDgQh1SJ+G864HXAn07pT5Da24wetIOhGhTAOTrPvlhzSC5FoOu5
OmorMVvg34YRdXs/y+zlGTdgJH1cYQnIy7w/9DUBg1gGwzNPSyRPQWCRrdnQxFrt
1NwoHfp5nVqYJGCR6YsyOdSUMU/qp5NRus/NrKeLhwWr/La79oYr2x9d9lgcuoD5
oaLF/sVQenOJrVDOv+YRF0X2WXFeSQuQeuPRUMwccM/ocs5Nnz4wwWVk9RDuWy8m
46KxUscQRwMwhwgg6lozmqCEqnFGCFqu68/NdNr6K6Rggg6GXLI5JJPrqO3Th5YN
ZOEDQuGPZeIIoqXfh20GPjc/g3od/zhob5lrmAw36z60Mx2LgDJ4oR59aefCpJQ8
vfQZyQw78Zzu/yZHA5cWATN5ahdnuqmoaXH88KUUpsJgIZgl1qUqpWxuVs8enF/R
Nafk15b/IBn9ANMKOM5Lc6uy0XzTHevdadyhEJV1S9rStal0YTXsTER+H8Tnc28r
I52HCP4iswhLvpghz39iVHlu3twLK3QNdajOBzqK4xNyCWLAJh+q27ntSciHa6hn
qUsMcPWq1fJOrIf/jsGKHy+5DJnum5l3mw0EkId129saufM6425L2SNdPdf6Z+2m
zdHaWA2X9bdYCabR/6rSWCX5ZQwYutsCy0DsJBFBPu7ywLXOZ9zWwl5Wl5NpG31C
4Hd4ur7Fn4aa/UjX/s121wDDbVIJiy38iDPYifBNGaVwjgBTIoxX3M4ErYznqhSg
OWN25voZ2XMwHg8lglu2iknA4pMFVE9EmQy8zgoyEOzR3Cga4bPqEAKay7bmJNPz
UTo+zeYShPAn5SjovLIy6ldLb6/y+L+pqLM5NLkKx4HGpXL2Yuc/dqeFp9Dmy89f
JFddCL0k/A1WgLqg++s6LRZLjrzxEJrf58rnpVvbxFlHP88Z2dmwk1hwcN9FxTUm
RsIX1NR+lQS22yC5EwyFC90ayv3oHm97x0Rh0YB0EkOszXYpnFz+X5y9qov1480K
ujWFGo1IOJxQs8A4gU6E/dgwJflSBBtppEeaELeVGmq/9VCzcPnnzCvHRNBoT3o3
8fSytPowkqLB6j/MqSLcYwy5GWU+fYCdX2K4MAqwf/w1UBpLaXJmRGciPVHMXXyI
fezFNiMsQRi/piStcydNYCWGe+7UTadaESEo02PeeCwwYlxiDznNR6fQe1znUPao
CLSoikgO56ydK/xKHa/DOJG14LOjCa2tlFi3zuN9KGe+sd7NSsNguXpMmhPEgnEH
VBHQiSKBse1gurFUxsf6gI+T9Cc5FLdJ8gJrztdLK6mMEzv6Mk8m5ScdsCT8ABHc
wzgT9TVi05argdbRNN968+l1WTjeyQvw5t6GouFlYX3lBiT2HYuweDva711fLVYC
u4YrLRIGEbyS6vbvwWk84NsSJumj92jx4wqk3W31+dqks4b7KmOmCdnzXQVWXsoZ
KB4qnOBy6KLDjurHn6Jg6U9pg+AxSusJZ8s97fyPxxIMXfBJPKUoMM3sme2WWPA5
g/pyTZvKo+YvOSNbG9B4Oqy58h0+X+SzeIFVTg5DuQkGRrAwQFrtaex/incNXglE
HpGs3lf3oRhWX49jwnGMvcvd0rps+QZBtZLyGEuCPhbYgdInuMnBvsd4kjGFCkWB
hepr5PUePY3ZEe/98yDlnaxjkKNnmFyoFqhHuSLkAuynLZAhpnuB/jBsOQuwIu1f
at/FN3VOWvI0wK1yX0VO/yWgPVjULZ8uP63nZJ1JzW4NDnawivaVwHF1Xb/+hST0
xlBCCMZktj6Liv6uQXaby8rPKthdB0f6c+RvrdGAzXldIoZdwSdp8DDyXvkecL6r
NtRwt2wXeoZEPTP4kWAGskXX6bspY1v5aTog80hdhrgjL2fThikAuDndbz3PwkGb
9ummZMtSlZHr9c4mjymm7hzauKD8bD3a4mAWMvv15EN4MgrkvmjTjIe2EpWAl+/F
eEic15mU7p2w+FXjgbDkYIDgTr1IKg9OKZjJXmOK6RPoU0qJ8jVRrealKCtSqOMG
rOCBRa7C922iKngr0II5A/yri2zjtYJkxLTJ+jM632Q0FUHtPelyx50Ear0uPRP7
at+UBkqJawXTKxePSMowZ9JxWuADtFOAqxzWx+GXealauw1xJbNvewuPD3Oycw6Y
PGTtOVkcbihTnGnRn7WizlwX26w+/bbFQNWw5ZAYE6kNRuvCLnmWkj3PkgPo8fMq
/Ho5prfxRLDHWGDe1YYYtr3qzBftPR8fwW3CkQ6WBzNpZfbwT6j3BuqmPlyCynCx
ryDk7tmuuyiebqlf4akj1+rGEyJkuS6VqXjLQP2OXf84MKlsEDG2+dS4ItXwFKkI
nyIb4EnoJlpj+xgrvPq5LeYDjr06a9IHajZMskcbqMutgoGtit95OfNqc1tsy5cB
0TqMBGqhuRTynP5tfZbqDlSg1vJ8ZS09ADs/vq4D0L+YfFYxn5g0059vYuJAKwU1
Ad1ZHmVZp1cqcjf1Cc5VMdcTcjwRk47ZqvCRav4Ms3IkKCYDzTt+Y5dOCbTp9QJR
KEqmmHWrcMxAdkGB27eMdK8iR/rJvVmjwH1v+dmww+PEbd2qxm3HrjVuqwvEQ5AS
iQjlSQtrEN2/tYvPYL3mq6sqBc1UmFFRSPeMKlrqHxYZ/iT/D5vKOzlF4WZV8TSK
vJfySRhRiX9yg/HgqLQvaTfoj9/FZDYFoPMYMGSdj4+3VXlpKSqoG2lsqcmIcdMk
afPy19UJeBDY2k5pcxhQa3CcRxRr2grW8eosQlJAIWZNxt+qev4ereoceLS1vqSV
Njnqrrr9z0JLshwbU0XlWErlBvY+WQMsBTOKFN6sJsWakdOJmEGpzR6dcpGBwddL
5ykSJGxigfsep356VyX/9jf5jmtsQeBBwn3QOIgYHR9FTll/91VGiC69emSZd61g
79fyWtTFSe8Ef6keZ1SHLHT2WJBca3ONl1/LSAvRzpeXvSnLRcOtzzrBPO7/Fcnv
T9aRbkpMFHvA93OpjeulbmyzycfU+39E1bc8tA8nGOSgHp4TKzUkIz96k2tR+asz
lyfk1VC1/r8fZpGEaMTTtDor9TUpf1nZWrXRNZvjpaUplXgRBVIOYQU8DY/IuEi4
rf2466yxYh82kbXmDlP3tC7TXs3F7vvfUIEQo9dg7k0xW3wHCKCO7c8T1NaQ6f6r
bNrA02XV5bnQM1YUHhr8q74ry9Ddd1qYfbI66yZCkGvdknjwiJ5gvceWbe62Mbkr
lh8jpJ4lQ5BxJu18eUQrbMALbIFi0AwTJfTOXinjTm+9a5Oz/B7P0Mih61YJSGT4
BsVBuIRTsMKSViqPBNNt5ax/BzvpQwV3FRYGtz3XS11/+CTfAV++OWumUHBWsHyL
bENCq9AoPiYAL4t94RTi1+DD1Gw/6oZpKN9eLmoQ/JQx6Zy2Whp62tvmKwC1yR2m
I+RX6M7AO8429A0SrVHiF4S/lR+jkiSWxNB1SWe9SJ6MKtKc2giaep6cu5akd69K
WGL+scOVNwJAYaF97WIt3OB4QmWN0hpNHnl2qJIwXoTQ6OBEC34v2XTZEbO6nneo
VuhKphZFJ1sJFrE4RRo02HBNP0kfbfRZhzCAcYrET44GDEYULQJvkR6XiRR/kY7b
/EalI7ykFqDYaWRkv06QSJmC45dNEvd6QWhJCFwJx/TuczVInQxHDbHzF2qFLKXy
tmvJeNaYlnkqe87H6pY36ZTEfa21poGb++cKF5q4V8fPfZWAEtj8B5gkvG6BS8Eg
kPUReFBq1Y1U5M6BbbgevkfQS+IufMXkhHuP8rYljpV94KPOVsyHDqEIzjSQFvNk
JQ5UcayUvUAYNu/yJY91ELvuuyzDPbejJSaxLwCuWqJssQXtalww2LW24heUKgRQ
EkQz79FRgbG24c5QG2jWspArbrDiDqfy9HHleFDFMgIiXq5f4s7pzWAQJqKH1AUi
AKE4FiCH8KbSQy5gfja5XvvNTWs1k1A+kddT4lN+hIsAc3y4kKLX0krHE0XuJxwc
O088nEmIS+iBdwMm58LrsPMCq3hhYNO4F/ZH+d8wqaPAEKcoew0fekPFpRILh+EA
ZpgJPKHaKJaa5+3uszumMZA3ijrYIZWCwSpgCw34Wb6Wxe8PTPaj22OGyGmn5qDb
UkhobpMy0D4EAW77kBzkTNNJfnDs8Z0KkO23UthGP/i2iYPuodCfAdkACKtYFevQ
DSEiJZ1OebVfPyyU6fcGXH3ITNEe791eb5dVv/0av/dNQiKGJYCNktQ02OXHR/yQ
6b2Eiba/uSPOgjntJJOv1q7me+JfDeQe75iNIFaH13OJDbONOKG8UdA4KoZ4gGYr
JqFNVzaRSyM+ovphnbOh4m1yc5cfMKeQQDIkT8tW2MVYTKryez6SGrd7wwS084Ip
yqSJTxYT4zJ8Lns6kOQPHGcWZjq7Y3TjW/TWAw/0pdiacJkWnwVnV48ArmSkmTzP
Q1myHxK2hi9KjDwIY3lMkYtXffw5RtIKR8kk3clmWjOLMQTnG0jAHHXZ7tAFdaG+
1gBMkO/p7ZC1IPwv7lqcspMzHcQW/Z4kA76a+V1MpNbMXU9oln2vdwsIom4fKkyA
bBs6o+NSHoUdxVF9rm+Vbyq1TcT+Kpep980wPrSsP4a5yXDS/osGVUHhpr+ao+My
GMyHKT9gqcyKnqc+Ejm3AQNwHWvTHLXFXFcLFKi/Yp3U4ryz+Blom273ixKTDLiz
IsWcKjVmiuiziNQjirgdQQ5hto3v3jFL4mYRTZ8Of0Nj6HNxOGleyPs5+J9nj+5m
qjILrX+kn+KEtog+yCBTPHiXIE7e908oYt+Y3bsmmco6ioCiHOWQ0a4G1E3G/n17
M8Edo6aislrsE5bp6c3TcpSQO/fb09BRLYdDsMB/dP3jAVwkePWPACX/d9m5JPNQ
OrBxNg6LrKWbqYG9TBtPquCJSITROb0uNfpFlmo3aZJQsDGMPWnMR3xVVgA94RO6
+0cfQC3tQk8Ekiz4uRCPGu2pDN6tqTgSvOXvM2KkMd9HECpO7/6j1Ucm+3thGbub
Gc6s7C2g8Ic3FDE9RJ22uhF3xtXCqi1Wj8F/DKK8/ojz7BzqNJEIf4qIL4ZIJsq7
/OYkCQVRMGKGxJgqJ5tqP5RnjZIBacltR3X8NOTBisteiIjJtbLEK9hPH/1W/hI9
R34NXlrEZfo8ucbgO5VcVoSKd2movaQg5aksCrgRNZvprXfQpjCHhBbtHkTJTXGr
CuOSNR9cCsZszd/yoVqXuqmFPEvnS7qdbGPHlJBSbhwjtXeMDINUCVPWVqMlVOz2
GFW4kKWL3aAHUJwBMD7jT/jkRtS6MW5VI3PuPwzIamd8+QLtQ5xf3Wg2/cMcN/m6
ZG46v42CIGeynWZwJsF2oEbiDlsER9r+ZpghcytEO1bshplGs6IAUbBjwuIksIHo
WdAMAqcGF/BjCg1DMmFKb9lE3yjlTffZ4+L0huaVQxdQoVvx1A36K7+op1LHaRQJ
mtSFUJPSCGbNHTrn2RMg96bjnDQTYU0Y8DQ6XUjzOFJXziMsAQCtmr3G5FutQsrb
1jN4flgqX4i8IqNF+J78dybuNpZ+lLuRyMbJAKWqI1j9Qhe4o7fPLSYwNgg2q0F+
+ZDzYr0WLdT2YBq9BAwh/upH3PnI2bRtVtu48/Kr2q8Sg9rHSSDA2QUJ0AFeYS8o
8fikJj3aJ9Mc+IfoXEjR5C9+2Z51YtwxGNAGOiVzMDDbJwkqZjxG68lq4I2Y+xom
lhqrws0FwlkGwJckjxQ3HAUmAslFCn3zPOaqGc5s2CvRXgQMbUJMD6oDOdBGcFtS
wVLFpqrj/7Gwwt++YdFf5EqLRA+v1QHU+NZ1VPcxC0uYC8NoFpjkLo8jt2nwkwm2
8mqh9EATcaAZHZQDN0RKicXUIye+XmLMYRHsilhXTZprcJDSOHnQ9FyV5By5E9oh
zJApshGRkoaQURrAihtypPrmK4jwIurBgjnqmENE2UBExtxThUCMmwQrlP42CM8M
2Kvkv8ilsCIgGJtri52QcIHCLEgDvK6u6rMmkBySjyKk/TJ5O/sNjgEWd52HF31l
Hivk4temYpKXXxHPV+yzTmPpASSujxUS0y1iu+/Lww0owsHjdEwNmJcE1GA9HPdw
R0IAfR+M5h/98h5acdsW+A3pLk4wODhLuH8KVh+E2qPmotTIw3nf4OsVE+gHbOaU
89ewjCDXTStXBmgi3rhYUw+EjbIApYYqu56nLwJsOdVZCoHnOLIN+o2QZ2pnM9tS
6tl4HGEUb9tqGPHlkAzVOjAjXx3P1Frw5c2aFEXaXpuqkd9jnkfRHNVOeXT5izFI
ubDUS97pK7wBgFYJKBUVAk1M9AVHHLTdtU4r3TKRIkFSAncRTkVreY3CBcRs1CI8
rvgGg51njeO49aSx5vKmn/0lH1V+3XQixyLuQ+m+71EQBRUOwO8bJdDlW15/ILbg
AstzCPZzeb/DZ1HxUnPzDdBcUGijujK5VFMJNqRWGOwz0fSrPTA5Zoc3wizmyMLX
lh5IUcfBzvWw5y0eKvc0FMz6ozT1rlJHdSDDy4zzCOfGzT88Hlp1JwFJTOHEuHQh
D1F4KdJaa51GrwdQHjFNlRcjmVCZtCRU6HPcZcA5zLkKaU/pSae0eOVTjqJGj6ox
g3xLkc90mB5ZQHA2o74ddHUsteUx4x7CDkoz+EcbdZEyTsHCj/OaiQ0ari8St3Sp
+/U11AQdCLgvxNB2i4L4z0XPfqkbILvB051JRAUXdtfFF0CGuIt+tJrNIjZDk70U
27X92gc9NVI0ochKFW3jd/2FN8uOJFE9VzivMvYcHnxTmDMOfstUii7OjUAfwqRG
qdYaIdZd6wh10u3ECVjGj+1AwZgdVJvvmA/HDGApDRaJdTonXF6YtQJSYa6IN4H8
dka66yiJIAQILPfcke3Re0dznIKgWkmbK9W6awDX4OpMc0lO5xlmTyntWcbznIJs
Yy0NhtlIzNdphDiUnqltIuycoo5etzkpFYI5pBx7sK99RHmyA//IvfBP7HFDupS8
pPK60XFbb9sItMElLhGkF3cfFiiZ2QJqn8hBScSI1I+LIHHaIQTjXgfWV1yiGSlz
lZR+Ruh4Dl5HhIMV9Z/DtvO0GiayEy+FB4Ej4BjBM92H/YBjc+b9gsU8jjmu/G5z
MYb/2HhOyJON1dPKtDdO+aTsGn6M0ROOakK9Ycvm3SmItyM48jCBuobJuNTPc1uA
zVPHWYtDwNZHXM7YlIimWfnx+pn+lOHM2aQKW2SSFEpsmLeKUzXWm7V/nWDZCV8/
ciy1t9mKkxR7JBY92gKRSD7aGdtU6TItyDEBUGv7IK+fwStY3WfGARGfkOD0jfWd
yv0HtM9PY4nwwnPrORHvPeeS61FP05Z8RDVoZ68cUaY1N5MZX6hp1n0KKK7m6qZm
RzNu5x3kvSsGRTkNAV1F6Y2FTOSICUcqfJLLQ1oM2coGM5v/Ws6Z+Xnd490Aehb9
Zwn7eAjMY6q0JbcUVSHCk7QiByydhBeNxIBuqFhHTkl3DKJ1/VVaffRZhb1Uj1LJ
E2djvY6ITuiiNCpz9D3YbdONk+hPDbwJKeQpf4BUqSPUe7HbkDdOsJHqaggtTRDk
/vpcWQN1a9Aph20TqF76B47CXfI85FeWAeNjpM6wZGHgRYZNGHJz4jcVhLvYC1pk
pN3OieCs850+Qx+Pa+KMb0lfOAfstLTzDrluTLU4WhYiSVld9pVPPlIMzBhwR1MH
ghEtocExwg9eyuT63OY7qY9a7wMr5Z20MCpNwvmynx8upyp03bcuB5cR8yIAQfJy
vkVW792GDR3KaAAMhpO+LV0xFn7HHmeFvJ3650yAJdGE9agVEWvkUUoCNUFCNE8X
cjtLsBlxo6P8ZyRJrzPQmazIQ7n7bDUerdilFdZDtjkMmidkMpHKLoDlGZyNnk11
ssGLeSQdigLQhv9j7NpPuoApoArnUrJR1A9/7HY02x0rRKmtdC7PR1zTpPZEhgLe
fBYSLIYcjf11APm7ab/7B+NqFJ28YNShaiKmU0a4mElmNRcxvBnaSPMstGDIW5cL
d3//MlQpEd8EycCsN4tKwSwccEEoeR6Dzf5HUHXL8vWkS8pWJpJTXJ6bMcNSTdcX
n5XC8dlCWvUTMkdKTJlqMHkhbiMVOPFr8BpoIco58S9YKMTORHYASVpXzbGBeZx3
rT7mP+sgRqvTA/38jsTpGF+zQ5k2vG/Z4BM5hX270mB2OPJufzLmOFLpkCKbWGQO
xcKGfne2/eBZqZXqS1YEJgame5FYb4T6bmCh+GtcinJAUVcQmRpWZCLDRtY0RUsb
d1uSAkI6+3w/akOuiSnahfP6UQwfVaWbshnu7FgDS6w2lRDTAQjjBDG+zSu3pIuj
8dvecwyK8BpdT9rjX2vSCIbPATeMDTbHSuaa1GfMyaybziVWkOb7Yrjz20Gy0JWW
MZ9NUNbgdY+XotxJelE5IPOo0dKOU/IWrfWrh8MAahxS4Byz/lZJjr5y66s3E9Ho
huRd4QeiLgQfHCJ0zlQCVxoKpFgQNf0c37+TyUO5QfD4nX1AjJtCvW3iZJhEMASy
eb4KcyW5Br6NgyyLQZ0QgKUttkIrYiXk6pJH9w56G13oXGLZJNAo66tAeMbjcn/z
x2TuZwPLQwWsVbfDGCDngV0owLzfz0e+1iPNQsyIvkpwbgnL3jEj1AeLLdR0TBIn
VGUU0CAt0Y0tLyNbpg4t5lnK1Kem/JqJpXEtClkkMw7/FPEvDlbgJ9DxZX7ePxK4
cwuuYQJtgNFCneQENnlRAfip9i7GwGbzEybvkqVY/E3AT7XEdB9nBQayIBhWtOX+
yCIHODKAdQgj1vXkqC2grk2hN7gfq/mEnIdhPhsAgcE6nlcoxYKFXa5VldGyAVXD
dBmzc1uTA931xisKIGn2SJQwtM76RWSOP50jQRCGNazSl08VvqplqvAnwlQKSBUo
u+XddnVxztE9ozBT5rSA511BgHI8JVVEN662AKVYb1HmLBc4xWBvsEDn9FlT73lq
W6pgbx7S2BBAxS6YD0xiZXG4Eo5lV7SMYPUBwqukCXbanz1ZQRGu1DrytMCYzkHH
ss60vFDnzQsWV4CR5u+NNUJdqqXi9+zoHpQXZ/Ih78JpErqxl8x68oKOOkcI/iNz
1/LBJel1DCKbZT4ujMYIxUGTJlLXII1PIHiVuTmCTTRlbDAjbPEi+l7SKhJu1pkw
nDXy9oPnSkE74Dx8vR1IVcyTKav1qK6v7mUp5RVrCByDtaxndYtGO3XzMnqNVcGg
r02hDz5ao0LQD3SJGAqOvqZNN4/XFTs7KGOGwI20hSpmmUZJqaWK1z7pX8mGzBuj
Z/VascUZ2rGm4Y9gw5HtzPMowNDALslpLrEQMUVPftzQ4KNviYvJT4TiW4xpvspf
6lyyiegVdPZ8baSihJ8cmbyFYpP8rz5mVkgxoE8nILt/QEJX2Jg/P/ji3xsEiaKE
1rIjhDJtJeDXZY/qnPtzjNZ0K/c9j6Wk520wuxiM7GKg+5TieyqTug09g4WzMN43
iPFH+CEg5bFQJ34H99BuRSw2WMZgkaJaodOf9A6/c1g44v6BwVQuSDYJLIFQRif2
dYCzyLQBXSfICMslW/7zzSFcDa2zOp8XHpRvrNgFvEQU0tL4Xf1ztH/8CjVWiuG3
9z17A5iC76dO8Vlye4YlvUBAPhsiRzrejQ5OqAEQMwaU+eUqqEPGAeK1Zj1aul+X
xQKGJ8PTjj808Gx9Z6jUtJG+J3Umi3+uiCTot5Q13DPmxd05sCPrsf4Ih1vYGdEm
MJ+sjgddK7m8eN9UxKjq/ylOAZ4T6Cox2n5/JOt12/cn63m5Ivo57YNnDTg9jWDJ
Xf4d/NYyE83MdOIfBIb0GYFIeQlaIan/UXya08aXNgkM6WH+67xQkXLKHWFaI9ep
TKGuZeddMgZexTac8TF0IMNcHyqndI93qsyEwZ7u8gyDhDtve7e2ILYU90QYY2G5
XeV7SCMoDGc5VGhMsoDnl4VC9eEN69Vpn89HjDLpvpdfgQ2NCoDgg7vLwUpnit3n
m9acNTETft1VyyTh0BAtT6Jm8pHeMCMal20gESvp/uK6HbLU5Fsacuk/RafN0ntz
zSa2l17hRk7wNRPxXZtrDXJ9jDOCUT8jgQtiGzTNjXjRFLH1V/qNP7sS/J01H51L
8M3t7CsW7j+g+Kfv3zmbc0KBkwNeVDKwofekA/PpxDIihgHqUP9X7fSwT1D+X2nO
vhLYgh8bBVvS7IIbiWKAp5h48y86nWv0qXdy6Ka0t5I/a8CgQX3Qt3aQ1MRPQOgF
bnuYFTNRuTyiMMXky8fAjDVxiHcEj/XmwNTwvNcpEDho9dWfXqrMFn/CCNsybDHw
IjV/ROogdYd2EQUIa/N+gVnXGgRAGJFbJLhPu38vATJ+av1vjeW9I7q7v1+Qo4FH
X6av3Gv4+bfvFdAvJkenTpa4QHzEImCGI6/uBeEwPVO59p22wAEliHIxDkQ/ncW3
53HVFkRDaeEMdwaWb/coQDjDH8GXAtAzFkxX2mZRXtRKT6b/3FheV7/DaE4FJEBA
WFrVhsaYOpEN0fP9cMflMWRPlS2c360Z5T5eDUwqxuiEfkR6EtBmZg20TyaaPRTQ
UkTpwQIsYVtkalZas7phj/9SdfXNDrAzWSToXy17a6xTyyQrIoYRnu5i0nDjLYJi
5SAYWujbPusYWEZhfmYuRaYuixLWHidN1wW52bcX2iOGZmkVQq3FXj5eilDVYqVj
eMttt0pnLzVWTtsUC64nqsBNQa2RuXNrUFAl1Mzu9a4yP70kdId1OxdiqptTDIaH
+1OrjpKPaR3ewnsImYTMipcZhvCTxq7y9LXxBdIh/gkMDunwNs9L0ltps3sI9GeM
FJlqRXT9i9sioCgykA+Q0YBwunQVQURUfWIilQvpsFfwHLmdUoVQwnWdynBiFv1X
Hp4w7UG+2PwK40pMJMFoLcZpuSOvrqfSKhHZG+mKfn8eQ6IFP+pec85GTH4eG1DZ
SjpbS6aTadmnxMhOFlDD0ErXThPwpHWz2Yj50+aC6ZqDGByZlOWQI49PCzM+oafs
xp2fkgDcXf6JW/fXiAeJmpcd7Z5/1NCprzb8+NPYAxn2w/JoVuOdT0bbJZVQIzeU
IJbIM30cLfEMPOwnz12RUMh7D06u09gXH/E4URo2EJS5mVSzMmPxk9ryX2jpIKNI
U0lzPD+a6FHSPPA7dsl2MMRyaYc/z5T06B8m+IpN3D5ozC700KqOeiK5BhS6Msbx
iI3b6GWVOe1gitrcBJpN6znsKl39wi78n5mLlxurTKUEFdHfxMHRnHoyUfc/6XHN
daSiVeHtNu2eyFa0g+Qz0SXueJD3JhklodtmQBxlX+liO0p2HTtVsa3g22CVtvya
5R6ESR1Zb+/KSxFPNe+9GZSCVKXl+/Mx3yvUj/QZsgmnUzyH91IfnhijpyNR39B4
1BNBdVtSg3WLFw9j1u7NT0/KgauYfc+yic/Li6ximv02PN3pTIszb8wmTi6Mteqk
H6wuOti9qtT7Gpf8flCtZ5b6uXh2ai6o6ZeP1ggLqyGcd76YFtwXMEjZura8TN/R
1ECwArOYK5uDChqp+aucZ3A1bfaNrE95IuCEtS2NhDHAuVDd6xh9J40szpzHByuE
/T3tStdPj3UiUHGu1Nj0NZlXmM/iC+10HC8ePu8Zl7ZEjuVFtH49Ku25JSmH2ltP
tfphi93oIXLcc8uGUu7sVPCy6oWs0ArL7e6y7N9PFyagFqdTjvlTKMXneTY9Zty3
+7FBMD4wKnx4WhZ4b6BaunWMpryk0fE7Rp7Y2N8TlL67Ah8J2vslJnSTloH4E7+G
kUTL5Gq1e+PefZKudTmLKzmKTrEMzwp7XkIZRvpn5wJdoD5Vf5qUGowBhLsPhd7r
l8I3dBfcLNHabUU5RbXXKKL4OUJV9VFH91NPpF80sYLq03tsIfKVxUtjSMEWu0WB
RA576H8kFHagHix2x7LoYYQRxb7Zxol5I/HrpKV89DtfM4kJD94aWcV7BS2XIvdu
EK9uDKFeR7RKWqSzIRgwkCa88vnrY04GzaXs/96wbhFk2pnFGjF4o/hO2poGhbZq
yvxr1yENCbuZG3/OTcJPSwYlNhg0DVRjGdwtydQ9os120G5/bZbNdAWrrHR4eGIy
vRogfRs1AxvbUcDlMy/ww59Ax0KQI8XV4Z7UDjDqrGjbGfwdObL1lB2QNKN9Jx1a
zio/aqVgttVrBfT0x4mEQGTuxWeW8F/yOvUlPzsOidTKlrSiHdDz9ROJ9SOtsm1N
gkzZ61cn3Xzyh7p/InToTcmlHwV7QubD01uJqL190JFUC9DqOJQOACf4ii2xA0sV
/zCuDDak5Al+mih59RUnidlsORidH7iahNvHGd8kFKN8Zdkjqa+qWzXm35093s7L
koeBrEjdp/hBucT9bm8u2L8DvV2uYLByxFL3gkiQil5silZH3yKWny/KfhYNcQhi
+qRA+kWJCM8s+ztBC3h0n9NSXBgvXHC8Db4+xkkIay3thwqK53qPnz11M8pOO5XO
jO5/dmbG8FktD30dTseCGaIsDqmyQZ+rW+ceuhekA7ycBuW+WlR9QZ7AXM/6TiA0
b37JLW5Dr0l91wy1FPKdxprAnRWnKO1Ud+vBmeRkQn20c4c1ZYpFwEj0mv/gdEUr
D7dtA6FHw5c+k/fLg997NiwEG0UyP8SJ1BcwPlLKjTnHtZxJbxei2/RXrzHBi7We
sKTnsQrMsFrIFThYlIrQxPd2KcWHMdTbOxQqeLV43nz/BtfTssdjtRKy09kzbWSF
un1iLf5vUoehMqXB/hiqdsEgRoqNWne2v4HSem7Mowqny84eoZSFzbfxG+RXbDzl
u+1Dd0VqhxUFsZEZk2ERh7GGciRDmcnpvKnYopZtFMFxQZxyAa0uJgOgpkAe8P3b
qaaOjQl27WIcaRECgSX9B4Lg1K96Tn9AD9ClcCHpF1Hptq4dhg01U/EUdGulSWG9
/7ikUzH6NHwg+/u4kSAsfeVDj3eXg8a/kqN7wS+VWbyPFCDBdeb+Ro+WPdPgk1Xg
qHoZIf/myT/xFWseaPvacJ8dUp5DsnnSVxmLOqr/ZicovYKKcwQ5lsEwS+LK7A1O
ViIWNvt0dsrGmbu/os9foLCCnDdeGa9M5bz037ybO9guzdpu9AcIheypZ1s6tjHl
BsT6JCp7xmvZkgB7N2MeFosp0WPJrvLYOnqj39OP1+Cr2ClwILAOCnTpAJ3+37pE
ofQIinb8kwP1Dtr8j3lNtpYEIEWA/cujUcqQTc8johNmLgUbpqy+AwcSAFyMFSE5
IgyetpiLbC+l8GAXPdj27cJj40o3vsXZWXfaDPaBQ18/+ZEhlEIiU/yhdDNoG+Je
kpry1YKy3ojKMq7ByrWlHihbtRpVnrCce9ALz6z5h8aztrhl/y8ykY71KJylnly1
HNkBZ8ysZdkL2S3Cs0AU6FxDK+ScagZqltS97R4fwUHRYzzwYhzIuA6EVd5U5v54
uIe6oKsq6j9fEtOKD/Wa6JRC3AG1gvFZ3Gp6FZ7HBgorhFPsNQUeXDhSozTIcqFU
mumLnZTLSKAN+4a98Bm2wJKtAH8aGvNBw34wTwE4KR6gwmZtsOT0TdmDYyf8/oUw
7yBSol2dNq2nII6LTSeg/o8lIxSijb1g6g8+2nnRIlAo6WC1lnvp0+y9UEaN3fpC
BZ+hRxBLR+qGW2HPQ91FoohGtPhhHUzU8aSuqenNDxv/QRHmMLfM4UEV+jDD84oc
x39c34VtuYecEtl36jjqiK1IBYzFUlBM9R+PQyAYtj9/LRXm/EVK4VRJ5ZADBGAg
3NqjR496lNca9+4T8UhDRQrZymEAFueLJL2jZ+jbiZoKdJWzz7S83t+vbL53JpB0
ns1emCr+9OrkAKpKvJ3GC1tH+kNWd6LSudMdYgZhrMhE5RgQYF5DbheUtGZHFVe4
7yVjmLDQBdSjnOvgqkPqUwEWugEatRsKZg5hWpDr9BhhYJ87KdqYjJ4ngVEyeajt
RFc0tJfwsV4YDAK6HmPGJUAM5sRL4kgaVESQKNN5CKadKrhOhAKjZHy8ZTvpFvkl
mvpdhewqc1BkoFmmnZVzMXK+qtZUpu44pVa+EkW7Dlyrbckndeff7/t7RJs2RRHe
Q8CzpGoAeinXZ0RMfssPSyQT5k16OvvpdRa3mZPaJ6hLrkjUay55qO76kY8u0fm4
ZZ6tOyfus2wOOc9vCWP6r4RT6rPXYmDN8Lzv4GVMgnhjCFIckT/yEOQJegxU+xii
j6ISC+X20+eMBqyDLVPl6Dm765lZvUsZ5BfB6g9/+hCCbEpw8C5yY24jbb3Zt2pQ
/UfCo+tVeXXWfPbBBzdb7qXaubGkBKC72M7bZnuJLK9APm7EBaSP7TSz71xMInNN
s8DWJe4fpEBXHM6bCBwWe9WzCTNcvC0WTkFrblgtKSaKf5rlH9k/GXM0Ycfjwg6J
KLfGu5/zWcvhiyf+u3GHZ7x0cbI3YihQdHCW9EnthPyf3oKz8qGS3Gf0T9/thdJj
qBbaZfPwlIw6NP6M5dPzHQVTA0wSyzjw3/u/IotLw1Pp9+Sj9APKn5530Cr/Fy4r
is8aqdL5UeQ/W4T9PsdRN+DQsw30LlzpkLdj2VoR1mzFAHMs+WtSGcdleBud04su
oYZBEQyICFG1ELNGupXEGQc0EwFRti3gTu9tPjNiyrN79Np2NqHddeN8usiAxpro
AL3n6KIf6tDFFI+ywGYCxwcb0O/7pfwGhufhlmPKheKtInCLz1B822N6SmslJXYz
7p2JO0nGjoLiZNz/U1t7VzZENVsSseO/VhbW/OQevcGD4xbocr//6DoGTxm/0NI4
56WJYsaDzpGwYkVfKZbjBuaKx7oNWz8VZrm6D1s/d3Qb0G19rnZaHlUvtPFvMPKi
m4wWjuH4Kx+znn0/w7kzukRFn3QD40N20QG9eLB3trQs/QxiDk8O37Ssf7Huz+sV
AJntwR0VKx+smlvwWyFysuBY5/bYHG0dH+CYTXftkzgZnpWRZfSZXZJvz6LnO5Ov
2yczVacHVT1LJXWXQ3cO5ca8JZ66fWBdZGLL6wkR4ZM4h/slSrGSEhTuvZGUBySF
s/nU1wrMzPxRZRFNSDocApB4qJKYEfH5Zts8IC/OEMGN/Rm1NNsYVopnA0CFjzCQ
PC3pk/fgnl2LMO7V625xHElE6LWWkTU9XzjLC+jSJUkRKrxEbxqEJ/GYKMzuFV0K
yu/SsDxtGJ5wAdN7G9sD+74zPQ9w4GX5EjDIJafSNRTkXlKVx66Urgs4tq6YhISN
/fNrnrTez/gVdmooyw4r2pmgX3fzirHyxgk3+ss5D6fHG6CbHdOptSlczWFXNMCs
BlgTXXFBUYv5RAfVn/RTNxPGA91Uk6rYH6/sn3wGe7iNtmy1ZxIozRnGxhiMNVrA
w0CxwDPTBSGhaU5udesbLm5/K6/FDoIS+tpYCfulzKG3pjVCMlRXPVtqXksdgh5v
ZDOD46TiXRcZc5Dvc1KmYQLMrQ8qXNMHuGWH7Z2rlqs5CQlxS4Qq7ftFHOPc+Z3Q
0+rUg4aIT+p/v5GOMuaUW5DTgS2K1wkrja1kNSVXkLGO5DWmuU9O/8eq2LUEzjOC
MtvNFRHmTDT50NQsmyURxz0+jHfI/VBZmxTujJrXWcAgJ0aOCUhYNeIB6bpNThZl
D+Ntk20TK2yu98y49gd9qnXcdcasyk19WnqCGqd69jQj/kQvThK4a9kKLoV4JvEk
UKbBxAjazrAaXLv6wiDqLceElLsKLfkqz/Psn4KSG9Yn/t+WGMZuEnkZvngm52Kt
bQiW1j9pKu43prgtbY2TtO/dm9Ig2/dvhydcMprpOR9ay7EhMIO6bI6ywaxXVfLM
69SpP0L6M8XUVRuRouhJzvOlRUSM/VgAnSWJcNSkVQEH3kvNAgdaKq+TnHzkT2Jl
3FeFcTABmfmYlbynU64yKGBmmrd41ERf6Yuhd1mz9PTFown3oKrBk8gLJBISOk43
JrPjanvdDOMERddXjSbrdaxZksFiLogSXEVcPLerfKr6MtTk+x2Obz+L4fdFxHFg
oJpB2+qAT09yy6xEhREI0cgGBsmVaJu88U4wJ5F9p4vJ6JVF8M0pc3wM+KhIDhNr
nbxlR4pyy/UUx9aJvVEaC3Ja5vAWG5DsYIcLx8uiWCndPhmkJ6ZAigLRpiu4hVDE
w7z3szR9TLscYGI3JRmMxVPyivuJskRfnjsnk1HwGtoXyIbuwoKHoNI0TIAuxOp8
eqbJ4zf+PV+8mvFOuSJzrRDkC0OoQLcqN9SF5kpedixvzQRqKKEJioQjKdQDavMX
4OqdVIj4gnkV0/n8sijlU9Ur0VM8f3s1yk4XvId1y8KLvuoxYL2VRLVO6aeWFKnV
XOXt3sUHLPkdNDw4ffsih09hHMRGY3WPwtN4KbOcpe8BCl7iZPMblwFpdzdn3HhG
uw/R8rtPSXlokcR4jtcpn/QDAEBeqQB5slTapdrwxwM3hi/VU26NCGTYxDC0l40u
BBdNk0uO3DI6hJms3y8HQBjyspKJ4D4Bg8QxyssrXqEr/D3DjTE9VRWIk+EcLavF
oGOiDI4pSF3hY4uh8Cz5ZrcePzZ6z1sPNjc7lzf/JzZ7dI8el5cgVZY7x8ahjghi
gfBRDymROAhTTeZ6HWFdy40fF04B8RApcm9TeD2vHhwk4BE1ngYp+rJIVwUr3dv4
Xs5oOn3X7vEC6355rkeYvZa0/oXQA9lkUrJB05OHe4X6HC2XgS3vGwVhBR0t0BBL
b52j8t5lNKXljboVpwX6FFZmBaiHN6J2x+84GEXVhvKsT61tJ55vfO9/e5vOLQ8R
6MUO9g/a9tYHDkndVKUTqtpOVBVJNw6NeYTOQQJoMKC+pK+o4JMiciNYw3hWjW1p
hWMFUs2KICeQRteaeCxsw8Q7zlqEaDABUqMESTrDJRNnYIx3aU7EO/9luLNNjorh
NoU65J6Rhyhy0wI6sksPcQlDlu9I4mFzXZvY0Kf2f9MsXrhEJF1WzVzgu1LUyHbt
/edCKmOHMNx//6wXvtKzmRMzsgf4EDFmXcCyX+135mpBeNL8ShV7D5Bw4nz0LCrL
zYGln7o9EMrZmMTzidDVUy4iR/f4COtUWI0cft5D7LaSTLHaeXw10XsxcKgICscb
REvO5HnHeDF0SavcHJV+Vyd80Xvd9ztcJ71IhK+4Ahc/tctVnhrOBWZb6/QJBA6A
XrD1HB70P8NepuyjBtwjSNGOvYHM7R3CWkAtbhOljKDCidQLxjv6OXdpaAelAPj1
6fgWcBvu2lb0DbybclXs5qhiKVCnAaLXiiM1iFVYdk7+IKlyFmP/o7xyEIp86ADS
vv76gpVZY9TXNePcVEeP/oMLrdTiRONAsBJcP+cjlIQQ7UHAWLD0lXkh0Szl8Edi
4auYoJByHXvO46WJ3sEEdOJ2NmEE76ZWbsbXfe0Xdg9q3YRo5KAjzYynE1OwBV/6
9NDWcUKU/REs8E0+QSb8hXjLtDymYDoTptzq9fqSeJgVnru1juY5GdAZGf5B4N0V
rXFXYwDMHsNovxHkRi8N+Juh1CyPa3yCIKHpjjT3lwX5jP+dYHVsCbJjajC0MkKI
qxUTsKNA5RrCuZ6sbpT2Y3zWX8RC+fJctkn9sC8UYeCRmZ183s4DMSsV/nF8j04A
DlWhBT6U5kQ3ONmTcURzzviaQJ6k47d6vftNnlRAxegx8gEfzazQgBjG7uBFkqf1
HCMjpM9RNwNrz4iWsWpmU4LisSCS+QGdazQYZ2TdkLsiDK4EzouHd59kcci20XGF
uX+No29xUklQsZ5GTIsO8JLsXAItnEM4lxf1LO5QnaTmAiDuc1iujEEkwGwjZeiZ
dQkWq6L69ZbORZ8c63gJOpVu50DW9CdcF5eBAPfTruhaOknpYQxRd8Yug1Im/vVC
vVJ+PYPao3E47HEk6rzi6K0Ryq7DpMZsVzkaq6NujKUS+21hIbjjUvvPhru1xGs1
nMTzC8aS1NNrofYn3HQy2qlaswys6PoZeBXMvPE3pPk/HD0kwqyH3ma3dZwfXxEg
jZUQU1jnHhnaU+RgGepZOYfE/KUekDkLhmy52kpa3z7tSKvyKmyoeEl1Qw1lekLR
LKsQUtrcT1x44e9bzCuMdSp9Kq5ea/BVbj0oNZK7Ysn8pADMJz80/39SJLXLTOrz
jbA8ik3P9YhGPpmGqE5HEF/8phpe7cXr5VASWbhvF3YS0VxzeR6aLyZ3olplJKXT
SYCJSQtxL6kHNBXOCVFMmgRqC5HTBpNi5yUZXyzmZWC3OQAdhXRHMvmjuud+TOmR
7NV/VO/erX3SpxkG96GZlHNV7ppeIDQ5bF5+h0F09eQ8TAs6HSRN+kZRNzRUCHnz
IaK3kZEtiesmE0xVwC5IZ0wNkR3KweeXIVzLsmN5WozpwGTvPCbm5azUsD0mIH8a
JzuMv25FS8V0QJCutQgI8ce+9vwGS5VUL4SWSpIs4hu1erxS/fBc8n8fDQJrQfjQ
aAbOwemPDc685O1GxaRTPZwNNAHsZlQ4eskAjF8IoPJMK3rm2Ry0H+3SOleGkIef
t9oxflMqnK9oZdyiJM6/c7b8kJOUOMY8l5Yv0z0yqsoVRiADayAcj6XsvYlg+tU+
ZQsxrKGTchHoJVIEmvRvGyK5ZF3iwD6UAU3tW4UQqKF/oj2i6fWwOlOEorTEl766
RoWoagpMdQ3fL6NZ+Ghrs9Abx20BMzFRnfu1v5UzYA3167tPM/ZulQ4Gxd/CuxVo
b5XcywYgX2VsIMRTquURiPwBF+7ZRZGpnRElVgMRVVWYycTK0wLD15q4gFKZF+K3
KlRgKOFcsTLWaLHR2sM64JEphpEZleoBmsExefNc/r+XQXh64OErk5RQdvWfmQg+
yX6+u4UpjpmnKOMPTGA61DzhRp1Iu/PmvyySZxZipmkiB+pUpk0aZZ2ZmSjVXsBS
F9td7kutlyVRgh1ha2SHi0wk76bcRa5uT+W4VHYIzIrGKC/K3sVHLJFrOSY/NgX8
DMVYvcwO9AeQpyGbC1ywo5ZtXcWSVstzoaKsOKl7I/jKEmLd6IISAEIqNIQeTeC7
GertTsDrTwcy8C1oYcW857IXBYrmg51G8eFd8vBgbxzZQK0C8odUJUWkQ+bLuDOm
7xZJpYZ47525JAtGfnq7d2HpYh8zr0edjXQwH9E0wNggiao5T9viUZV3a1l7vzaA
0A4xiL7OG0VcjFdwDobliSzwJL5HLNFS5T+R1oNvgy1DwqB1heziUOQuhdsamKz2
4t24iL/UrgtEXFmsr8n+WF7Q6l1T0elvXlFacDEH7+OfCm7a0mWwiacbgv55Tf0D
jb+1yi7416og0rMdTDsMx04MfR5GrOTy/EbvrQv2b+sHFisGIbacLP4tV3CIMw6i
SiuHNtvpl1tSf+ozhwN+O6ijW2tRBjIhxiS78CwPPmtX+Dna7s0E6Qn1uRIvyDFz
jYPOjs6sS/i8SIfjiusEejPIHVt2SVJLvdi76+Sa6HDyu1hKK0mxYEdct9E3xFAP
KOxyH8XzSHE6SCGS75GRdzJD5tdsdHapySbFWZdLSfczaM64S4RncQ7JbCg5St7g
WgS7flwxa6nZAa/DFVCfkbt2KzJkPApFxwU5Zlf+v2FxqVKxLgEGwH9hCvTUENp9
9hakRv0oEauRhRJ35jcGafq0SxTqbMdjRtvc4JUI5yH9yRdKO+PePDh+RiNUYgGI
jOBPqpPoRBA2PNPo/FWzEdCqPDEYCt4Qat+7ZckkmE84dikSrePaLH/xgCxPKP93
pa0nqkoWwXIOulYa0fdxnvc5RAjjMOV48hnEYjtOb7vsFRHizQFQlpEDf/rvGTwE
PWIGXJosE5eWTYYOwY2Ucp+W1sIbNtTtz4Qc6asPsJcxjQpHrSm1aUqbduNYWKmz
dvXSOWxtc8TP2VcTNxBXzMHti9o6MZrwE/dY+GH6xilQFHW/hlViAzriGy+a0U6c
BtSvD6h2UCVSFS3Lx6DT2H5PNQ1BDUiTTf4ZHL/2OS1ObNUY0gaqWlNVku6IG22Y
Who1WssbjPxO5GeDmyMlrWyYYjjXmSmEpDCeuNm2z+tufFUvrrcokDXn1W6sWn03
H2vadf4nmuhDCj57GumdJmRff/8eQcHKs9ILySbQ/Hk1YJf2wWOvbKvrCNgiib8G
cAAY+4+gL0OmJag1VcfImr0WZ6pFQ4Mvs6QF3Xze0wnEkjjglSGPJuI7L/TKBwJ6
gxuA3knIFKsfHbE/jHG+QRUOLdgApyO1kcnbN6/QD5Rk40rS1UR8nR/xMSJp5SZF
boOU8UNxqJ1MOgKK5puELxmy7BZOdA7viqb2uT5CSbQUCzBI1eR920h8LUuEP3GK
59x18Tj27k5v5qxXrKDGyfDDxenrDgMKy15aWJEIkBVx4o+F9gVqIWLp93Nd+El0
p5b95BRMIqD10vRMT1F62X+wTd+jN9kdpsXpodi/2cww+qeYzDuD7PyOI3Vu8aRc
2qtG5/jctNqSQcPHXv8bv9/5DpbirB1AKL6t83RgOCGOpGmqUX2rPVpKRqI4A8NC
cnrjRvnG0PMTarIG3RNW28eVSNOW9cMWIKXf261b3QFfAz3oYeuknpE6vAvUDxna
h3MeY/8jqwqDroDs+Gfz4LTK8nukB3X1ZwiUPRTczLoqY8qWalomxWzJuMrF5udL
uTP+rwk0l1x+JCq+JKKk3uT85Aqp3Ltcxau2dyAVWKWdRC+c9JZQmiVZM7A9rqrX
tmR25EgqX63ty6gGJz5oBdL+TxfY7o4YCWcKUPU3vtzUUab2mR28lFdUCCV7Ym6g
1RInMtPTFCtbOVgd4Sv/poS6oWCPFIRrH5s3vhfzNvITCe5kW8as5yoDqUzQtnLJ
jjEowq/4s6xM6pTQwD3ZD5v30KEi+6ALjUmQ+rylf67w5LyhaqUqDeW/5p0Wrf2E
K99jyzPFzhrB+JIC2/9zXXvG+xGywss89H0P6GUNhO+bfL3FyJUuCsyE4H1whiQn
2Ro277uNBb0EQ/3QC/EZmmlbQCPgpmA4Bj9rnyBaR/xph0f7jkBbqKbzTz7orYRP
Gzi5JfoV97ExazNV3HVki+XMLozGlHyAXc0TRZULNQCoX1wdALCfgejmY+LG28sg
pH8XyjAbJtPbxi5b0BzNJwGdlldhTaouFM6cOsJInEi8QQbvj7BQ477rT/6TttYZ
YhM5pXheFyvPNSBCsc2sLZvJL0gAWBr4nDsft5Y1Fbtsg9+KCWKmmCKLL1w3b7p3
zJLOIi7Mayyou/YeWl6XCCiWmrdG/D0j22wwf2SYb6rGHyycZe5eaTviv6jWbQ8+
FYR9xPgpOckmxt8vHbE+rRY3zUtdrYS1XZwXMXyu2/ayTt/5xk4t80LfgJ1YZf+m
qCPd3o7EsefdFmGl83D8kvv4S63IrX0CJhkj8IoMu/6JsOf8ZHQrpV3h02WogsR0
wbTf5FWx/6MXiGf5X98p0P3Qx7zCI9jyMOMSRPRryi3Wx4w/WvYerRWOFCvwk7vF
hy5cxCvr/ZhNQTyPXptKgXDLRbjcM8fWQlpRKgiNjHJ6LAgxWKeYOdiRLyA4nhvN
VEC7rU/ffT/gFZ/A88fY6rHakHP4pjefJAarRyATeudiSq/J1lYpTU1+Ws0VS0iP
XSynWYU+wk038Zzj8DQgNUSpXtdzgDuCEDyWjA/1erlh8eB0lRn919LsVPMJ7eQU
eX3mYorzA/r3Wz9iMzRva+ouqdgJMSqx0Jc05/iFLtsN9tOrrzjBks+MEbP9dx75
4dOUZUdO7PUxmHUUXjRMqI9Fjl3SFC/LQael0FtVOrUBAANHFqZaXbXLxyntw0mJ
r2dPONproboihKmuAoKOVcNUXTGrZ7sfj1BQHii7+q2OBqQqyg1l9TwvkqmAPEnu
48IBX1B6ClTyoXAh09S1K71H7L3ecjLKJQbVMfs37YYFSDHhPv9TMNnKbcosO4dJ
aA7ZSAYbpNp5s6IjY7md6kYijUUC60lE1BJH0lcRK+SOct39LM2QcDBQ1q68uNF0
s+hwfHNGW50shVFfiYWmKuoGTpqzUQzZs7x3d3inntts90fm/dfckX5+FcaDAfyP
650iafaP6/D7zogiWOLECEEBM/8hVIOHz0pAjpjIjX4a6VV7y+6w6MxbdXWPckNq
NKEdZMeXX7yqTa+4xViOwQ2C7Wf4uqXaCw58gE+M86/sj5JZHDA6zNhxuIugadHz
OuNp2mK5krFlaQrzHDpZA3Pr7jxer9GWW5wWsC9JUILQVS7K6LF8Vp53sAgV0xss
vAD/BMQ+frJjFZvxZp+liuQzkg/DicW4BLYD+Un/njDz3ynrpZLDNs1PeFsnTCDK
Cfd2N3U/Vm6Xj6DjXjdVPExBX3gbMIgLKFnv+Si+4EugnsjnTpr0YGcpmpcC6gWp
3dDbITcYkvlDQsndqh55NpkaKFTwP7PLWnkRh85Iyf3SDAX0I3mXzURW6QkOLX9W
zA10gPHXBpqQeBnXTiFq+8oQdpOo3RpY92+pTiUxlcsXowYS0SJwBm43bU0duOBW
XEpWjfB1wXmXvKuJMY2GR/JuoPKYg4qVK/++vUjsbb8Zlmm1oBZRzDrXX1U5g+mq
Aaf1CfrtKm4SCclagIrYsR8EKqnHUlGL0j9ziRfiOnMw4iUYMTX+NaXHh5/N+jxB
17i+RNkySvU3Pxeoyat5N5zZfLW0ouR0OLIvwAngg6vR35L9ogWA6T6nvjAFG6qQ
o0lkxwSj9HerEt2CNykJQ5jCAmWXn0LptULMZH73Fi64hNaerwSRzp77IlVIFvxV
h+gyB1+LLMDk8fFOMkaSphPuKgZ4OLFDjqmSUn6atWPfh8GrRgt9iysYpmEG+YfN
/oQrz+jtNqQYvQPK6lfrRW+dcZ2qNIpId88d76g25uLkmr1qry90VhqEb3g3B9Si
U8OH1CNFLKIAAezS/+YrMhf+e8gr19uDZff5F2M3GaRdYzLiYpS+Eciqwsv4SkGI
KtzsR/kmcwOiFb+gOhFGWTYBhCc7fcFsNmPP9+vzuVnfm6cjIAcVZPyZrP0ULlIi
htv563aiDAIwusKoJQpVb6IjWD7NCAX4Uw6X1iCikdeJ1ee0K1Mg3L/1dfR4NiEH
vjqVed7cw5DORcR0GPMV6Q31nacqAzh00wN66gpB1I2NIzzznF58GT1PhlDMIa/2
9c7kXT6md1DI8JO08T5fg0diYlsLuUqw5odrGPrthV2oEy8SIvaKvC8zLntKaFVp
ocWw/IYOxXQdtnbCCEcujoIYinbkp7L74oh4OFTNncXGqDXoSDcLU1Pvhr0ZF65/
+Q1Li7o5dpW1snDrzRBQP0+c7YTKm0HRgrAIiqXfhz6ItA8FAHkX0l85bJR/LrUr
Wn3YCNt3QqXfUaB2AO0H0otPIlIG2EN5aQ57PiES4+OLa7PxaaOMY16w+Dck0waT
xEb/W1OiiQEZfV5JZiQtI39CfwjbAWBERIEVzeNx8+M5bKu9YeogXEK6awZwbC9C
2o9wRUfEUPBloYxL+AaQO/wEMeCbVManDBeJyWZcaxrVReaXbJgaKLitqOeTPRX2
O6sHkK3Zs8ahRQUT7KRYU7Zm0cVeI8GuaeKWg++iirzWxj/1W+glUBJQivXNrQEf
IhbSBVDL/Vebhbhyg+vccClKrXxyZ3YQ3Btg4IeWy6T92ylb6SD1PzcD9QxUlvCy
wkP7qauYxd+5JAkY/1V6KumsmQcz2RszbBr8oe7cRrbPo49ofFc2wyxGKYEppYVV
DmMEcxeiCWeU7/NwgH7lPw/OrPF6iJEeCqplZJrNglUjT61gS+txIeTEluPU5yhZ
pOTj0Mu5dvAS7258VLSfGNK2EpxynXPfb8rpwhvdppro4xRh+MpxrDr39ABvyBsn
QMu4UokdF0E8+Aeoqr1MDk+nkB+JKvy8LPLwuthakcn3Fhbjxwaiya8s05Dqbk7K
wYW6YQgrbBbqmP868F6S27hRFS/tSYeqe5Al6kDaMZVJrYgd3mRROWYbqjEZEejR
VCNt7s+ittaBKpKn7ESWepuynan+lfJY/wZNydPJ+5P/y48CioOMi0MuFosddtIG
hJiar78U8LajcsqWxNgHTWIuABtsxHh0p6WGIIwRU3MOhgRAdNYAdFGdd+mxDQTy
3AAQOkBwEVxFOIsjiyRkgqGcV2PIE9+bnqsZjcEYbS8dPztZ6xl5GoYyluXj7Ikd
Hlsdmh7xQYOaaEBo89dmZYSRuWBQrkjiXJo8BC0PxJXMHGfiqJAMpB21ABqLPKr/
6d1YNysoXMFN9B99YFldu+eLFw89lpG4PNIFhcx1VRdgeFwf47F1qrt6QipH0yav
pK0SczmxXGlvKsvUvZ46fykyl3K8P3Iw1rT7bSfWD4PDGDE0Rj6G2KPtNhPKKy+5
RwrWTbuXST+DeCseEvVumVGG9QWcZaXIu2yllPsUGrbTeIc9+W1YRFK62oWbGhdx
jjrZYTPiH64D2AhD/2A5INEd8klQZL2WaUr3bkFxhNyrg0Z0v/FW5Mtt34b8UgVC
YB+7eRdeBrNElpYM4SR1EyW/tl3b/5hK+wkrbT+ii7zHwONlyJMyRFGt3gISRg/4
GpdWXF6NL5MiN4d49RgbjpR0oJetpbLqXfiu9XajsDsroFEDT3Ade5MFNmse2DDN
2MjBtbMwDXIxgC3dmjxYBrNMln9LfPwdtfOq9UkQqgv+Ir/xz3l62tObAWx5tp4a
uHpDby1UrHOAp1oV61ik8hTLUro+fiRqzlqN0OV2L3dSHJnVt6piVZkjNK91Uv8u
+FxoR2kNgGtZLG7LS+KllDXdl0w/hdBZjJGpOb+U2Mm3TktRjwa6jIq390MkStCt
tLbgQI5ovQpfSbWmVHOcssnFSnCRctdTSOTP7n6rfj8aBp8AWHAQAgTKTjLbQDAq
/KTi8zEQVMkMKUhPad0OGNZywDByNVV1f2ZNa5JTXRtt/lS+bzsqyRHolkoX4mnt
HytyKiB70hZfO0xBl6L60i7PkpyzVCBcSJUR2QWDtKw+qF1QlND3sJx7UIWwU+L+
Gn0KczJDlMtkbuCnG8U3T3qzjHrG9TfJtXQZH+PRoKRMhscAT5KPOuTNHbGXMjbT
rzDRWwkkCy50cII/so+sfBLr7tFuZRnPlulCDk0wnNxmaMVDP0f2ZLdy15bdlwM6
ctN3TLRgqYju9rTiGVs2eLHcylMFkpPgA+79E+PLQBmLor330OYdiWXlm7cQPYcq
2CfPNULcEp52/aKV6HuTNrJLU8Mfw66ssuzhfOC//0GjA4zhfmziBywDkqe9YLZM
2MuHrMEQHyrbOrILSmiszHrHK6a0zMGGrKwofK+GmonIhp2NahV1q45AcchGl46m
ef1sVQSqJhrfGIMHR3hzO6fUGo3+Xog+lIWnoonNzvHJ4a0pkYCRKDXcFcQfPK0d
5vA2LKwIEOAQp5/P+wTqUno924fKrwvEOSSzCFHQpmoUz4Wi8f3MJJbrElIG6cT/
e3loar2roZgreNq6oaAP20GvOEgvzM6rd/N7y2uGHYwhrZ9YuG6YLfQ4kUmcNOtO
RkJhGOTEbw6uij8TCY85BWW/5rfP/60DYmT/PoTQZVfY5OhwwrqlGpe7FcSGPZX6
Mcl/fw7+EdMwQiLj7wrQCIQSITiT2rVUBl2O3Nur35TEns8G4KPWU2hqjvTN1aDl
BRPVe5yPdG1F8xXC3JxQST6+9odKr7khQfkEYumAaQnTGT0awDU7pKAFbfPUY8+9
lbqqkO9HI5mu1gl0gQouFc/GcGjCYd6cn02Qr1iGQmgjdq4RK14S2hDR8VMA5QU+
8NnKsCxuRz+jD/itPBm1cU83dXfEHCoZ/5J/sci5S0q3XwDJvu9kUO8w2cP85jjf
+OEARqfxEc/FTmIoBEAOzPFlEnVjXhIDPUWkhEIIJc94eGpjsBiA9wEvNJAWJAcl
HXpCJe6IgYQ516VL1JX0fph8WPpUGDiZq+FR176OKlTOwrFtuN7ovzYBhSuppCBO
FtsWnt6v9NCDBgJjb9pi1gh6c9NDTjFUTp9lOE0HlUVO9YLCDSy4QXvU/pWFw53q
odd6V8qiy+zGb6rxoEXQNLnIOxTcI/pydCDoOBOUix8qqM1iCLR3zjJ7xA3ObLd6
oEcLWWJqLSFHC3djwoUvLAJupV+i8OvApp3waOKcLd67L3DORpdGlqvdSBlJpWEx
hppmGw7UDMgMbpLLQvdKxIIsoLyJZN0VeVWPKeFPbN6jGpFMJnqrMGn+gvOo8QTR
Sg1KFLg1UlCv2SB2+qRc9GTHWz+qzGHA5wzMw0rH5TbyQr8Z6HMgoPmFYhaiaB7M
78mzLQovX5ebr1mBtQQgySzu66VHLjcOf7BvkFFru80B/BQGBKrYdpb9+zNHT0Zi
WlRo2GvSEWk4sYf5yaHfmafz79NHivO0Ho4xxgqa6dLR88Tf+i2YA0vLHIu/PiyV
0+npWCuU6/qy+iyOao+DsZXYHF/N12cM6WXl3M0Skm063TRGp2Z9CmScw70IDCW/
2A4uI3Cf3eRYIrIPq84eQ3HGWoJEIkjGHL+nN0xtnwXRK6SkbpRWA7fs78Y3t5C3
StOIWlNpKEre2WrPH4abSbXXs2Qo2eu0+SmwLhxTj7ToK1pfosD7FB3f4lyYmejN
7iT5RY9m4stjRa4ofWFaEfkwA5rUJ1Ql6J+iwX+muPVlUIhlGKt0u1pK06weR0tl
yVmMGmLg7zR1p2Aw9lOU4tIG53DlZfTJfmmcePYySrM7zv7QMdSziCHA3SS+lTok
Pdc13qrdysX4uwe0VVi76zA1Ns8LCtcrNKJ4yPws0b/b/CD5R1OJiuOBExT1t8b9
wMf04+sqhM8LybNGau5Fs+8a7nXESWd8QnFFMq3ATDWL5m9XYdIp5TKn7AH21GDi
lRyHyoYwVt2OP6W+hZArhYWNvorxOcz48fCZtmZdnf56OwXWXTJaNgfvFWXQJdAY
cyHJSfSO/ZrF0L9d5z8VlcfYMEemVFj/RUnAwFmKv+bwZZbaVNp/ZNjb20Jjac+g
8I1110Rac04R7U1S5yYWRAKxoPI2+d25a5ezFWSndBSbJQUR69wAuMosx9z19qzH
6RMPVzuIPwSD4+5W3BbBmbkgzCZzJD91jt8D7IdBNptJIQeXfsnz7C1W/XDfoIxm
+FI+xR2d4+gOi6P+EE7ImMm8dipe8wXg5KZZHq5VIWiOHPLf/3iwAre00sE+ryOL
sOxPYSzM/yiVM2skmLBnjwsoWlpUkA47ZTJwOFSbkx7Guhzzhd76N931TKjRPHDr
UOcR5LdZzl3qxz3mOKE5X9hmhd94hp2RQfLjA2r6gHBSjQZGgwZleW7YDnwokBzT
choMnQBwo4TSffcdiOJyGvLD4pkGIshISy4fjHgyqcLtE8ho+4bJJMW0ajuRCn+B
QwjPrd9ROlu3EWxTvYB7t+BvOuigJW8B2DBTOQvRS0uaf4aMjJFi1gQZtXgcf8tz
zrz8DWRXMK11iSiCasVlmqfCppqUZxFGS0Of+OUwYP/1l/tayuHEY63lvLL+gUGN
lhX4SMWFp7BX8KTY5k+cEyOqcZ3nlc5LypP5/AoQR6Ul7432YPGNZvCgY9kT/zxT
RwUUIZ0nndoH5MvsiY6KB2l89bBwFRfymFSPHl8yA4oj3GIGRGmSirgMzXzmwlTG
tzLaX9JP5YWmmp8D/q88RXzSgNHPUyFR5WRYzr/WOgdQnO8GKNcxQgJj+70xAC45
jKzvMbu4BiI1JqyIlgWJgMJkxs2yUucG8XZdOMROQSAroyWd/ekgp7/4euMmBo2B
ASGYsVuzQsNrdZ7yOgbzXQuALsdUGpyUVqUCu07q6XaAy2Pq8ILSr2/yj6JvewmC
Rp+UH5uLBWl/4mN1jQQFtr+YxQPM+NSB+06pbprn6ZA9/mJfl4ye/Y6QSuY5uTJm
WpFReG4HBKG+ZliyZ7Yx7UIuir2D+4i75dW0nIEGUDjlxtFfYdDDDshKAv9p3+cr
eT3EZ/KhOS6oGTrJihxky3lMq+oRCRk8qxC1jp4XfgzVpINumMIXFFDRuLrITnC+
i5Av8j2p4IPX26/ZipEC2eqboT+G7dk874wycewqORMSnSzNUTmkTQbJSmnIAjak
6VnLzwPTkjnPjHDXM7YdjiHSH4OLTOIK/vxiOce5ZrllDPWwqVDTu++fGqSFIQ6B
F0UbffYvPkVeI5mhEUH1tntUlPzOuo8XUWhpgpeGs5nmo02bZnW0l5ADw1yauZ3j
Uapu4MByKdPc8x+DW4O3/4yrxwoBuLKS6iWZZ23JYm0gPB+TJ4dH78fwbeogaSt6
u7jPkhn+k0EqwPG5IXjhuFJS0Fu7ZvCheS3fnAm2q3hXL/ZkUiFZG4hbK5ClIs/i
a4Tz/6FWSsPPl2JHXUIYfQibCYIqxLTp5Z8rWm+m1TdvQW/Tz2+I4zY8fXoCNKEG
e7L05XuJcdIaUY0g8IibNUVimPjSfWFTTPOH8wUNtWigrP8qZ9FOKQnhrZp1fNgj
0TUgSI2zYz+9hBLKyvIkNWjaO9Y7xSgZoke5hfUGu+XaP5lsaGG+uU9EpQD6g4+I
gIzi+6PvDN64nGEmp25lNqYdFtHfu9QHOnjDk3rNMIndIYmhv8vy+QI5jxdVflGm
7uySBRRp68VaE3bQNM/tuJeKtMYoip3+q8WVGgKj7TUtJyELbwNTve/bChD3/732
hM8CS6Fj5BVgjnYEQhULaXY6zblxgLXMM5QHuVRi4XPIQSHFgwDn4On7oLtckRnG
Al7JDUw8aw724IwhlDqd0LGUTnfvOuxTyebDl2nOjjcT9UUdQD67Qli15tHDFRDd
vfR7a4/8LwfSASmTCz8Rc4VtgmYo6uvCjrMoS7k5rYHlW09eTwZbW5wtzfCFD0OG
vDoeUidHax0rEApvcSyifdTzj78qtCrmdzPIp2GprPKiku0I2mqpCeRKRSN+oSt4
8P0DbJsM4mrQp28ZhwSsACIK3R51WNOMjpX9ffgZRuEi9KcxVdwcECartCG4aKu7
woDKHK7YhExPABD9dqTCWkkkQfSxGEkEMJUln2PlYPCzh14D3jloNqLQ8xVfiqPO
vp+L3Mf8z2Mv1mM1rUKeFeAPiyaLk6Jyqrs74CU2fW6DIXtPS1WA0Go4u+cC3TSj
Cq5uS2an2fRwMNhdSNa3/bkTPP/lQ0aajIE7UN1+uKKgVdr71zW5JxHO/vxcXzt3
RO/WfF4Uy/HpPWChwNy7AxHAXddbZPtou+GrkE5Bbt0ZXut04sIZxSXZW9vpzJhD
QRm8k4VcD6S5xzvi0cHVuL9mDvpCAza8J9JTsWoX4hupjRpsXFaP6BhxcwkgwYDl
XCAn7qoif0Et9KMWFh7rSdJ1GjTICfLJsV6gXQkjbqJfQ19Vu7KlRZu6MCzGBOZ+
IeF/a/qq0tF2MRbjuMWuth0beyhf1scIFPZvYr5/jAp1Wj4u1bTzm7F1L6FRNzAa
eh1LuW6PjElj6j7wKascMAak0IFlKCCLi7nDw+K/YV1J5Wj2Uk7eAIHmqHlu3wUf
b8jjXVbnZzuobnTAThMxEqiMper0aXz7KD+Q4gD1N44yMWzOzyT8uD2ztS82JXz7
+jFGykx/Yk3uLAHmiG91LPYpa5858ltX+uBgu4VmbKJ8UZxMY45UnhRVcy/3Rx/D
vUaLYMdxzq0e/u7iWR25vYjZNz4oMLXKslX5xeKaRV7/OAAbgg9pWOvkBTxOTxT8
814q8oPd5k/ooApVXaRuJkW+o6wwiTg3Gqw3nX1Z4Dj7smplHqSK23yHY5e38t26
Ov+Rl6hKNDsthZHRbFxjdF4nJizeq4IZR66cDkqrvjpnTWPRWt5wnhjzYXIgrsqq
gzzJqfIkNJUWc+ZbNteZhlWKRX8R/K7w5Gq7VL88Pnj3Zx0Uf3a8ygA3QXa7xVTO
UHJNP0Pi5r/G5cTDSfawMCmLyd2gyMNM6al4Ct0HDCJmbI2j53W08UU6iDEeVcbr
57goY8krq1qHMm54FnaUYf6NkefJGiCs9UOpLUGdBFdBRxnQkf9imsXwbuJudVTI
P4rTMBnWCqx3pQuV8jysegyfnJpeb/Wvt3J+G4klZG2IkGxENdo6tWlk1jgB/LJx
qjeHwoHqs2P/QV+gwJEcsnA2GJuefh0XEFcs6s8qMpzZ//h2TCWAEJuXz6nymtZt
6mGq7qs9Lqd1UvGHX7ApIhamY2KgiPdYEbKWjMZ1fNlw1vAU/GuxebpXoDl+TPuf
MXGQhGH63qyjenr4z84qgD88+lTBgpAz4jRpHFGkDlX63Mxa4MK9p+sKlZ0Lc8n4
Ldo9DgTrQhe70OpVlEMNGgjRC6RHRe3obDFRv0U4F+m6C/wZZljMcp0Yo4LIcjub
AqJB/v0D3/Eg15UnFqQ3DKZS+MR3poA18QrpMEPBCZw595PAgYr8omp0zoXCvCDZ
RAnrS/ni8Ifm4vrbb+gjXdZLAoNHdOM5+70hmVfG3ucCSM/0IO5TiCNCAdaEk4p+
32m7VL7rW7zYBM9TN3/dBMt+QoU3f0BtYNjfQE5l4+0VFySIiVc6CjXS20sRA5QI
tvEqC82vZsdBk6y1m0n6UL7vsZW80w7368q1bpqsyfpF+BLy3P6FlL1zf3UgwrNe
UeC8aE2ZlaMYGIjTdjRim9eJ1VqyrfnIw7LQQsJ1KX8yykh6TL86jkky3MRBDqI5
cLkhiI1rwI3rCzFcyxDCAOIHEx2xvjCS8tVTUyPn18zU8GBWnHbzkEuhnFpxl2zh
5a3W9magZcxT5dfss+RX9XPvrBlVk7bASLIFwq6bwuGWgcAsHYPXSt45FS+LFXwj
9oqUf1wpYwYQOWlXCoh9lLOxgMVGAddWnXl5wtD+x72H5f8RaGbQex2T41Z8rzug
5bNDRH2vb7l4R4aLsFIxG+y7TbHIKKXwEq0oqLppGtFf/rNqFkSRbCRuHfKCMWLO
HXCqaS5/DkV6fPE6WIwkI1vif5CPMlZucafPuK7zs33FMEbk7RH8OfNWgr3GSUVH
spXP80XuuqTxQ8H0en+qDBY8GkQrW4Gn99XjmqD2iRRs3tpfF9mfM2rZHLNbegfs
JmohO56h2W2t9SuwkTI56OhUAjFjNU7nQ2LPdJudtkxo2igrK56VyVs9O6kCJ+id
Jk4CkkOBM95VXPvjqy9FLV05urNDpXPwPWoYoeHFrR/KpvnrKiqaIULYlP89PO+j
gE+5fgax7Qmcz/XA3GUfZiRcjOGxvwH2sB0St072sxCCrVMCD0UtqHaAx/kyr2lN
IOHX4rIOgZ4OwXEoo2EfDAaNpym5REZYa+bW3u2YYl6Fvj9lavTNHtHYRYMJvQh7
8Sek4Lfc8ySycgQ1JE0ecz9cASB8rDMiQHTTUgDBOCuZgw1Uru+jcjQKNNtfCGA+
CB1XPc8vc/XXOMCadrBaW/zTC4sXYaAa5L5JUudX+Q4HiOtOn7P7/W/T5lYsYmac
P8ySyM5F/1mg2V2kY4OwBOWCm3ohBd3FtCNiVwsYjHlOta3MUEljoR68hr9l1eY1
peo1jPzXtUPxe/aftt7p5c+G0F44bztixp8yqRbe9ZgUqWbQ15fFdfTIvZaAJ29A
2uVZpiRGctg86nPqjUKiBe1hH60E/BPXzqQNMsI+g5mBpkcHbpZfudTSeEmTlawK
wwl/TeM03okFENrZ/LBCNwvYIsy0ALh5VpGum/4YdCn29Hfb2Qar09xGKYQDUWGO
2zUczswp3QRqFxiMrLwGJPSiZESetoOTbG4ZaiobSSzX/tcEEmF2/q4Mfb9qfHMW
kaQO+XK5vT1IR+9ObMyqfjLJ8z3AuBgLU7Hl7eHwK7MjCSvvYYOe+iOSS4Q+13Ue
OsIiJyXwnmmJn+oT14A+aG09wU7gJQ7XZuWue9TX3c3AFBNNNJIXlRmuPWU6F4cf
slW8u/xLKkTazKRHZRxqf37F67do21GpRpGnWa3kKdmLc1CsrScNraczBXkj02wI
3f1DUEg94P6NWG8r4+nailRe0vsfcHG+Y/6SOR5nJfG+CgFqbHcGXhxryVzrFAUy
nf7cQlvZHw7m9SN5R/86e/jwfHG+LPiNkSSB0n5qYGsJmzdvFSJ35ub2sX7l7ZRi
7wJSdpdyIte1gtHImzcJKHf9qsJ9Wt9qMw9CwvplUIfqxgTgIK7W8UeKpApDlbzW
sHsCPBznxwEuuH17hdyCbDN/4rZ+D8LIDkfxqco35+mzLNmCfuUhR5r4pKecq0qP
B8wDYq5nXv4ohBGXGxjktJlarK5TiiKl3Glxwp3mCQ55LQK7JvpfAEPHSIjPowGz
/7lJPXScyzztEWoikMOWtjlOmiJSXiVKJeHZxRhXcjn9P5imfEphkytWghB76+ss
XdjYUQqbpKH4zAnM+FKCjiXl5GM026vl3BgkYjDtM3+AZsobB3POVVay0HwZ/kzx
wr1NeQn6t44R95ThD/ZZ70JbybY57WBVhwkZOUeNTXOJw2wcpi5tmJbaQFryr1fa
LZgIFNeUMi5wge0WIxAlV7H4c8WDqwcJ22v5JYkgf/JazVF0hMMxDzroFR4cEwmP
aXsyBmeh3REUG3T6UDtbsjUyHAVNgQco3fk5x02LBoYg1AezSeP6iY++a/zqIRBO
fKTP+DYuoZo31QISdQ+413NYINbJopTMhIxOjtgkb6xaJGTWLy+JUalPuN72cP4v
PL6kT5D1GspqD+nlOsFnLZ93z+4VakpoKin+W4aBfUSrNy/Yci+wXhsoALL1Aqqb
uUmx80rS3h17V68TDPcoAANqHnOYLAsh2k4X3v1DxdCat00cH9PVXechRCXJNG7L
XaAGRSEFVZxjxDAFvyMTKWSIs2Zj+5O5U3RglFiE6SUof31fbpVmXSbP4eaCM0Af
W6ifP7/lmO9pfeEN9Lu/KCv6D5pPYR9S87nAGO6aEyyGL07TuO7yv1ikefIQOHFD
CK7pqGVDba/mfksahGCpApFjbWrl/70vYOnVtJDi0bzkxJxGr7M+nhyYRIE/qc8k
endgq32YrNXvrqAsjCGoKB4zj9KZe35fR+ROBw3PySXyU/m06dElzzUuAgKHdvGY
XZeyln9yAiWctJFfRM2TcPmlQL1iL8RZwiC6z9cSE2cFyyqN0bN7g9M4s19f311a
6AbN9duBRy2g0PGCxIm7GLmCeLmNuvIGupIwmPxXT9Xzp2UOEaempEa5ZngCxW0R
Ch5qneu2AiN+1hsPsCvg6MyPcVa0Jsj+JRANetTn1U0JVZHzE+pMCRCU0by2ae2K
w05ganE1yD8gtWzxiNqWX6BAX2isIOiurY+omhT61OYMM3yvJNreHkWv/sK2pc1j
PhvPsIkaNuL+ina5E0kskWDJ5QgCdzRjaYY2/89KbjGJugQ9yy89fcPF1jzjuW5n
zGHj1bmKZPW/Iue4xDqnCJDodY6xe1p5YQd4dB1NyDSQdC1Txwi0ScfVCkzRFh6k
rZGxfOwOQr8U6DsD/GrjDk9o03jyCebZxmO9kerVEiCMhPAtz1N2ilM762ZUWugs
CrURztw/vJPYfLeZmO4ousgrfoH3SEKOdNjeWxbMGlAczeZTUVg8KnhqACaiZ725
UNkgTMnKqDpS0M0FanE7LgSwBVmhvwKChgLR7tsH2wqxbX1Mih/ML/KLcJxCGbOX
T1TD0FcP6BHeScs34wi6duFv9nkOzb34nX8H1KM5Vy6eypBKNgO7+1kYfa60kJB+
VBl4y76X4gJgiEN+ML5xonjur8h2+UTKP5ka+Ed7ZLrYDLO6ZDUI84XZUxftCHne
5lCTZqZUTc7U6BlF8NLS6pKHOd2X5r7F53wKZvSeX0PNmg91jn1R/XA+fCWCJrQ2
gdWUhwezHV5U5dQBg5O+aT186DsVu7D/bMA3FHWXMf1YxyKuuCCQ+N7n202JZc96
3ZmLsgQC92oYoWwX2bdr2RSptRa7NaWe4f0Yfz/o0sPh9bVS0GtOuJje6WSySLmg
jqoFJr40wye9OPAVPBYBmTG9b3WdqnJbpyj5Qpwn07Opb3NeI8x1Ceb/vAl4DmNJ
keFsL4j/FwdEmwgBjzSimpq7B6xFojxvnLhuzeXIjCsDbVP9Se2S65x5hEEXID7u
S8H7lzZhHMbunm0wBvVWPih4j1RPT1iOoA064+dlMzTrYHDPe5O8buh5w+4yNyqd
PENwFnV5RzJpTrRPtoZV1oo0Gpenlieh4Sk6NN4XjcvrrRbCDJrbQxCiTMjhDSRd
CO9kXmncCwWRw3QuH4vyWiujRNxuxhhsc1y74yfDmhfmFmvezo8xi+PqRPNSyL2Z
4zcbpfXg/TOmU1ByLPjooDEfdijoPvpwbGlZGB3Ql+Yj8WghN4Sr0PSFj7h829Pl
EWEPBkF9TJVw8yZcPKXDLv36H/6A1alTKQj0PQg+UTxJcW0g2GCMakuFB0ykqFU1
uFnSFCFA5/qGEigjkPIFbzgm8xwTNpBCzFggJLL8niYvh6nn8Xt5vOOBZYUgDIIH
pGFuSC/p6LiXZ4t0UBBEdBEKnYYJypPDFKrxCGQflkNnS+SuZDFWxpwI0zQ8OIES
6P5kjacHqomxK84oLldHc/V9fmynk4nG1wEdALlasLHs1D/NZVIpzxioFaj6PQen
3PSfCrApvgiPA7TxR/J7C+/uNHPFcF0j3s0FYQMuPRnJpWaWgkZk4QmpXsf9N+N3
vFB/6I+nQt3R1DDzCwi1M6txaSz9YqmXjpaGRO7x5kGflXuBrWgzXKq1W3w5VUqO
q2aI5uxCTA3j/cfHVbxtwpZ9n2SYOmfVMH28EH9lH2auCUADMuJrkGL4qLuq9lWh
Yi/JPREoomToLo3azqeNH+TQW4cNLMvpy69jXhW4fgUqTDQb1bGVMavkPbfeTnZw
34pAZxKwnKCdXMa5RRXx130bPKjVoTBthppoHL2UTk3JrReO2FcQGhtinIWSM/yC
JOKr60sGKJioP0YAwkxJOWhXp0puJM3/U4c+7K9thq6ZZiQIkhMjOCQBugdXFpb/
shLZoCJArDr9XcgmrDrdclLr6YQHCeZ7qxLyo1kwdELSRt/fP99I4C2GKYFNLz1m
QU/jKBl6m4B7DRSgJJF8F5mXk2zysQatZBpRuAVsmIH8FEvwyRMCFpcBiZw7XSLs
REEL859d7ksi/LkdLBSlbX+DlH4BkKYbXEFeqI6te7GX9NSkHN5EpSOU9GyzpXho
WEQooiY9sT09Au4XhfH98mmTXZILa1fpQ6Pvk1LmgsgGjbclX3N7wc5b2kU2XAh0
4ofhOMvvI5S17wFWvsXR7y3Q0OSiY7Uj6BIwpoPEAs2Alw8/CY7zIcHqbqPSo9ew
wGgjKhZS5IN8CbFz6wsz/LKw9nGMKmGCcpXLnPMmvVxb9htcOVHTTK9HB4xJuWIL
7tbdi/FRKA/r35mLZz4l07Dz3rZwN7QBzSdCqJgx5trhEzJ07vieaAYRtT5z5up4
g9hpYDFLwymW3MKcsBZkNcrQ7mY+gKawBDWGO/ly1ks6/BMy1aNHVDTNoCipcoRt
m6myUzPnv+kbIOVDNRmxLxEExGszcufLxf/ME41jkfuVDVtId0UJe8ohPYDjU1g3
BFse/BbiN6ieg9E2rAlO7ivwFCGYvKaJ+9v3Gq8KoOAydkSJq8PbdSgp3iDagC3w
7JJ2lIvXDC5lCFZ4z9naZ7aR1ZBRAVCFauOQBPrfLVWtiLdMorczZa7BK5CO/hVk
XHZa1HkDpchCJyZqSHdhML2UE8qZJc/Rw/x3+G05xJoxF6teeytvZ7LJdwV2QdWw
RqBfUQUEXii10WnU+mLbl6mkLiQ06293rwx8Kojz/tPu4HN7jlAhd406Z26MvC/r
oZI4hj6M1MbMSR0FApWJayLf7P0JS5kHwmP780AHbVZnQOKzmckBiwpmLmH3TCVG
p+iieNynfmGH/9zmbeMVLpyL3AIga/hC1hxLSvXtRCfatjLx07JLkTovuU0PWALT
k7OwN80AQHl0SR8YyMhKHwUQOOqIlbGSS8c1JwtmNUme9ELA19sS+cZBNDRC2JPa
T8Nkr9emaWZgiAHcLzK2DwDkRaCPV0M7hJy1dtZ3HmxlJ3QO5PPj+6kmv9RvzluD
Gd3f4UBLzhPpYWsbTDb4vrAfrNtLsgJT3EF7D/jXbGLUqil2GBB2vsKrJOjl1RPY
bejJwONF6sAooMb13RXw32bFWiSnkQi85fgvx0c49/Nc96adfiRATfh+XTJXWegY
mPrjD7gtzclO/XQA/m7a5brFfwIoq0ROLIXoLvOS5QIsGFhlWrnKeuHdT1fVkBX0
zBxwUZSvK7ip4EHhI2kwU4KWeWWvlPKYJzv4t7GvF+zFLXq2a0dRUL6ymPYhD60R
t3dXptFMjcYpVs71bDoi1UijihICbOLsKc6ZkO1QUEXQk8G+flpJofEaa1E85MXq
xHMNiakeV09t6rcg/1M7jlVb/avkHdZvZ8mCxccPKUlRP1JvugCAREfJag1k4iHS
2mUo7pJRo7OUsS075k/4UvS0JqD7ZYA7J/06pot2HZlvCTy/L/slROBFyfhnt0UN
mskrHnwLEHptz3bEb+NybUaPloOYXlmToBKSJwEh4unLGeunQiREXjgztLE2NCag
HmItqynd/PRYYOrFkJYyGKbd2Uhp8bzxfYfBu14GMkDB1/qTr3TyjbrSjnCgW3d3
rPsp1jW1inJ9wv7To35Kcr3nqyK/chYR2uupqSP5WKBIxozp1/sfeJygH5VUHltv
GZ9ViTVfQzK2bv5dSywyB9kK2zjmVgOAO7IjHjZuWMc9hGd+4k3d1itpdivLP8s7
/wG3V++Hh1Mmel9FRlwUAN+onKQ8I7Hxy05C6vt/l+92UlteQ8GZNvuCOZONLz70
tHFJVsYVF3r6Z4azvRUpGLR7mjkFQJ9VWfuSv3lDRhEMFejEWh6sokG6h05Kjaba
uuKSEvEzd5Wi5r1IH4LmOoPoxucgUFLHYoHuq6DyxRL251l9tCopIjIz5g3srhHI
2337QLcG5fSSXWE3v/dBa7HXeFbFa9ZJR8yS78Cr4mi+S0gkCw1KGz0ak1fK/Owl
HC9iBOEEbz8yKsIZzjyktm6snFNddUdVdv1BsSAeB4HQIznTum2ECQf8BGoWkyhX
rXYD6l1HL1Er5MUtlIUJBXIQPgmpGLfZe9ksAdo9B4EtKapR/U1tuuMxNP2uVnrs
6i1n+rcU5tWpDKjDkD+RS6/vLhMyS5YicfLv15EwYNcFFyHsNf6Tl7rc+5qbCtzJ
s2iH/fbK5KgURgiy6VO4K4oO43/sEhrfUDKvYfOZkgocLIZuiOCPSivb4TyUoxoR
3NXGAN5A9gE/Db6U2A6BrUXOrRQn9SUtM0ihUlGBZyLP7Dpdi5WmO+BiLVhyn5Xf
Rt6aDLH1pZSqFmvskR6wHR4xmiZNuRucAHzIv4pgjFO1zd4dNExlhda3jxEebpzN
PDnCGE4j2Ct99hzxsYLrZFe34yhcCsGlMxHcCJsny9v5RIjQej25rb+xIysIgkm9
x8KvZ0ASI425nrp+nYFRmfos26cDE6iSYn2hny2pfnickn/0iVOTWthds70Ni4ps
0Qi0cX8dBwz4qTcjB8yCh9svm+b3pW6TlAXmoiQZkrfNDtwunOnMNbN4Qx4pGYzw
XpPBQAEbXBFwSJ1dXV6BzzoD8woYtuxSomt9j+FGL2kXRT8hFNKuLK2SCTMJGcVk
n98diKjFFaZid8zD9Nm+dH5y9rFPTgXKdpkhNAHhcbGgAWnqvu2GxVFPD8Or2oCW
mnddwqzRGhZLFc5gjPbONcqR6HREsASeiUJpQ1PE/52VNWk20g7v85Rsrn7l41aB
J1qHSZaBft2zn/CdA7YzLlvjTuRrMmXOqIXTJXlsv90GWPrUP2WmX8ZZxedx9L58
SxUrnd7znYkagjpJ3UY19ALnVLTpugtKBbfFx+07kBaAmF8umVbFYh2rshXifA7Q
tVrj25OkKAnWAVg1LN6yDX3KQ1azx+4JTUHu+EYzDqf5vJtcNZG1ATD9GhQkqktn
E7KaVhpK5zQukUfX7pKSH7s7SW+wYJJKzkOQkZbb8PX3GkTrvZxwjXGdRYINFB35
5q7H872W2RrNXv+Ulsf+5Hc93Kndt7S4FWGYHvaCZwTuoIKMLSNlJXY/8dRxyAlm
lNijTSLG4wjV9UiBjnwui3UvrCwHToTmYTnfFHsLAOTdpUlqpVRR4NagsZ+7ddDT
l+E+CvZZXAxqkqd+AYaDXfD3sas/ObgZhb/0BEDP/Zdf+Z8sohY+iQhPtiSzWAke
dpGp2Qb59vF3I/9MF3BPkVYLyQKHDaYeGaUwFMXGW1WjfInKIOeAUK/wcg8kT5hF
TglJzv+Dn+0lorwJHD6LJY/ZEnl9sJSfrwYPmiQao+pjbJjvCbOGJnII+VLxhGmR
AaNFTjKksv1i0Co2Dqc7ydGKTDz/SxNi37YAepFn2WUWi1Fah6DY6/IzWngVJHlE
tDD/JYkFXGBAjXHvloXQaRl4sAjOWWPd76OfNUyB2JjwULGtwH5YCyXmCORDy5VI
PubhUnY4RQV4vF6OHWuOSasblt8RMHZhSF93YDqCFUjoXeLjA6HKDbNjQIWia6se
I6os9F/FrwRgECtZ5Ph4HnP4gm4andKboftkjTcqDkhMqKvRrFIX6X6ngEFo9lEM
rgEY9WwFbZ31i2DjWa5Z+QEmi7JM9wpjc7J19ZCjJK8DHIYzJ9YVeoe0XXpibCCl
uCg8ByA7m9cw7/6gnkwCH5hBg4QYYvsxeHIky2U95yU2gEKiDsyOAp8V4meCwvHG
CQ+XIeecJENkXp0gkZ3+jyFb7fw6IeeZgOpeQ7gSiXqb+DU1/+ueqm72JpilHqS1
HLMIQslKB1JXtmryJju928buyHD0z8Dsl5fvRCqKdgS+2d8oqajZaF/4UF1NolA8
PLg1yQC+pCduTxaPDeud+Dpr3Sb2VmVo9Y46d9Jq6jg6S0osYvVE0jY8B46EevrM
3DI7s77PrfRIjxO91TBYQyMFWlzIogWJwwY6wjBy/u9KW3brxevH9EYffT3Ya7tG
cCKkvmIXQRGQn5caucPAPPUyMxZCAAyTMEHJz8n1ll4AE875aKgpPDbAiioaD2i6
yMl5FIy493HCfGub5bX0NVgRjGIIKQIe0/9+v9Ow1EesY94sWrRqtmp78JfZLQm2
QOIz1PoX7WwfOE+TduZleM9G8jVAKdvADiIG0nz1rbWuaf6haEhOHbkwkDyu4FJd
I3X1rVABxyRv85iWW1phFESyIKboaqKzvZBq0Uud+Kso+L3hRMXFeLbOw1IT0R0w
Ea7l2KzuBUolXdsWBHxdujNSe3Li1uCoOkMQS07WE4aSuSICWUVi+HFS2mkyl0p1
2L/MlsSSTQKPvU7WGJobt3vqp8wLymjUQEWqgJk6pD9ad7w+11l5yp+gs4KoXQSW
6xMlYDQh48N51FHoenT+FusWaVXsc/7QuuSzz7oduI4N+ix3WK8YjmvjrXX1fKP1
KGo5r2OuYXfkZTXguGJSoJPEx0oR+mpSd9O6D5zvylfvOxILteiLAuBcwLqU4EBh
wCqTPSb6VavUOye2Sd4+avQUsBaBvIk/NtpCCQg4rD3/nSmpzihBDcmxZSIefgPu
3A9QMD5fmfIcY8f0ySi9e9YWE6v7U5ja7PElElIxaAZUXX+L043W5kIUbm95TS32
pDglG3pJtthjltt8PIU6scNoojsLrnvtx+ixfHgc/xDf6nzpHOwrP7FodfCI9Yo9
WXWrnx+sQ/EvPFzMSgKAuxY9Dogw3lnv/Ri44X51PiK0Enjy3T2LTRcoyymZ9IY0
Z465ROt5Kb5FFyF1Uwh8UvFjfGdKaeqbh8D8xHe3Zr+TXj/KEOd5Ye8bp7GibYeJ
SHf7E74EA5rUfNo9TrfSmEZbS9l9Xdcs+xl2x3ZTwzfE9PRVzW7+c981yXQ9KIly
d14LlUe1/QP7xbPHzlYEBHM3L08vr8UYfLB28ZpUBRPIm/MkDzETurNE0nJ127l9
TX+zYMz7bS44uKWM5+fCrM73wJJFsMPm/LBwqNuzeiF8oUoVD8tuOYe8X1dio7HG
ocAIwBYVf94hsVVAfqfSWZaURNQ/huEYd9Rpr4RgDmlHorSMi91fmfJ+1JiWGxFm
ZaEweQyy1SDeROPymSOwjGaa32Lzb9IjcJ/hNYrdPF4Epf30+5SdiJQ1fGsSacR1
myGW9N2h2iG/QcIGhX1Pt07BnBHZUqt2M1iy2gEMr7HzvVjaamTZ1p18VxttM42A
9a0mBnxJdx5O7k7BdYUvxMXFiGGevFcY9AkUoZIF3Eb6dGMA38D6YAO9z14aKq2d
ZJbiZYa0Y1DoZo2NYR1F9F7itjMaAYWjCHy0Qy1t3j+5F8vJS5vkV7LwBaI2pVIL
eJUjWWujG2fJ5220kdm3fF+0tQYk8w+BOUCXIxOPL9kZziMZfZmLQC+l9kjMwbub
i7c8Xn/5BNF92JQN7vgQnGrs1G5bDdeLWSEb2ugXuP6TvXidrxxQLJS3Hr0Y6Xhk
EWlXRh1kQ3MihtUOGNfQhJ4QT+RqBk8WDAc/pU9JJ0X3+l8MmkZx2xjfxrQ+4Rbn
crB44MihSS27Wd/tVbX10cP3NnjcJN+XstKvdR7qrmeXRigEuA0xbpCyxJzbnCpY
iM6ouH5VQrH7KrwCFhbAeVX8aT2aWItTIOP5yPPIsvPR1HTxfecLcMKpW+Y+uQZ4
fKRvUZAc6bZSJC98TVGzk/Jb8b1mkY9dxSlQwbHQzlICurk4nq+ckqYFFVvuX4lS
uTXKr1QU0bujjYJtf98VyGUbHLjV0ZHbu38QCVXj1NeCp7lBKsf3cVSlSW7i7tjN
bYnX+SnFppPH+U6qsfOIFEH4uA3P2LnWZo4rSCS6ztvVdh7RHA36k4GCZmV5m8p7
ZELEn4oB4DKvDkbdzEz280yYj0m5rY61vGIcIbjXTU7SdzRgcoD0WPkGrFznknvK
D3ZY9rVeFdn8h+Ljr8vYCTXxqAy5+K4EnV+UINCv6nKw3CFelAMKfuwY0Dd2W9/A
sMBLeAWUMVHzElVQ7HFgEqpIXVhkv1i5j800c3lKo/lwg0VQ/Kc99KEqaDBNMA5D
Bp3RufrKM2SDS62RvtyFZQ==
`pragma protect end_protected
