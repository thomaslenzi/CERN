// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:07 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oU3fmW2OUfQVzvsJVb3COxzVUa3YWzafCxV8H6xk6+5HJqeilBCu22M2Gkf+nSoy
AIqkN9EXdxi+xaddHes/YMOvpgx4U/Z/ph7SDyRy2l5C6KbMHd2vGyrHmKAERBWG
3FvJqE0s4ebNfZqOzmZI0KKJCZBd6CRbiUYld6RY6iQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8992)
OE1opKeb64rffyVwa+VYqR1ldHiZ9qIXXAYGxzFY/BJGLRJQb+jwjR8a6m0oWwsv
j9lQIsQkP6s7FdGexBV4TQxsT0cQxH/mdKl2h4uLxEAt1unStt4jro9Q+0bLg/wS
BOCeBE2B6Lpq2sgIQSX05dTjY7xF3gakDggBFhGEgQ7IHxYy52TG4iVPiMiDNh5V
aSNe5seJbIy4sZGOEb+LTy42SQsQMjSZewveMj7yaAmuo9KtW1W4EUQKd8c72I4p
ojn0D+nG2l9/1GHKAiJgOwEgEYyZBPokEvVkPBxRAuyeye2e8kU71Q5t1YwS1zoZ
IUVGTCu/jQL3vi6K12M7rxggqxee2tqew5aG+GjGt7Aj7dAydgvnaLt/89mgy2wx
Tze4vbFAv+9j9wQz6WybzYFDoDGZJOCfEH79WyAECp0IeDVGS3DSrOH+N6ONRT4N
cDVKUngmrI7HRNwnRfqBZCnQG6sUyAau1tJleOjXBA/c65NJ7OpjjdqE9ZvCmEZq
cLjHL2VjAaEqnifm/cuHbIctjvCKn7nVCixcFW5LbJ4ngMhIyw9if8jIxKcMNao5
AgKob7VD3UqFbxVcklo68ylsn27DZJS7bZFD3MsCI1A9ZBfP0IhiEnfDPVwnNmNz
lAEsEhpP6vcRSBYM3cv2wqY0SEnNKdwg3K9rhe9T3FHMULbeLADJOFmWcxhbzSyC
Hf3dL4up8UFj42iSE3AVPIIT4FxzdKeWFdQRboQI/UbN2UIpuzkFe0X0gEEz6VSM
7QpmaTIHzdvvYXVWCloxEVJy6oLioeJVTPJufvneldquTD3tUf6ANlZ2tFwIpE99
jxRCjPg3rYDHf9y6K8nSgdEocIbpie7eVjr+kTDVVszLukxZF6X2WdqlRopt8wJF
Wtr0bzJUcJSSSqZ2b94pRurx+SxKd9m9MQxK//2Z6liblDqmvZ5H7w8V4HeAuQLY
V1GuA95zaALIk7koqoU+aLoR+p+al73621OSiRe1mhancOan8VmyyJv9iZ9H0gDs
oF1MrBRoYm+dGKzNXWy2dVooAbyoB6LE5g3+U/RoARpmgT/Qp6w5bF8NX2MUQVLj
pjSPlNBljw1FM0/grh/HGI0HmyPu/MTdYLsueOppg1Xi3Ld2ROB7AZZyxXhMzn/1
9euANbOUMJkU0AB9fiTuCRqPQflHo3H7DTiU2Vjk8KD4mUCKf2rvdfnGwqFeAAUW
TKZJVYw8tNz8fjecOkBb5XNnqImtMaSwnw0k0XLEF3xq7D+Kuwsc8QLPx3jQLT/n
QqH7VtQx1hK/6kLbadkxDR5ePfZBw9NAPhdvncoRIo6ZQz7wFSZUF301XwVRvAcI
6RhsoXUKm4ApnAWX6wMjIoHKMYzK9JU7mz7aIgIP/Yq1xQfaft3m70BigpdFfFNC
H6Zw5KZUVSlq0oHizXmUh9LJsc0clzvHl4N0l8jp1EsFc+Zazco8Szz+jYydTkvB
0gfvIWwJIR53CyZMUws7xTtU0OIFG7FehjhWis5AX9IFr2+vsDArpknzrGDlgqDw
Ycojzb/w/PvHk6Y2CYcrk3lMCqSEB4VvaSwd8JIeWsWQo6VgTo+zt8XumU+xtXND
ZUZOPrZuKi543OViTctporlxZKMjbgsYfYTjgQ6UrO37bysuavPvjSxh5Tv9ecai
Z5Ylg9KYrR6Lzd0uROpSeMxWQyumM1eiV2Sa6pOTLmo4CE/YPUHATJwG6hPMeAcN
l99BEfh2Yw/kOjWdPaYnv5JnlNBxIptBJbOE/xt4oOOPcGu0PpaACHmYJB39ifHE
lLaHPyxaYdZBmdyzHe5MDIGRSiEbniflq8OLg9IUJDVGZc18lepks2n54Zuz+Wu/
vixjSSqwMlIPXEljyMj+6ov87m9F+YrYTNkPH4Lk9DEeyu3sgPF/RvseeK7svkLa
PFrQohtnFJSMI5sAe7Fe1w5fALqCKzVzCoVURyB/Lm2JHj8a2AJNoR+8zR1A9g4J
SmJ65ZeXTC9eF8ctedP6mujvfJL/9rgDC3h5gNv2Fgl/Eugx+fwW6eWCRjZrY5jp
AWBFSZqFYZpd7q4VHxqPAAQR9B3P5ec5u+W23I3u4G7blo4uEkXJTfStTRg8cb8U
YqbYfobAfAL+2P5N+teK+3bmVyjCzAZxMc6F6YgjoRtaXYpBrIvUOBK++AfP8HYY
kYBAls1IOhPuHBb0sV7mY0oNuLJOawxF4W9lLAjEkn49Wa9o36QbzTlxbue28MLx
1XhFmpWBGdfoPOe2ANQsnlLlVZdZuNwuNRDHH7ES991fvoRaREgAFnVU0HMqck7s
aZG2oT+n5vaSEZFHAs5DXZ7EHaZpy79kKklI7nroBwBJFtdlhJs6ywb4G5JwgkNa
FTZ3kn8Rd9wnsVD/Tao6hB2GBsv4138QXHY7C8xbKvSxu5tv6gmYbMe7lbCuD5Wa
cJmgHSSFKqxsFMzNuQQGj8EeFIpiodfTjdkyzxYmSbWwZxlrmXIvs1kxjv4b3Pu6
Y+JEcDzQaO/0BneKSfGnV8TH+WBVZkfCy3GV8BgZ8EB9FgFbI5R/NdX4MjkzcGAo
gRinQkNhumQCobYU8IOdo8UzfgZp0WqzTBTD2OZXlVohX0SV7oTGRr/Pw/YborMs
LJ0z3gRymQZBjoL/U67fl5rfGWNk69e35eAwS2AWk+r6pTS/pHLajxFvyJBvl89E
V820esQI+zqDT+8ySCg+y601pLAh4dy8GhZi+lORTFrNwWweSqz3qamWb3afXe1/
2KbDR3VPzfOHs1SZBURVMYCkNPYb6geor2eI6aGsWtKc5+jy+EsLDDJfwPPq7wQ5
8CCFbNvz7v381e7fag8jFQD+3I/IDfa+baUuJvq4Pxp2Gd+BNE9lTqHgXpkwYZQR
3Kzt6wf4d7e7MGissw4MNyCHtiNwqsnTVAjSfRSZWAsio57xy4pOi3VEhRqmfZ7r
UDaUBhtCq4EmVIq4CTwm1WuYVyrXnztdK0wzzMzOSWy4LmsM/fYl283nf4XPOvF4
QrRXhh+NhgY6M/84XoonS9KRdJkOM1ex4enSCdz+46YY3AuxWbAJK8MH1G2tK6Bj
kiwl0KY2cw2TqIGCSuXJzl2bmJOkMTePwCVVd1d3yHzgpziMbSur7Lv17slvI+rU
69+pHJd66eE+ybAC1m0scTLP0jH+F28+R7UTtq754jABYxl78mG6gpa78FcTGbmJ
N5ntVVfSDbihjQm4WZcrnhG2g+mUjyczfohy11e/Rfi55+1PLxiEVQSGn0C41i0Y
j6hSqRdESVL2rkoojEy7ZZB8hEMuqVVLwB4QdXWvc7e14sXrMmCnAaGEcO09sh/K
Q6owvtEhZrYDfoSYbpTaBJF9UIaLxPVwibZiIWTyOaQZXtRyQLnlA7fhK0HeYYsa
F3L1zpqMNPd8y/c7VQPyXtwPlgzhZdpB0SeDxPV1TlAwNY5kxlWW42WM7DJyn9Wd
saW7zLimhPsGh0QKzmjRm6+EnDRWLyCCtiLhkGEvkbjKxUOq7khaZLfLEyVRqNlN
94+UmDdvjhfOVedP1cW7c/DAN64coSgkdAzR/y2BPv6gtdWv8/0ZTkLNE/fuNq4U
wMAVsW/ZxurnusXiAD5Pdew11jGHUFAjgn1luFiJyRFkp0ACBsuet4q5VuGPJO4l
c1ZfN+Lrm2YpkdZViG2gLBXvm/lfwjfC3sd6Q/gkPZLtZiEekdCNFXv97rgx7Ee9
NrQXbcsz9o2Cg5HVJi0GEOR/1dZBjRjQprqZV7BVvX7IaJYahZYoWcZG6Im0eGSk
CcmSdkObOQxxrPtbIA/Z72ydzicSBwEfFLIlIrFvIAQ1of63d4bQKcDejdxK2Q2Z
F5HE/UtDkbUYguZOaD3lYZCAFZYJsaLWuWaykNBL4J92s1Yd9Gu4E5DcRwU34aWq
yPUgFUfUJVLMXPa1zAyo98C9RdY4Gsan8yASZlQmlvPvKSinuMW3xBNHgfkLYvWg
pcmu3CfJzgM3Bs1Mp8fZ6d7HS0tbzS0ySK9obhinrha+9XEXWHeEyd07XNgRM02M
UCJBzmcOjPJMhkFq1dh/cf7L/6J/hbnRsfqdz/hELoHPvYwiz50ziFok7UEze6z8
vmM2JjkyBRvRSwcddiLLROZ9WJgvwEqNyecOqON3mWxTwW3J6maNj4BYtk68nhlA
jqxWTS99qb6W5BkOKq32ujLm1rd4Rn3FCZIj1ZL+/NfWFXOslRJPxvjrnasdf0VP
RajHPiAjW6td3LvP/5L5MRGGwkziVeirKl0F/blF/l9hULgPKeOmFB/ufK81wHjn
OyWWbSsdt90bbz3FwOmBIxM7TQAYEpo/QjkhIvvmCf+7wxCyOHKSPoj6yanDXvr7
g3/ljBjpVnzk9ZQ2XQ1pRXA5Avp8eGXuxw2RhzN+9Fv6oh9nbLGbvgzGStQ4Ydi8
ooYe2QVKXBnAJntFZcUgG6M67PcLJiOOCQ15tO6vVp6eqHCPGdvquWCyaTwPaEsI
bxJgGrwX+cma0KmzWUpZXIg8vpD7RGr7RANGUH02DBMwliO92WltcxRSmt+Yti12
xKb6VN/FZaaO6skBY9lHAOnwfZAAjSkgWHBoKcc2iEdolKdis/s2XfKFtZ53az6f
4JimKYD1EOgDTwOvBUIwcyFEEpFd+pBvtVZYBqvQxp897aQWxX4Rz875HC/RhKJU
vj3SfeaEyFPUN3WMHIBf+CJBCIJgED1kQeXwRkdgNBi6PsCfFCFVAnzvaA04NDlq
NP/aYEYGGGh8HG5pI/YXEivu1P5FxFLz+eqxdaJDLN10CrsSET7xpl30371Wd8Xf
FyuUVV9+0LW9B7u+INZN8tmxItYYVIVhtYHh9j7knoA6pRqPMYpKuFNwgboIR5K+
HGR5VI/mvnMtOigac4OjcGlZduG1YbTV/9xrv1vulZspw9lT2ycEgNOpEYTNcMqC
KjQQKRSNA1Kci6J2NMb2nSPTqU48OTGe7vm2JwhIMJdPM7zO3baQ7PUIvjSoGltg
m+niQaSS2M+W99O2shU1GC5Id62A+nYh7vZo1uM2CCrL9WRuIaULyR4YKc1WgMVm
qZyARLy6OyWpPmNwhVoUJ8+mPgpfW1aLVS4pr8jV1ZETY8qDSH9zVuhD/W7K8Jhp
hVt3nP9TXhqCSsZZo0i0PSfDvITLo070E4a829YX3+yPKk2fTIunVqv+Kay4j4P1
73dxS3Jffc5IORoaeQPP6UFWNRRcpGeXEq6s70YxCW9tSaB1DGBiQ8MXypi7pYOl
sNHhV8ocs6+QKE+wckYyEEebEbk2x0bpKuMsYZBqqVBWM2gEJOtVEpytJ7cLl6zB
F2BlrQ5ypMcOPH3M0nsSz8yrgSgm2IFQXgk2sl/q1ktqDwlz7XI9soVe9R6f7+A+
eH7i1IuUm+I1wRAGlgzZ/TryNYXvj0SDmvVkL1YGAJBoJ1//hY0n2zr+ssS2jJ9A
B4lW1gDVHqHHxT2xGkBPMCNyzcYp8vhayF5K6AcHmQxLN3a346seSL+62TKsRWAO
Zr2ecVNhpFUC4bYtYwf1KNRh76ojPjGeTgsfghKEZzviG2bPig8gqGijlk8OXPi2
v4JGyh/yI7KtBKk/sevZZF2TWhScz5WVDJjAPsxg1lZfQ4bXLTrPDR6d/sQLB/h9
5LbawwsjlSCoFsI1g8CvHJr9JJT305HXberztQuyr4D+l8z9FrJDYMxFYGv8kykB
gBTStJB7OGLLdAgcMpct5Q5Bf0wI6/hyEc0YaykeRt0cKJMULVtRerepm0JpPWes
/bLmREQIPZpqy/9Dh6ZvhFZyZVSCmsdMTo7RlgsdRYHNYtvZzbxQIW0Rkizi6ItN
KYaqrEYqQEtQpYaXSosxu/C8SHohGCrrbnyFjPmSEbwR3wcEzilkI6tKLTKGM018
4tYWbSD2cm8PXNB2oKl1DYK38wf8uOVA0RQHwXr3ChQ0NGgCw7bi4DAo6Ii6infS
6+gxTwyxWjn/VtyLM+iNRY1GAiHP5rcYdzsAzJYQS0CVe77dcKepakDijiJ/0lKV
+q8TYBeJJjD/SuFizFthdJfehooKuENMP9R91JoYeLztjpKnlcNspinJPsazMiXo
9FRRCOJ+mEKwCjqmtZmgjtb+PuSEvDNVJRMHGumq6f5HayIyyVXh/n1KCZh0dntX
frCbL/uyGwFbllEsQ5xddZP7G/M61A19hl1B9eUYHiqPKfB4cuY7IJK5KPg+NTRq
CjspcVbWA6ryCrLMFcVOBNi1JPMEECE0dqoOwRxjY15O6VJLB8t2s7ogm1yoGDRw
eOLSe/UlLLhg0KxCtJCRP9eUz8fv41oeXiSumZGK8EpuTMduiwrSSp4nbY+ENUGL
NSGLfg+2g0FJNgLwXTnuCCXcdn5fDO/DrZsSY/Al2BkEShlDdc+BzhBkNkEJBsFE
jafHw9BZfD2RtGLGbiZRg5pL1cbGLB64YawojEq5BsxnJXMlYiFO153nEmcAvvUk
31KFal6vG0V7TucD6TbT9NBjIq6P9bc5R8kyEqPZsEyXovuKr4FiV1CiMA0KUoMv
0Q9xdjzCP8s0/FneyPD3pd3HCu2uL40ORzy1ZcEt48NyZUe8xJHU2lJVCQZ4Mn7m
t1WXljYPa+GKGfqa6UROESHBc7px2lA+hZALev6ucViPwayldMBGAgGuUNknESXC
dvWQoDQmjjNkJHH1MubEesIuPXV7Ju5zGZXO3M7ID8/Jxkyy74Yms9Un2OrNoPGc
62uW6oZDvrnxncBhgF/r703ZlzqjpjKBbvUYeEZcUbRVlf4G7jh32SAGaqTnetYt
HokX1uYMIY1X/mBQYrvTTE5EPEOjgbZRjiAYMx9v5x17HuVb6PoK/yRbJZ57XjOT
/0K0vtHiqqLfypNfG3W57+rk8s4VVxQ099uK48ubp6vEIHPQeSXhdz7Agjq7BcVI
RxxX4Guokw/kvegcMfwHeJdXC6JyLcH+1aK/JGdkBd5VoSa/kNr8udUVmbOMnn1d
xFWZd0Nt1c3yWSYdHocL4wlh6YXp4+Yx+hDGMdjRz3Vcyd2fGJPD2IF9e0fFaeYO
INA8jGZ4/g5BG4e0vAToyEcR6OKcWaLbdfxamnhmfVCCe49YCltBeyau4Ls4JztG
1rBw0xhOPABSC8O58cqolQujykOoJjDZF+PV65g9yRSbpwrg6Ht2sI0RDDm3yB7H
0chUjt2bCdidgoGPJUeptiZU5mJAAbwNXVyw6fZXCzFVRvXY/p2rEatph0ARyYVB
yA+Nb1jf3/7UreePpqW9cH6F0yNU9YAf1MK2BcZoZ9xnwT18PsgvSABhP1KCAOYf
Vq4p1yoGi3s5eysagomS/5b/EWys6656WwFOjP7eZoaEY9uiGKLb4dltKou+/e4n
o/9ueTwueafwC62e+QAbTGU6SROc0PAiMdKn4CNSB4oxR9nE44/vBCYw2ZgCaun3
JWq01K+PYz8HIdIt0kBQFE3aUW2Ese7RBmasdb/r9FwzV99nyoyUukN6G1L+wmJe
AWESf5P6xkQUYFmSSYd+tF760bz7sA9KDn2OH/BMquUHv7+6hgFAarOhtJkIu7le
AlimJhZHZxHyCKXvIAZKBGQ58GJ+iRaFqqJP+hti72/FKrSZfu7L7+XYq+8wy3GM
RGoF97jf0fV1ijRLxReouB+u9AJUzazYd5nAiMadeXzL8pNyDwL592EqXvm1X5ir
afPvirCf72UF49C46/x6rt5Ewkl1QbnVWGJ8WSEF0ueTJq6t595/Kh+aFSG493tZ
Gz3hSXmqrbY5AJsGgvR1A5XfnrCHYm0jnfs7iLVv2o6s8blqvVBU5q5X5aCZYdyy
9OUpoKIbDb3W74U/Hcq/Rf+cc6AlMhgwoQSP8CrmkIu/YY8p2NAdOHcCiMUxl80h
msbk1xE/e2DjaPcv+1d/LsomOIsDrZjA4hOwUerfsHlH2+v9kOtNDNB8/yDsCQE4
x9adFNumFDAqf6I1+yCMA4cJmmjNZi/hgGA7Gp+MLH5nC/u8u5yq9wdgSFmh/AbL
qSHTlyeLfqDqNXyBF0hK3jEOUwFjBZmkUTlcBKlOaJ5hbncXmNpbUyzsV8zsxx+v
XCntMBJyxiM/4HwMngdjM22zj0BKXo4kK6frIjACWdB1D0qRum97WfnSNJ847ohc
NFE9GPAfUtmtXhDJGxnbw7tghV4vNCP9f01lE7VALoTHhwL+X8sAMQ/5ZRgM6vV1
42tGsKjV6plupQDBBFkQuzEi4Q4/Io2/YmOWZ3k9U2kKyDt2qwOcsL3pr85aXI8D
B6rLWqbyQ/B5evdwYlv0myE30uQofGJO0iDUN/givA8YTo8Jf8jKm9UmE9aYbr6/
oi07GkpblnXGMw9jVtdA5WepWUk3U5pTgxU4k0eXdSA0ITDAgxuCYl5nWtAuYUD4
WFPUOFXDfQ4Re7rIMGQ4TZKPQ/LFDq777BsAlr2njVcckEukIUkWE2RMxGq7qmFn
NtGsyDoDBrRI3UX16vPbw8YTvuWVvpx3rCoIfIC28zINdxtTUZOaJBl8kk6tz8/5
6JL7/jgh5/FfI43+SxthR1HdZG0XyFKXc/cd8V26we2BJsZ5ue6GRciRmmS9NU79
KPv7LuR9ZYyA712e7pl1TqeGnjaLeYdGldpyPnr4fVRAdg9L5l2isgMSdTxwn2Hw
nh2VaByHAQHB2G9usZX1GiDtG7GzOy3AYDvoASlORxpHzxNjHVoEcfIlO7kmCQHS
nFAkIq3G8pJs1239dnsgOu8dlmHr2BJUfNWuDmr440VaLvVpTod1JfNDipxGRqIZ
eF6dO6y2ReYbqbvBhY2p0/H4Sl7AScPnZoUZkT0i3t1KeVzM3tGj1xb2tK0IZuiq
c3dgQFxjqjdXJXM8F1xgEi/ZcsBw0c4Wgtl2rpZhVU03UmZXtiPj/xrDc4hfWYRt
cpGiX0HHWsBhqu1ctUds4XjJq0cPNl24EK1w3jcHd/KaB/eC2Cnn3CRKtceIy/yw
ryvSe/L1v5CE3od/Gn134vr4rGNtmv6n0CqiXKSTAjA6gmpiCcj0TZ+MKozbHjXZ
h253/Xxkrzp74IJQC3JIIsxiefYRgmTyiDo5Ls0EhXDFdIrqGayqjf5OqFNVa7e2
iKS7HOdQzPsuuVx5UFOkH53G9+hQXkViCv/Hhae6p+049bNoEQCTQWn16ZpfDklP
77TCRUTZtbfKDsVI0kMSopiMR+aXS3k0rapt1f4tKKVo1NRGyHsuUmOjUCmEsyFP
e4yQM44Z0awLWBZu3AzBuYOq2sYHLnJRJFvk/hzWgxCJK+nL6gJdPXpc1KDT+5eO
XdZQfXxWG0xiZDTVlGkCh504R7F61eoYGC6wdoywoQO3hFy1GkKmqKoBP6QIqm1J
xstzaPBaqF959NQaVzt0QgPM6MXUfS++P2uc2oZq0yjADiII1ZBmZBn1gxANPyY1
lNGNq3NWku7LYu2v1ccCgMxqDekUG+u3gv54inlvlP6SDlN/eyIiyxOUtCe4PEOU
z1LQ4MZjfSvz0+1H5dM2Br92EHrSPEfNkYXtqSNlVVND25GQKn32SKIQmGdcO0xm
web8n0P7pbVZPdM5P5N2Sh/P4QYButpcQYufqNfvdQyJXstHdhtOzL67I6gX92t3
2O90pseNcoDafnLEbcHjoTFK+4lqKPo1II9Pjtukiej9UspsZxsVlD8gimNuTn7C
quYvWf3c7I6U5u9sWtZAQWBO3kDldWx/GvT5FTDRnhYMSZ9DX7zb3aMO5/kNxu7E
SDd1BiHYaCrYB/zgajZ5gS99uF4uiOfAmzGstLsvKyifsTdezw23RRlC2dyp7rN7
AJZNrsrf165FTM/7gaWG8tb+UqOupDbP+2Tjd8HQxa6F1FmISvswPWiDecnRcuit
gqt+sWv4fPHZ5M/HoCASBKSsS0sSIPD9Nt+ufsyNFm5389VPQkzaSZk1slT50s9l
3VpF247bXyIwD4sIrIjGnnWIoYNH8cRGZ0Qap+NWz52tTFXFVbohq43hA5b7EgUk
G5Ajrt64XC9G9dcu7icPgx2khElaNouv7PONmF4g3P4FXDe4CdvTcFy0S3MNsOA3
RW13B+/pe1hm88nbuWpFe4lMLaRlhufV1OcnODbDsHtjQ3zTf7DXIkRn64eGglf/
yWA1FHXDIk2aP0vM04JibnJNZaPhvQkSFlfvuELBmP8V9voTf+Z9KqMS3hqetL5I
mrzjwr3sdspknIntlkzvZxLfVOjp/0EcEhJbVRSjC6dSiztU9SPRyoTp9PQBzG4o
1iLtgVwCK8JQ3Yr9qgqPzTV9VwrdSukcbK495kpWbNvIcs7/lOPc4Qt6Q0jdOsMO
NCgoYtaORdfP76PSxs4cfIQzJRypjb+0vnQZPL2jJ9yGxotRq3AkKQXrezqe7IjQ
OL+K9gJLcpbtBEAOjklBmVoJbY8RmQ0kQeqeuIu7ka1neCgOkqstRxu1QF+Hwg6B
/punu/N1iVE4zLtkXGg4Ogzkblnaxy1Jfk4pU6UEA6YgKuPS5ZykEDas9L5Y2T5Q
OyuhVcPPDwuy32L06oaF7ApwI6/8rOxk/qNERA2NSid74oHkY7f/2rDw23fGTXC8
g3v8sP5hEgui/PAfAf7lnnEIW7tRcYOOL2NeVy23EBGse6SDTt1oq9u7sMz9P4yJ
ytEFgeDES3jY/ayysjGM2tz0dsQi7j1KfYeZHWX3xo1H7tAEacfPSXC3D04RMV/9
Euzt575gNizcZyQJARlVq03YOXHbU5Ws9V1Kd/m4c+eejEzbJuSjSF9esXSr64X5
RVWAsnb6PCRGsvKGn1GeNiQ4fBeuv04SQRjsN9SSHyfhUVaIZwkw7xAEgqd8Aeun
Q168ysswPuGgj47oAYJ9tWTAlCM9Tqm678Hs5O28WQ3NDP8+BNjfRyeoKE4grIq3
GP54eg2LotdJ15daKe31wp6BohTpgp38s8GSUMWDQZM20K6K9yl0up9qtZf+rBXx
QJ3dxEUag96+KfgXhnOTuxlG6ZIbuRM1B4oVFZp/haW9VEQXda0xNYa0LKGeHap/
gMsrY0w902ro7rt2xTGu+yFcR/GwaSruYhsUci/CbpguTszFRyoeSTR1/N7PyExK
6H4oP3FAo4UTIptmJSlho90v1vWxIc99hZPp+L6OmJDPfcZMYitqXE2h1HA351x5
akK6EnHfRpTW66h0kv9mt1Kive8ujTieieREso7ZKl7y+iNz9uGZBCV5vkfxGR/I
oikMYmz8aFWw8dE8216rCJPnTidUgMHJJgvh/40KZC9vB5lzlPpWtqJXyfG9Zyuv
muOhr8mb6lKXr2rc2z4pcBbOqhPdWPikwq0KNh5MbAGMSpeyHQ1ypM26JTiGuYmE
/PYtsorl81/7QJw0n0OsW2doNpPtXEgApn7ub7IbqisvHHyKwWUtcUjDmR+Hjfty
/qhQGB73yQx+1MgTIVKcy546K2hzlkoKJ6H4cQnBDQy8kqwRFGYwtstC1CLDtgSi
QYPsfBMZjZoQb9m3B7iMzq/DPxqqt6Ppj0pXl9cUrVkqI0Hpc0ofwr7dGG6CRk3k
oC2Ap+v6S1cP0zsAulN8ytqjaDNwNrKd1Rrd6SfpnOFdNwy8S4L8k0Ib7JQ7VofU
uCR0kw4wrUbMSiYbAUY2snzjReJgW1ewL26Pgd4s0carHrYtS/Jh4FNgUdgXBs2W
uTU+nWXlnd65lKQjCUYrZJcDLHu/+JowP6NqXxlGVAg/ttqzKuySN6k5uf/rIQI2
+ko+vfjw18WRu467j0w+WyVSfscgto/WHNUBlKcUBV+4SvU6Xn663qvO+vkO0z7x
J9yoSgvWIDDSaH2mMiBwcm4bUi7jojXjs0PotKzvtuh2noChTDUF6dJi6kLFtcaY
Jq6HnnJsizb7Puu3libT6ZwdmbGnKwuyiHQrN94B/gFtsZPSz1Mkcq0+TvOwdJ4R
EvQ92WNYspnabHRHq4SpYhG74vF5U3DO02cLyf0ooddClLaohfvEi7uc53rnz1/6
geDQuwXKRVHxHNyPPBlZVw==
`pragma protect end_protected
