// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y1y4Im7sp31Ou98FX39ehcxi2W0EdDE+HCg3eEyO+e+K1hCn75ZBs3PifaPWTPL6
6MidjzYHWpZccXW2Q6JtszKMVEHd+YtJ/GIrMkfhrAUe4Q0Xinp2jbTlQpIZA8eM
Drec4+KFwqWjkmaWuaHuOEjqQiLt9QioZkdvHcUWI/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49744)
aiY4EMoFtbE02CtuPZaV8UFKH3hzwGIcvgysfY2OJXw5O38iEYjW8jK+N7Rm2gQu
Wa8Lq7nTaygiiP2LSWf2WARt6By1oJl+KSbQwMPLsoVRAPnlSIEqvGDnJFgrgeJ2
IGPB0GAdKDN4SAZ+TzSNyiLxMLTdzbYXxa5uguOAKEDoNml1uO3MDHDr1UajDnyV
Mazp4K8VoXM8IL0OmNebRtx+wFGQk+vsMxCNmFOlKHKI4NJYRXuRN8YddPrrjZ4E
USGxAk47QQ8WARgEiZQvQNYZ/X1VwhQCUJPxEQHMe/IrOIYBd1mKO0PrTyKhmHb2
SV1/Gp+MKe5D0mIok6FyTO48q3Ts69MLD777Zg1GLeuJT3PKD5j2NrU93Ldf6AgF
TvcXjMnut8+Q/Rc3GCNEnHJeb0p9PDOPcehH8RtQohLhsB4xE1XgjCMnVLCy3dvE
LT7GnCnQCETwE45zH63SXJmjgA6q+jYLJB4fe6I1Ig7ySFew9Zm84wkxAqlZ58nS
rZypJxrvA1KjPqNTBskdNwJaHD6DqaUCCoGiPyxuVlwGJwU3WZbiy40lXCqsl6yG
nBNOmoNNxGbpIuHSTfFMIFiivDTnKSgjyruNbOV1IwejCOuQj7Ze+2Sbhdr0QwmK
g6f1QVJFv0Od8ccCMjbrfqYfJLAz+BGCcqS8fw4L0Q2p5cDZgGbzEeJKncFUbC7W
+f+xkjYXpkaQg8DXbGCF9rg+bIBhZRyONJg18aijRHbFeelEWJr8Nz+u9r5y2eES
WiOnapNEhglDSXS+YFRzA0ax9cQqfYkihA8JedRMrctfE0wUYLNoxkeY7sxGtmWc
MibZ/v8QGtNc7+3IHlAc1wwv7xglitPzHsh7UCpZdNNdeYUUk/Mps2HCFZnZyO6I
2FcNKbPCTRhyccVqlb8SgWbXv2Do7CTbRTRn4hSuW0LTsdVj+8GoeuHoTIQP5uK0
d4AkSPdeej0hKCff53w6Rlr6AaoRIn/XV2mT2pSaXYnOiH+Kl99VaexLyoRuPQAX
snZMNWu+aGzdmNeuRTSmWpAEQhZNXSjOsaqNwgKSVs6Djp2/OCIGitOfoguBIs+9
UHHwrn1p7hR1F//gTfHKRcIqr8RaJZNtrIy9+hhGCfuolsCQuQyETxCyipetuBhF
RuWRD/v+HHQ3qegpQegD4ibEWJPZ1se427VMKTX3ejDb78ljhmB3+OyX9EMB33lp
+ILEv8EPoTWDZ62+CyVewG4m7M3hZAk3NccVg/lxu8SxhdGLAZqYT22iyZR+BQL5
AdHYCT5I9Hp24qyqyn2A7dpypEqu84ITpHYvnrDmoH1Nj2V1QRt3X0h5vsGpCSSY
kG/PsaVvwtnwC22UuDnlIAQpwVTQpnK/SACK3U4wZ4Q+d7BXDFirQ0vYcdmyG3WO
2cjIQCmHRwdyzrJn1arj4xp0AxaildmOmVOz9yoBk48b96Bya28Xq+hiMm1A4teA
6qbIHmqmU5lPwTxkIo/CgYjsvYYzR+nctCEsCFC047k1rIsQrAsQX9R1AbAft5+D
CvRscqTmSGZs8J5AqmUdDwhzonSLIfMowZ3wf5l7z8mvNApzFhiWpNqQdHuiEtjD
sqCHjyVpbvNwhwAeXMR/PePg+ISij2WGHDd1p8NPNSkV77aikLzQcDgUlQXSlC3T
/7/yFkuYPxM4E5fZlY/+xC9BfglwF3RnukmH3Mzopa3Uh+VNWfnoE8DFrSEy2civ
cy8Yt3PkkycN76lOBqLPhzyh4EoAW3zilTiNWw2X7QX0tQhy3sWanf+OZw26UhKs
mZsCYLXTb8EhGzbp4BdFw5w0paSwcuOFV2Naswd8BcHsa2HWhk7dYNwq0e2WnQDh
5/bdhPHHzQ2JWgLTBN5MRP5pt/q1Lh0hTAtDkrtPpl0sbvPp0H1+BDRyFLsjWLsv
KrCzKuGNJc9V5Vv/NJY9NbdnIiIyyCAoWeAw3kAHkrv6iEd1WUslawNt3AW1tbj4
Yzx4mfcY54rBOBU3ruyj0Ft8veTxUFh53oK23mvE5EksibRaFyVOCiFuRDtcf3tI
lWXIb/fm6WohXCInMCNB9KeThHVjqzeRgyqXTF4Bg0u/m9DGPKevjXJtvTUgGvuv
WmCNeMY3fWuWj1Z3zFpBwfyKuEAXPPsAZ/AJH0JGTnw033UZfsefLV3EWU3BcJRM
tQvU9mfisSp1CsX2RB4iZSVadWJrtY9dpXBuTTla0qCpeXWhSs0BifMKhnCEDsUK
JgCT8Pj46ABuhR5J9vhtjMjZ5Mz0Hu3/6HWYWZ4lM2UqE8zoJ9IlSgRRdv63tLSJ
P5bAmCOxRqDDT310OpJDbXTXG14YW8H06DIdw9ajz/YYd+Lc+G2+/CGEwiFIJmPU
edKbPWbQYWX0CbNeQTZefROeXK46AhmjUbGi4xrukw7G0eqDQO8HP79WAdBuweMx
r5nKi3nF4d0p5ICN6r0E7+PQ6wpn7y6ENjCyF/k490eUd1LHbevE9DgSvjeKzoyZ
mbHbk+eZxg3iTp1BnWq1rL+MTF09lCDx9m/Yv3/RzMR9N1N8SJTsRxCCg6KQxLjz
ggI314sCcZaCp4HciSTxobFaCBtuhJZ4mnghj2Fo3GGRQEyJK3kIXWLcCzxAZw5+
E2Xe0e0xeeJf/bPj5qzd082YPMsUBWdZGWEqwFpvdK+OVhsay7q8RFsq4EqQWLbr
et6q/yzHNOw3fM8rn4Tx76X4cC/LuTfVNT+lV9WTOjzspna1ParWx/0B3RRW9ORx
0BXcYAIPsD/Z7Mb+szCgG1tQC2Ly5sSj4Y6ni92AF7DKCOuRrAMt0pPF4+5OKpjs
z3YeBCF1aF/mF+Joy9X5Z6r/Itt2hN6yEZS9680EKd64nYm0XtA0O72qbblpf3ks
Qr1CrUqWBiWSyMyVCmWJ/gQf/aRQAkWE6h1MO7Ctj68iPvMDoxuUKVWm8Gu4lwBm
v6QOJpgRAJR55y+rlmWx1jYILmRZJaEnSpyyxK7hXC8tOPMDRguCz2Z7md2E103P
0CLpDIjGs+kEA7jkgnGLsMm7hhNiYscjYDSv2I0Rw44KAxs/p/ttFiqgRkkPeD2S
2wIRVvtaDcjZwdR77pQ4oyqBF/cu02De3h2TeHWIcB0yFRGyCSJzVYry1792ITPc
rGvKVG4MYXvVVyPfevoRI0WqGY40oP/Vi0legPUkueqMTJiZytUHPPUfwaTlUBH1
ktdSlwzuM4kCNcu3Pm4mBBi6/Oef9BMBLISxwpaeTGbKoRgzXgvLsu3VjGreg1YG
+DCm+mL/HyZw8ROolj4r7POlwNSphzIK/OhVL+Lxc8Ham+uPVVgQBUlPC8hhoINm
AdUt4tDjWV+9qfSI85p2psOXUD5j4juh5YTNXHti5b2i5IdTQA561mLFL/khgVJW
rFnhRx+lfZr2E2RImtA1F7y0me6P0L3VfwgLG0TSRy7ytAQA9VBIu92pEBK2saSS
6rEubiyeqe9FbjiNq6MUGfxLEmJKHCmGc+nwqUN47dTsbWakIAG8mcVGLimJl/ng
Eiz+AvLsWVNIref6cKCfTG1l+KK+xjSoAufMucJmG97ocn313huR6bjStM8AW6hc
0QqcFdeEQeyZa/w9TzDPSCod3ZbPaxRJDgmk3NVOIjWBUE8zys48CSHumAtlfrVR
9oUwo4WDPVb5uVbxuo0bmdQhHMNK7tyEG31EZ9ZB/oXMYZHCWWdDMxp/u4TvxH1X
3mZ6XGvL9SWUTFsUx6Rc4qjXMhxnX3RMSIpfTBOqYGuJQU1EOgluE91Bws70HLVv
x4ZkTagB/vDxgJ6hv7caIGqQCOb1oW/XRkiu43took6dtQbTUU46JIN+SRIGRQST
Sop0EW7uhjzjZnq7Ry6Ux3iTE/J2YceZujHE/CemEXB8JefAaKGdXxRvwS/NWURC
EjBQAhQ1WG4SBEbIK8JN2j14vGyavoAGWACLk+RwgLznhML+nXc/mJB/SX2iGHoQ
DDXP+JuS8BCOE6ZzOO1oNvUDA7t3NPMCuXq3D5B6aHINDiHVSy5OJuAQgcT8AO/Z
tLHA/GBRc8ecnHZhlnIHOuNUKgigXMUIrEoG9agmtAp6Ynvg8cbs2HJ3oGXKJVfx
h8W9M7Rpat9aFKAedIAtsTO6RyH8+Feyf9aWysE2lgWoHqfhicfp6XWJnCOgDvCk
zp3AQDmNiK11dZbj8w0Z++L6JbsoVJ0ORr7GDz8AplvRdccwOXUotBfHeGTRI8Kc
jKUQnKArCMKej725NhR7lvMUzzQV63y1mhQEeol18o52ALIuOdckBJtf8VcBEYIQ
AHieTY99YcHfYrD7AouA5P5PHJpbR2zUWAtiKxjqa1WgrOo0UF6MZD2i7YNrf7kn
PFjlQrhsfUqZ/iY+TKgPIGwmI2ob7ELY/J7eiPxVbxBR9xlsgHV0YAu8e6HJgSak
eT++ND6kb4Y+fREpjYFvnnOdW2xC8DsAP6Dekv8n1nbVvvksZ72l/4cTaETk8wzC
/e/PApDZpXr6BxMTVwmm/XXFJzBfQqUUefFmtvnFjmVXuOWlbre7FdlT/RP82K3S
HoqoxcgcLVxiIdvDo84+sRYX7FQ51v4TkZme73l8RaH2uBIGJh10jpHaO3BriW5T
oOagHdSWxUYcEEROoZNJaNfhZ5muUworZq+Fn6Eeool7Aa2K5Ir9rUbyW8zioU6c
xV+vFCr3iW7f25HC2PvDmlJEXoaKLIricWdaRxJs6a0RiAJm/L5Vg6ZvXRiJT4YP
7ShQZgErVNt5mH0iRsSMAzFk7itGNqSYlPHb5N4JXP4GrOkma7Cu5xlU2IduZxjI
tL4zmSokS3qOb9VP+VsWLsMs5nId5qR5NcDZk5Lq+Bl1f3OnCs2+eVchcNlSgRA1
IcHdseDeA/lctLXrM+AH9xQ1uN9Vlc+TXlrQxDnXXmGJO5JJGXEfHNm19xCP34xr
HfXNkGWjuvc0tFLESJZEFtpcmUgzeet4c4sJv1UkBMvLxdPw4OduZwGGOHpINX6i
K+L4RB06narYJFrd2bZR3dUzq6PlpXD47+3AtlW/RmC3pVQcI4yASUA90wV0frNk
nZrngAKsudLrYL6F48Zm8cSI59uOJSqeSxGeP8MtLWcDlnH9pBK+LLY8TOLTtJBF
lbULoqYlHZxuThcH5QAg5KE3RhvcBX+z45QGXCDt5lRQg8o+JUIvHkWIwNkQqjVA
664XYevy4E5+KBOkw98+xks9Q73UWtopicVgT2KGeV8SiHR7SVf7huYNErdKhpC1
NOqT3t6sBaUi9O/H1T5ClbRwXfh3efVNWH8AP3aMmcr93R4sD4oyZmJNfIXZWOLg
xOasCJsr4EIJoUKHZXiKZdGZ339WG3fs2mSFTHrH7yoFh/Noh67ks5SfvzP/GUPt
RIzeN95R92mzBxnrtWIQY+MbQ+7jUHW9GlKmosmBI06j7v+qUputyqw3gYqGu5Fl
TyF45ck+9K1WeswPMxT+haUgJbJBLTRH7NDdvq/molwynT9TWFNUd5rQHGoG9ctx
FZXUnqECXe5KGNx14HM3Ngj6S8uY5JeLKx/67G3ayOeKks1dQq2wjGlRpYRX7tLH
b2F3EYb+Unf+ts6ogZFywhj/rD1hRhGykc8Dcvdgme5SQMgTVTGUHSyLmkr/4w2a
w+IYChs9WSiM4H+1h6ZY5N/RcOlar0JqaJ789aaX/xbxxIeHfnVrC0iMNM/CqyRJ
f7AUN7qzY2SiCS9M9oFyKTLZGQTyIi/GZPa0yEXE4oAS78WSyvhciFP+SmzV/jdW
rnvyFgBKl0L8ceYzbYmr2W02sqhdrQBwcjf9FgVomzT54Dck580Li1XL0KxVKope
fYGI+NYRUBngdA3WGFalWdHCUmANkcx/FykGPYDWIAT7ROZLcubgqRkoYM59R0q7
pYVIQpAakmycgOOvoCCmIZLV1ZPHg1eQddAp1NG1AtZSTWUN3UL1QrduX0g8TWW/
GJDpitdyxmjebfTatWuV87GWenQuaRMlu94HCVX6Xih+iavhvPjKgjGRv85P0Izq
IHYLA7k/8GnZxisL2kSCbrDDSqPO6/pbY8XggVriYgCh+1Rv82VxoakMmOmLv/ee
EkqfrrlIsYHZT5KouNU44kIhmdwPssHxnLMzzSGHg0XBn0GQ2RT45RdvPGxjfMcA
jYBdXYY3TmqZU4r8wSsOJG5AtzhcHFVdVSHDELw7c6R5MM/yOrs/FrZ4HYDWKb3H
vKRoINiSdmlK2fHmNf0IKDyUEfOtoUUhHCJZQKFUUBLQv4xaV9hzoWVrC7uoz6mr
oMcN07NORoJrBq3fam7nVALrIUhD1lj8rbv5r5CJVZEjzf1+x4WkfItLNz4z+j94
G4sYL+uIDz9q+yTZWkHjSsU7zBJSFugkYbHI7mDWgHKRo+/PIC7cpWtR89gMIcS0
FjHgI7VMdRLzvmMCPC4uYS9Eo2lQiVbtL7QTlXWI7Rgi95XpWWsbC12cAAliAGc8
uDt2e7oa8fJc7aDgKAU2o1CafX7rfV8vTgt095ui1b8/iGOVugcm+3Rcx8dx/o7Z
3TfwpMPq3mVsR7YlFSR9I+0eAonNE7yCWgseSEU/w48SG1Apabs2Um96xC7JFpQk
EOEXbG0rZnMH9gzPR0OP9tRzDdY3twZS6m2TJNTed6O5e9ckOuTnWVa77Ukr2Chs
0s977TT6qdB9K0qXlntzJqnJ/d2Cdmvtbaw4qsdnsBsd+fcWjvjk4uriNBlTkLjR
EcjuIa9hHfVYkvwPBmw7NjD1JA9fpcx/f++I/n/GEwyOBfsBespAy3IgNE4gWTJc
bhLvSxpXf8tnqmxFaGd9mIiuS2EJT2w+5fEJqNjd/1vg+OANxcf57bo03zSpNuCe
hn5SoDAb65C8aeNdQjJEJiStaSSv56umjwCTS4zq/Oo7GNLjwst+TxMw2WbyBY5v
z5000UxYrR4hDo/XAduyCVfcEMZ+6rXkO8gMjYat/VyC01GjSfwN8qdQxAtmeZnF
KMiztKVgO15d0GY+mvq6JtIyDOXOXrkhwjH5pXOUQI2Rcal8eAF0VDmwYmkbN8h0
8vCQMHHHhc5i4kjYSc8aaobvWaBCtBmAv8Bv1bP+P5KVkyKGvsS8yjVJ0IxWPw5P
JEWXr5f56/7WvJuOvO8r39RINYBfdEyt/j8MOeDPspaU96nxrBjvxvYKG51xMG9E
fIh/4P3UbLLmjlZIaFkSl+HY10tAjCuRMf3ELd0UoxM+3n6PnZ313fUqWqsM3orD
Rbg4z3UGL1qiLr4/mJbXaHKYrMrTxqw/5ko0UoCn3Qmv0VAXcdD6qeOw+x2J9tlc
5xOkxInkCCFfM4GLoxYbSDNNgC/ItffnN41qEhriMDizgq6QtSSejDFOPigKOQYM
v9mHRRTWoPEVqrjuLuXFlf862jyu3Whn+7KzrCaTV6/q3ZGW/zCUg5E/HIj+5f6f
z1hoUs9mRt7eYEcABDxOFlye7FBcu0UdJroVwnOqqTdso0sjaItk43YKahijYvH1
aEegKggqcaU0owbDwKhDIRGnTXZ8RRl8dqMzMnNNeXWmF7dwLEw/lpQuGf63HEz5
8K40ofDkZDQlKWkHUU08oJ33C68D0r+ChLAxHjKKPCi8tyXww4C4uuZqRh4L84og
N7MsjzlILNbWWaD7l8br3Zu50CAWy2qbxHMl974XpxBTxuJlBZ61O+WTBYUtlUII
iUcYasteeT4MP/t74OjRT1JsGGt/Q0NCjiCsvQ05vuOgUYkoacvczK9z1QqYCrjU
QmANDeyP7YSPOz03RcPAovZqfb+abhlYEVM6dT7yrqcKhCrDThjidNNfY7rnhFN/
C9JZM867Y69UyuNOSq9tINuAA8WJaCLiMHeqD0OjXgcfVQAZi57SSZi3rDAVjOvS
ebJcKHZxy0lz5JHeAdz8VNGn5f71C8xp61Pd11DRr7kXTLcsh62mIQSUdO2SZSw0
FhS8sANZLoIC06k0Jp3Ctd+UmsQ9UrSNwktB8TuH7HQUNhdbYmUDMkWKfjeUZ/Xx
QyebB1hPIEo/yGOUDOw5rv6DnpUhByQItnCT8P4uVM4iIfJuia53mybWDN0YWUmx
r1XnHjM5rzf1J7aezgUJK0OBN85gikVd5CcBVAk1M1QEmlydGOzcgoi+/j7RDuoB
50ZxgjVhGqGYWT/G7WVGHoYZ0N0D8pVBhNq296rsaYgalDKjGzsE029YgNTEjHRq
6hd3XMPYFILXplNryYYiXEhsYbBbFfmOJNiASHzyRIzmuXxRVKVsqVVp0KARYwdr
+iUjDF2KMVGtNu+hHdstCLI6G8P65u4VaG1w208mSDfDGhpwZeHqwQBrvOByVizz
ssm7UcdB/a//nFzW1oKgnbSK6y+Tt2k9pEyx2UpeFWvQufdqJUGAX8xPVROpDv8G
ONks6rX4Vdr8CaqbB+oeyBh5u+QwPTytMMXXXk0LyfM6usGzP6CN1Fnt+9ym3mvo
U7PEEKhEfcICHKwgrKjvLbr8aKmS8ETgqORQQhgaxfaDYYOqw53V+7YlwWk0sGu2
5rAWyNKm73E3TWk692Alln6mOI10Odzw76iuFYsW1W0jy5CCUJWaLm6fC0Lxb9a2
eGUmns3abYy1BvzMrcGIx0g4N44QmCuEXggKIybMKjNHa+OL161+EEzRnrzOR/7T
7wbex9Jdns1twz+uB1AXtJ3Y1zg6blGEIHme5Rl+kUq8X9aTrRGwCjGMAHpeKLXA
yRTHlld6hjZM/6zuRI4WcBTCnVkfTdWWLAU+9tGnzfWz7xrbrd6DI7MGwDbYoJtm
wnuXEP3bZJK0zY1kgvzgDPKCpTMx7s6m6Dvr/0wPMFj4LUWPYnYePmXlU0KxijIL
BcQbznvbtvi/otXzpKyYxTDFPAick/rBkiqlNZi8mmOZUo0G9kv/ieMteDJ2ioiT
fQNGNp39mKH8NwNxLmC7MMksbEDi5dFsAoWk9d2CaBuo24wUFpBrJQB/FwaZVI0E
DHA1b0zuPdnl+sMdqCEn1V7B9z+ik5D77QsjjMxNoKOXPOOZPfGsWXDz5Z2l+dOr
gW2tq1k3LlaTUii7J+RH0aEcy3G4bom2Ggkt/Kta6dbwIRPnzT3TXwDJwb+avEf8
V19vudyJrOOUBn3SStuYFGkTTPEwY2b1umCxWIA+tGv45txufVxBqJvSMfHxM8eE
kGBBynUhehb+tqBOnX003f0ZJ/GuFIO5guHNU3rys/D67npq2aieVXQ6vLzkCu5Z
1lH8JIHmIaRtJskxfo+++OyIsu/ktfWhkLrPrnPP1TksS7rr8oTQX7jgH7IVvSun
ykryNOLZrT0gfmN/L2wABZhMTgvXXt+mVLDYfFpbjJd7qRpPtGtWRSg5CF+IAEg/
6rCrsD52Jc+hGSaqWe9oLVUD6oVgzynDUvuh6KVts2TLs5pldUB45G+FVxoipBWp
AH8IHrNO5J2NykyNHxD1iRRoTx7cbjSXRbq+xolMaglfN/Oxk04kbqsISHRNtc7u
vbmrk0Cq4G2Pg9vjzCx2TEbcHtxSi6HNujrNP6Ayt5NyPJKJGzGHJMkie+7ykDxc
97FaDIeOigUM7X1cIUn0Eb3hJKXqEG2+1q8V16ITd2dRrTohQLlXN1FtSN16NF7c
sO2+wZSAuXNUsH1+n7nUrYKdNVSvtdIrMspTiDZgIznfd7ImArU8mzhhg5kzKlk/
MHm0344DIBBrBExy2mYhAYSzbfJgiupfiul8Y1ZMZ5sQcNXK7wFBY/XSHW6BQveb
eNwxkAvnPpmYmjrQd2y9FI6pt9+iTkPEHabihbGQanZ5XyR3UwmbUW7MH3gna+Z9
eHHX9hvTKID2dlr7DqXHdaE/ronPuLwMIZrZanM5zjiYCEJF5K8ix3EVgvpzQ7I0
5DB+LKd+ZvRnOr/drBa2kKn1mZeSf/jvh66j/KnYoj9TA3/HMUgK0Y6XJJHR7zVy
K+ATi4AMZzDvJtUY9bSV3frScL9KmpVMurT7MsJsAMjieoshe2/g7RcLvSaPS099
6KXWwpMfPWFX9VCNSxSOT7dwp9QPiasFL/TuT3qLbuYgluViqaZxgZ0KOJHCXYGm
TfDr9JiCRiQMEx5YNl/3GGnqJVSgcb/3Q660JCvXh26XUVr5vWsO9L1u+3HLuqji
mK6n2zli6prIWutWSzYM9+relAjUjf3hVFEHL8yt8r6wo0olTxGdCaL/NiD9ss35
PtQaxGqGSMriCSBD+uQhbKalyFHleXqN29KzMg4rf/zb1vS81+nfHkM8xbvCm+qo
NMC7mMQH0LPkL9HXMjg1npo1REn7TaSx24ViBFoGnHxS1nDmp0IusY//vS/Z6hWE
BJotvumg3U0ll58ffV6DESYRRrkih3f9aJgfVTTR00jNbEiB+AVfeP/Kf8VhIwD9
Czj+zxJvd2jyBBi/52jx1hvjg41mE+O6QJGuW/48AIjfnhwkTcW7+MMj1TTlqrYT
fsttTKr3McS8fBmoBM6JdagaOkqkE6SM8hRQ4GtW4acljJJ79t/dr5hUPnoQclLS
X2n6uMjVDgRNfgHyR/og/+NWxZZ1K9HaWVg/Q23VmPaic0UbFl4Ui45kljcbIjER
vdxvQRJIrmpnoDL7OvIC6yxFCHzBHe4v97V0gylGUhwV/M14kkGfa3/Y06sQ5iW2
nVbH71BbEy0vjsVL+KObJpcolCj6hxovtwqV/63rHNTw0eizx5IY6MfEwbsdGG0O
CRt5nu8A/3GcaUfaTZxbZ/cahUA3X8R/iDZPfbNShjr4hNHM4W/dmbRwNHKZ2Ufu
FWNsOcMULSaNvesCJ5LwgjjIJR6utqSMpEUZdwODKV1bSNzR06IQDdUeiOoxqg38
C67Y0etgWIoni9fy8ed2ncyqLeG0CBBmELDOTmGI55n1rroQl++f2xZ7vr3RAwUZ
CFvfakrOtY9g0p5ybpO7TuaaJ04QD1/OvyMTQiYCxs9tnbGkGLZn8OchygNDtPxT
MSOJ2K/RtA9zFZyDhagQhVVr68JuSg8RV5h8fF1iDpgU/UDs1qWNIhL61Awa9tQj
+ZFxjVEQ8WKbBw9aNgXDiwFSACvcvFZ146T9mewGgJqVh7b8gSsP+KKOW6uWXPGR
ma2A8bP3wN9Lw0b1cRwdNLM9v1V8tzq/R8D5dw2tiE6wyGmwjMhz8pCcTdrjxM6a
FyKoDTXwr4yUQbdPrj3CWn+N/5QOWyvWFcKwluuLZutwu4r1WB+j88g+gzQRVUwp
2a8CAngAKJxjhEoQk+bRShWufxTvGEtdSYjnH3l49DnwOcb6l38IIuupnN9JaROw
DuzhgrEOJi1idITPqwUi9Sv9CbO9QdG2fVUkqLwfmJvjDwGkSjXxm1t/OAgBruEB
QShknCRNDLor1ZwVukCPjcKsDdLdmuH0qWO3DT/NUYh+HgEDR6OmhIEI+6bDjbTo
fO24/kR7Ijxid6/vY1WfcDC7yCL7lEaC+bJhgz123htIfXLjoDQESqtnTnpr0G7e
AVPjrO8ebmA95ZVTYiZjcggkZCMGUiMnc2jZNuCWfyEH6NY4Fnw1MLoF8tNnlGmT
4SOXXQY13Rlq+eqq8TFP4uy5QQ4dVrEl8cj4I+Spdea0yXwUsQkrfF7tpEp8D9AT
k5X3vViL7QFFmp3Ob4iyafkMx1aDRa0j5c/w/bovKLKdyRmS4/F1E+OpaqnrJtv9
7YEaLbfCvXUX9k0s7KpYpJIf8mXhijyK1KYO4NLY32wtEM57e2thMWYMJWupWEGa
8x1/sH5UiIoLUqwnw0xBvWOrlbeMAklSM5cUdG/Cs/ufwgYPJG6iQu1qRSLghyR4
SWWNIok64ZbGCkf3oV0NSLcPYMI1ypCaHy+SoRVBIVc9EaA+501cAeWl9ZjzvHjS
SsClGvIMLKPJDL3YwWkzY82p+BrHUp6UESm3bAeXNmEjU0jflx07xtTKGuNI9t/D
hRll8VGx7dFylp12rHFXPUvA+WkN69JqA9NK39bJ+Jvsvlsf7Y4Ivl+5Uvr5qJ9I
+JSJivf8bmvgbmvEQ2AMsmcxPetyAskeTO4oA5fqjGYEtYoWUav6LLqpR0LRjPLD
r/9MvMIAZ7NQiedbHk6j2h6nrNSKZxMPYDlP4pWIJWTbuz/RjpXwcN7ghnvCg4o9
HNf5a7xPybD22lQA23OUoHoZnopHWimbBAnfXFyer/fV/Zj6SjqD8Od6miTphhls
35pkqPdAmbDSC1UPZSNDyp6Dh4fy9OtZ8XmjfVKJ1KpvRRscC6EXDKNzAkVMpOWC
G6tLYoi8tC7x/HeC/44GYzhrSLqk9NiN1VXSEHNBQMQ5VBo86aLj3+R6Aa7eDIK3
AbNQd85GOG2bZ/sZapWqgB4JIMMH0rr3kp58TMrfgoIlQfizAZyF48U7OAGjd0L8
If1ieHR11l1uta+T97113e9WZ6fiPygPZOzcv7cYuPAtOrTkjepbqPYpk6FCRWdD
ChL7AEelWXfwGTWh6x9BvT7dqU+hpQcU0TWNlCLWNl/+7bDcuAjZJOHEPgNuZjEK
fVLB3MifPmXvtRF8mFXSeDvTLO5yOGUprIL8MIzlNseHj2Z3ypRsQI2kCaoSa4D1
bSNC63wt9yfW/4cEkpQybNRasvy18WpbR09R+a8ypg/lqY1Xe75FP69iGqBMnsH0
vXzBdwQxGZDoDNIwSbm5ZaMyKle/3HZQwekLkhDiKgKXYPFGiotxsFmS22CsfyFl
cBq7q7r7Sd8IHCOEuZYBoQDoCRRajQ0g+VWT38LKfDMZPFZO+tVcFiXhcb2I3nxV
adzBG2TWyFLK43olK+n7pJKmWw4QTQP0bK9+0juyHT8O0k1DDJTwMMha3B/dkD1V
OY2d42DcUtq8IpWyyLnVIToZdsKoCxxcV+Sc7osKU0VzHUoJwJEzGzabbKhU3Qjd
6LqILL1K0fuGoaSt4a32jbYNZUdPwf8B9cCDYwkD3iXPSdzkWr+YwFJRCFE3hhUz
4+Yp17jh+53cNsxiHwOTh1g4SEYuFVADdZ1C5YNN16vYKDZptxMZ6FQq/jP1FvR8
cXHGDnghNnNcad/c52Z8y4/kBHxngZ8fAA7QRsbCvi8l8TMLJ1ZL1tUC8AY1zc6z
PcktiKp7uXXodILrWuX+KyGV7ItMIhzSrU+zZUJJp+ipV+JESKev8JyJThzonwqm
iBg1cd/WwzNcqZ7TXxcGPP/ra1OSZNpj4z1nhIw7mnzEMFdmov4vAy52acwew/AX
jS1ZACVUrH0PV/pOMro/w1rCl1gJCBxAMuy76bcCs7A/mzbP+1EaUm41pxz1nLL7
DjPFa8mCjx3yZ6tevpE4wJsdAXANGKdxKSVdF55qrZ0TyBALvVHa9unUKAlyiGw4
MsH7UAXkxGOjFKQVIVdWy96XD3GY09zXPJnjFByINQkJDLw72VeC8AKw70JOCMN7
365BhF7Dear9zf3IPn4N88YPCrZZNkMAeSfAR7+T7ULMMpkZniDCusuALou7N+J9
POYCKY4EgT3C7t2nYLtNd5z7P2Ral0imfy4vd+lcsTWGhNMBkt5EVusbnFQdTHis
iH081RCpgBmRDjE+z9U2ITiPAk9BK+6tJPpp6azJIaKNqCZSBajjjdYbUqFPGiag
OQe9aqm0zvD2PNB8FzpzUVgSdhxn0qkzIQ/HtWthN/LeTiryDYH0mTKoeQTHtNTN
rQc+t/hh2N6VBngWJdVp2kE5EN3C3+sLC9l4Wbx314FplYWRlk+c8HpyGJfFopko
NyflmgxAaizfuTwDa4EaTjHnCvvCwgvgSI6GsfmV0nXKO4krujblpLY2d+7ZuED6
/Uyfx3ko2F4C18e7J3S6MC3v19yt2c2c/LKUkwgUl8AWAgaUc316df3dyREGje1N
/KlX+4nVhixxxgiw0mF8bLoCopMCgI53r9RWvI1vy4MD4J73G8h385DuzSjDGx32
sq5aC0pONRKjn6s/v95Drm1H3Xu8Q+iYCRpPvahDB4RJj6ELm2AZRxwqC4pYcfAN
sFuZbsq0yoGy28siywXa/JoYz7itBA3QHcOpOUtbik8ogN+a9fZUCAz55JtnpajD
jNTFVITfELwPDDLrHrBO/W6dJBP0+k1/sRwgwDLYViVvPkQiEv2dOty3jcEtsvUf
VOumWnxm5Yd5JUWXS6wzRsq+b56Re+OB/IKTOu+DNA/8ojkNBsXl4ViMSY1IeTV+
bmpPqNSQf8FDtLpDt1UI2fRjvs1/Wgw9c4yvF/kOOijImEQkJ34oAE3kKJ71YAJp
6sggxCNIqjRMS4jG0tyfBKa8G3Up7+rB4yhgbwLzzeRo0OPJpG48ZZxlvV3UAsqi
yMigI+0thx3+0BK20da6x6z5I6c9h+ogAcnOVtAByI6unjW4RW8xo+rOIOnKpXX0
5U4wr+xaNF+Sppu9dmrhWi9WFsOtFfZtvHJiiMEWwVg71dORn9LMLff7/UJlqRVP
pduBrWpQkjAf8Gyv/eOJ1tzQKxvZ9kjRmjl5UtpZtByS5UnYbetsOsVL8Dbal/Mh
p5KK8jf2Ew/wLWJMikNdk4tdavslSnV5PwpIrOiBWuOL+NzOrMlbbQ2DLPaZCkl3
nfz7GnE4TqniP4sEjp3irvE3oj2X0oHQAupMmTnp5UuPVHok7FG66PCvXc5Jphi5
gmXuBa6rcnerbs8XsHsgliMeetir0lTkZEDQCvn4rDofbgvUnpFyNMjVgjky+GKT
bcgJrzOpDZkQ8SvoCWrIfJh2Mmu/0IYvE6UNMZ5APXmWNrbplfD9a05/V/aBbh4M
sci6qwv05ZLxFnB8+46+TOMu8+f1PtygH1lvmIx/LyWxgVpwywu/JJZj+66RAADQ
I+gUrWNoaHh+rOiNcyKTu5zZixcm60LwkmVxUDAiMFvBTxN6k/0ndwD/Y4sj9bwL
NbHnkMrnoLkeIWCvhqkZ5u5866hoNwjt5Ow96eTLH13woKh8ww4gnJJo+LCMNQMY
myhIzHNOYB38x32uIxdCqEtuMDaHANJsFbCb5sG7jPFzZM2dIqjgXhRJuIeNwvtw
vCQBETP4c4LTnoCCrtYDrK0iBNc2E0ce60ScCKRM49lZqii76FMWiXFYvtwF/uxN
cFzfcpZVDio4t8SzkrQb//Dj4nFckextpDCCOi1Eckl7k4Ah3RpyHoouzme+wqyE
4f5lAB2smZeF4Qn2CZIQ9b+y65k/hs6drAGhWG062PzSFHvP1J1VrmfcTK3VPjv2
AXX56LTKd6hj3ocLFD6Mp13cu8tzAvdNFpw4NRgDqIJWFr8v2DYzySaH3GF5H8it
W4jcvgQGhhZ410enmTgbQuMNyrcM9tm2cSiO0XG+JaB5sVNmFAQ1XBotQfkFIEno
whsQDSlwO8GFhoDfVlKCub8Y0GSvjMZG/4pZSxGw+I0XoPHeSG0YctwH/OX6Gf6v
Y9ANFoheyEGBfndzUxp2nT6R9kEvp1Y79SdtKrLbps+hhNs67CU2fmBRt/WCLhd9
ipY023BfY5IiMKD3RkfCRmIHTLnobG4UTmY3Cufvmwk9ub7oiCcZEJfrzRvWjEUH
1xqMgOtdoDzGgEFdHVAZ6BFrfH9CA5Kexo2m8ICGLmviwsWehrb2bzFRRUKVMJpS
Xuvn94tk+YZ4oeoFaiJX5WR/oJ4yyNkC1xFlmfXgFkfcHSnMz3pzoZLTj2Saz0iR
8kqNh3XH5axeV4k5Jwh0DGgyHMbaaRsh+QprqJOjsuhvZkjAPTLKj8DLVu7kQwPu
X++8b/3kqdR7ijYRLfqEOCbZCQdpKTQkj44qiHg4+O1Ea/XAUKvBju1oYRRpiMIT
P8R7NdVME9FjeeL7bTSoCJ8EKRDvBDnmZrheSCg9FcT+3WmmdGziJo2vcsOF4dbg
evcj42NDhaqbRupoBBY8v6wBHUWWmGi9530DlQHuS/LI/fGH1RlZFOymfceeWtDp
ft2pt7pYBcmZzdjEsvJZNZx/ThaIPPRwS5ghJIhNegQBmUIciprn2Nxn99aMgzq8
ybByUCeUwYssoiRO1gNtlY/kqMSp0kBnzuWZQRnwArsK7iYUyBv6GxIlKigDc9OA
AljbqmZCjDUY3RMlLaibtVUFoHMBm9QMUc+xlB57hMGsKp6QbMHycaU2Lq3X4BT3
Gvfu93ENFnYEFXj/YQEw38CQT0pTFGH3wdpoYdCne6ech9nHRDzquL5GoQxUOuKZ
TVE5ofJynt33KAAVi9kDf6y+frAAzqhkS3/2shrOPKopS3wMHU+QcavArBPdnQ9X
lN5YZM4O44zw83KudEff+Ky/4yR8ra17RVZQTXVxW8uZ0KW79jBVpcScwpmZfDQL
0FTotxREM8Q87hqE2Ey+kPLS0Yhe0e9j4tFcferHb9tjOMtXVcoj/rowXNe9syoH
D0mhe4j4qO5dF/R6Zf8jg9Xs9MSLpB7CNqYZFdxoiIafGLbMD6G8BARxX3bK7iIE
xLHUeAjW9CMgzlKaPW1tqtOIHIF2i0PtzED8awGqjIXM/lcfELVlS41TSzNeIvTm
hdF5x4DRQx0N9Z1YkLuLxjhyHLfNlaWhX2rozJQBczRtUwOrUAKoMir564S3OaXy
YyhD5iBmp0K9pmYP4QszSsaX7GcNWIn9rGEuCZ3EQ8/Ds/c0qnqhuJWHUujgimTw
tfScpUDJAygZTz9NL92FuYYjor6KR8lbGZQgJoweBLUlXzNHxnh21uu6Pwz6iLHq
cbnpyERCx9i8IxES7QdeqYFan+0JzsKp7rA+H2iI5aHY6KgFxmjEvePesqXEgrvn
r8Ibt5z4nVtsteA8he1DHVRAeNWpLw70aTDRi4vaNU+u11Aea/RiB64Ihzdjib62
x5Lu4pdOp7huZDafUIQHwtJvUHtGwRhWUWaabZm5MLVYbOtqGIjL8sqhmMQw5S3c
JBJQuKnSfZ/ck418S9t7fLg6Gidh/UQzidbhtettAj9tEhUz+4yRbr0gaQ63EaAh
RWIOF6ReGFdqR6RIbQUzOQemN7YWlfSQnE8v6bWSG39jEPaU5AUXoTAre1T1SbiW
lMASkG80eeatcNbQlmRsMgZqJuapsEt8IwdPfLIYr3KUrHdwmumCbPI2NfAp3sqL
VGu3VSSJ/+tyiuHQP5AsqJ2aTZi2VYjPxqpIRcGRRRTwXvcMH/jsSBo4V6Jr6iGX
XABadNCNdqtRROmi1RM5Th5io3HvkVvXdgOaSEikBgjDpTHko2mDbJoWPMXA+E5I
+ksQZEuwvMJ+eeCXQyP8kL2HJJoJvWVnTRJttoGB90rfsAZGi1GMCHQ5Axi3WrPg
SZ1tOI+2BicOgfvVVZYlnkmHLy7+YpxgWUOg2iqqfmEZBU09+Phk0SsbbRLoOpbL
WrRKFa1BGGb8KCXXyTtKOKRvwcCWD7pxIHbyoc53c8kH1QmDekgKzKpRN/BFfT14
2VHM2IAZqWCinrAJNdLfukAMAbc1Te6b1/AMDXbbMKWC6XxEYMjAFj+Xk5WXYtZN
8hS2WurJVhxXBouM4eAm10KKu4ORnHqKPWT1SwK4gzgWxNY9tczzFteQoxjaNZ1h
yGwIjEHri38vNm3BZTJTLMgTKGM7CoECVxNALrb50yBTfrMK0hSC6lyWmfxyR45D
pcng4zhB9UhPPdHwhWtGjOGG1yIfz8hI9wsh5OPLdJzRqxAk6PuL3TaTnM7Uj3Ju
dDKTF70dYXbFLpKAGcbN2sJ0CSIYYRsOoP9g7UBSWe0O1KOmZhCyVkt7FLTYDOSJ
TRUjRvpp0RwPxlRF3CpmF3T0FIMnGJA1kJV5k1Dd/wfJirHTaRQXxlq85RXew+CZ
bXfuw7g/4qcKowl7VwF75qyVUK1s9QW0KKsP74KXvo7y2C87JuwDwCoCGJHgqDJL
xHCw4sg7abFTFKUiyA8udZzn+TTYPl/kmCmQbrClP4zcyr00AxHTIvW+5aulf3St
iil8jL/ZcomawwVcEudocOiZr2kBwfZF5UVR54PGFw+RgeR5Lq8eISvfcxamLE49
DbRiYR5OU2KyKStVcjZjd7yWL3SlplXT8DolLq3Hln90BWz+SsZbzwtbYVzbPRfK
lRa1vTGWaF3caNtiAK7VlPRN/lmbNpf6BDrLQlwrSnYtA609/mDlOU57PqszHauD
YhB6BoeDRdS3BXZ+jpeSRLMm/WERsw/WyoCXUh23c0/dpsiszTkjEYBGH8NGbeEr
wccRGt8w+dyYkzY2Z46sKhU5Z5d4635SQi/cUvquW0da/EUVue6myEJeT9yXd8NF
G6l3rYMl2BKvh7y4co970cxMLtp+sE9mCjWeXq7wtM+qjjhEePAApUxb5chlUeZQ
RhbxPb9FztuiophGG5aNgyi9dQlEo5xuhnMLDRw3IykUEX6J5YwRtFjSKwrVn1K1
uES/EsFUXdH7RDhp3G2p51zXQVu68NSW5cyJ14u5FzisS+W3AgJ5phJsV96hqHmU
C29Gi+6njonMQhHPCfcrx86bzB/ImPPXZ1m3Xvk0X5SYUDBoEDR+pZkt34UStgCE
of+fcX8IJS0IC9Trs8KKtvazZO9f9FT9Klwkx6ekmt6G/65wZi2a+xJxfxOlc8iK
07CNX+5pY7twPSwC9luSuS/rKbn7of395PDCK2TZQia/LK3/Q3A4h4jvt6MXlcqJ
iP7M4+2STW/5ww+6Iq1QDd/J8H9e1WZecwfA1JITmYjvkD93DEEL00jVOII6TQuz
drDjs9NMB7wFppuqdfuCAC2XizrXMVq+Ub3q0bPM2J+679/mtQNF+/7FawlDax18
V0ks0EFmmqYMUpP4hbw6i/QuQEEZcLoPannqgypCeb4M7fFqGbKpVDMZ3fuETi2z
SMCytIAvA7zGymQVR9l5to/yoZOU7uMsvuhubj1xF7CLW8GhTGgAnMuTZnUpMV+p
coQEJBEBUM4qo7KATjh1FSx7Zd6QdESGCKMxd8aHReVBTrsbDUmtvcqAuiIFad/3
djnVPjHZPRy3ls4/mmmbKd0rFDPgvVrbsvlcsYtaw5cG+3KI4xM1TFpHjRbuXC4w
OUkyTRUHVB3th/C1pVs6wmmRgafF5+kh42u3TqsE+Ho8wPpE3yShzdyuGWxttsPe
j3iQgVAK6bC9nM4PxOB7UeNCu3jsVxWdlVJ4dMlVIjrVZai7n9/nO1MIP+fsq4aH
OhpzJURumWIEGMSOyvQ+mTeI1Ttd5clL+ryX35JgnQ5FlGl32+BtDMaE9s2MQSUI
ei5nNMBzojbPqyutdwXqXa4QEXIAgcAsOxg4BVLULaks4XmpvLB2BvTHJEAylAK6
piuzVyu9PgThbRuZmFK/E73LeDB7qMKfR6cEbyMTDz1nqRp/Ik52dUfEKcggBD7N
O+UWDLWSOOdgPOrKqFmxXbEOsOghfcP4oswKwy5qkawH61Vjtwbw09ymMFJypiQM
r2t9oJuLFIzVMTIHL0tcCAOdya9JGwYYttXTk4wg2kh/pRv4IA43WTItQPrzYhKj
rSAkR2+Sh61stLNu336UiM7E5eFzu/zsFUEBj2SHlAVHOYfq0sC6XchFgB2paSGV
JBt4VQmTRWxXC/A3qlk1Je85furMgwwvcd15zIyDDXuGiPpYjdUg5X7/93Wa//Zk
HJqm0pC351XyPul4pViS450hOuLxNu51yRnWyCjCaMUzjdtqiqMjvm8axZSSpKH8
W1iQkyFrEZm+q1/xRz1JOTQ1sp3tsc2BPp45SeKdZfrzaVuyFHwwBY/qK9RegviL
hbSKggOp6uLSO/GnMP0bjbymp/4ZL1kDQW4X99SuObgFa9RUpnJz7qyz/hPqQFsU
wAy6xkAfaeaNTsr+ThiDmVHHqNqpKTzW/fX4nDVN0XLn87TsShR7OBFAz6d4Rhjx
bf7DeOWbxUIj9pzN5srg6GhNp1aBFIvxb48Ss+2+oPFqVi9tC29jobU1yZum5kDm
+yIdLohBtMoq9FPK9jrAfzPUTYkSVnFcbgnvIuqgeZEv5s18UiV416F+ZVrI1IW6
RzhenwFgDyi20f7en5xVKl1WfmcJANLeOy8FOy55CMgFhR+aaS828fOtlXFc35cX
6DjDxykkDUObQ2GsxXfG1Ju3eUCxr8jqiDDq3QATVq4gL54K7ekFkzxIxpOel5Q4
SjXJP+uuMjU0EEtFoqfnKJWrnlXIFol+tm++UxHi6n5hv9Bs7oWftIWq41geJRgk
ATXxKwAuzAQfhzUwDwnHW+PPp36iDJo74zgaleCzFcPl9Er/XqqBWSU13Veq7FRa
B/v1sdX45l3fp1oHpsY4MUsh4A27+xE0hcXl72H2X9b+bTFYoo8ddtUSe3d+UQAH
AGtdD0abNxEGZqoxxbU/PUS02jtKUt3sStzyTGMkOjmbn2ir7EjblvEDwn8q29E6
Spiv/ZOp6Z0o1LwulLyfNU9/CV4vnWWB+Xb+iHEWAjGT8Lc6N7MkN7Kf3C051y/4
x9n52mrK7JZ41kaMPVPcb8JTxRE1rQmbL6Hgb0uo1Qg21GNF6OTV0jYihqxWISJ3
Z6RW4SZ3kKFx09eGlxa7eyd+Y9cn599IIYA8yFYquPTfj9WkymvGjOoQqMqI0mq/
b+kpacrbMUhOlMDuzeSSRtdpyazgK8l7GwIBrucQLKI23VfFWlTiLu9aeLpkI+yd
DaeoMkgZSB51sKOZ7EyvnPTFuZT6OJWZlmqKn69Z583d7l3mzTqKyCihuoKEplzG
xukUglmPktlZVWcEiVcM4pwGr8ztEEUdo88ZoAAy9wpTdh8ND8nRnDsGrtuyEDON
4N+qHKFmb3ET84SNC/aaEqFo0xVw0XVRGCXgYYlUQKKiFBrAU3c2Ruk+aExiOnV1
sELEktr9kSogiBrzu7NO14sLQ4n85oteu+pwC6PztMMNH4vSBTw0JdILkKtlcax+
1lXGkFQULpJ5X+BNpiHQ+vRn1/RvmFY24pGQVKM7N+AcxyZPrKVDwgpi+SQ4WOtj
Kj+FCF45nS/djee4P4vOctiYfDpVUU9Nzv23ne7oH2nl3hA5ILU9MpRgzi8hCSOn
9R5xlRpPTFmwBlLG+fesQA3erI/4m06Kcoe4Cmfcw8gVSct6V1qfygDEUXC4PWOe
M99y0SWTGByQDOTlJs6L/q5VdCgCRlozPqjdfUnPJb+ySUxEMXBXn69VV4pYRbwu
RUM3WayHPAQCG9LdX+A04r2wvqwGMKU4fFBfQZrcsO1oan7SzyaRxBHXJyS/m2t+
Y+tVs7xUOAT82FzFEN4nJtolB7NNqhpqr0053eS0AT98kB7Y2EEQ4B97WRQ4FQ02
xyYXU65vjMEfXA5GgXKN3LTvrayfXbh5j5m0D0/AfKpiyw796sl2pKTQtwDemaJf
OM+oi2ewhYvEw+TEIVgZl+GOHx240azqSJIrU3GIPrzLYZbK0yhgUiD/BbkdREmj
XzUfHyxzCrAW2uA8xQhpazUDepiSOOKRg/CqKldpHtktPTI8SU0CXilkOdq9XNOe
PNMX8sXvz6kUAwD2Kb2Qm9lOevS93D2BZL/uuMLkp79kBcwgWYaxD5mLsZ1kx6xn
u0JzPgIb3Ew5pwtkO0bINpraUUgLq4atWjU2pMtzqBFVnhuEF/XN6Gl3IHR4CWKg
LQDvNg7E4FqsenUpDJfAxy/fMBbohbYODuQZJ1aok7eHINqDAMQWRI0gty2y2wcf
6jtW5+PjCdbrJ6hQEIhVNnJ40OnUVs/92qMiEgBEdHcUH0JhnivyBNMDWqaeHsSG
xA2YsPFjEB/t33DnSTaOtWKn86Z9ZOQK6Z7ipcyuFbcIyaY4WQC14u9pdqmf2UVj
mrL9z5EMFvN8n9wLPUqf49lAv/NOeIM2DaTIuumwYRP1rgk0HCNEehcaBrM/S//q
Ivu+o6gz/22eNo1led0GRrCLv/1odFSXlL8fGty9D9Ze1LO5fPJXqxjt9VtL/AU/
CvEH+LbMcziQsnVMmSce6HxaSqbKNktNIcls9K6MnXCHYonZJhIqSQxpEn8nOlwn
daVeD7LEM8bCGQSmrM24sv0RH/Jswllmq2wJhAN/bEKsBVmhnwHsjywqmOJjkIEI
7QeMYct2+qNWTdDtIB3ZXdRt6GQEt9ASzOpXz24OwueFkGPQAWAC1ArvCG9Phcs1
smjzW7UXL0fEsOZfde7alwlXk1W3YmtJ4hCrOszHaiwlNKE7y4Nu8shJHRcZC5uS
CdqFrfDZBJvVt6g7/uboQZx5rKw8oV4Ll1zMhvTLghre7NxOKX8sEnTBww3Rz8rt
AlQppOmAD55doA2nc0ODp+/MUdPuElrvEiKX9DpTLvhvA8UFZYnqX0PXP6o+q61J
A+mKyEX5KfWW0juRloE8iQJOnwgD8exnWax5QAYYi1hCWDzDeYN2gs8dd6882cah
BySRNKVwUSb3f45VRejzG0E1kRnrAgeb/HeSZyMspLmptJPW+64clQPHzuCqvV6M
Ro5Fv6nIeF57OsLp7gpw5UMV+XeM7XMrTpZ4PwHu3BEyNv7E8u4uQqb9Q3Lk5Bj7
sbopatntxs+eo8OMwTE6OR0C8Px5IkAQrcE4dScwQkGQLySWSBQHYndL8KLQH8px
xG0CmCjFsM43vYC9v0nC9/eOcvnXjwNdt78KN2hFNKwN5+z+8MyyDiCGvKcnNCI0
RQDi7a/r3q6yJgumtKfmJ+HQSZMKXPp74lmQBERoneLKuBUdwDb27IifIcl9OjUe
+0eIuAv8ob454fCFmOYx+OuXhn440b4ZMm+riGFu3tWaYoxxfabETrGflmXLluKZ
APmShbIdAT4cElCwofUngzfYl6SEzMq2HmAYAFxIIGnfSqQQ81zXJrk+72ltP5VR
IsOqJxxrrmbYxhOwQXvYjQKTsJoo56IdmjYDvTlogt24RB1Qx8+9L0iyd7pm7bdb
t8MWzL5M2XAg+8w6G4z0uSl4/1sXwMSrwk+kiMVuYQp5xGa85PzRqTD51OnzJfBq
lkYaSuAUr56JaxvdTgWeXOgUJ0AEK/ZL4X3dI/o8mtv58a0NRyM/cEBlEqYWE1Yi
fLUVA6Euy7wiNQWQEenuEBrNJdRF/6ELF/ay51DKrSKLwK/XsjM0lNzd4ZbpXBpo
Sur0bDrT/sZrwtVR4b6Wx4W730XuYDFcBe+U2N7alW2RVhToty8ssTkYafAd3/QG
SuBMLNUFgUQ035MPrM2vuTTMGWj2g59/DqfWR2TEurqC6e/eDHcbzuElTygTsFij
qVXYEA4NXB0QkPchr6neBlF1HzRrKzy7yFUNWDn+GkmpOv7erEY+yR6/NRXtu8PX
QGNaGadD1d5UJtmFFu7xB8jGKEliL0LdM10AdLXlXiMGI9x/bu/TrQajNIVNhq9Q
hhOlvPJf/iv+D/Nph8zAHf8cwJoU9/hAfKT4aJJAvUKEgMdswr2Y8CMP3LxwkFu3
0gVYnYyatSkwdiMb6cY2Z/wsolXhwkABAlq6+O8Tau2gU+DeSV6Gtu4sOIzs8iI9
HWLa561Sx3AUJU6Qg5k82U7twd+OlZcGZmMeXkuiITxDPCFukFU0r5jW9waXzWLp
Z4GaR1+sQFt3P+TIGYUzXzIkY8B7vJgF5H3E7qNlp8yJGARUWaSIkFpEEJqcLusl
TXuAdamZp1OSHxNj0Yx6iAbb+zCvSGltrUNKPmk6hShrCceTc84JoQMoLrw2Temu
yuP5Jbp7oLRGNL62SPXlYTCRsXvQRnDiHTDJ5pu/yvMei9OxgpmZs0+kNHIIIuAQ
P8V7FjEy4VlBZF4oQGDRYzOqSnfw7ta57q/LkTpmOMheiR+oYGP2xJgFn4ryjVC+
GQ6CaWg0tM1XEkrui8RDCHyY6KAser1M3n4cy/sY1EL+kZJsFJTlsoa3/F3mSuyW
tiqudJh3nRc0yeJgj/yB5cJZqW/+XishefykYfl4Jzyh5d5zjl4Wg+yrMYyNgYmW
cnXJkcYy5LqRgI0o7XcWrTVTtmRG54ytCptgd12iocJ6hiuMSeCkeQ4Hm5lnlq2U
48E3alAf+6/OEZDao4KP06+KEaugKLuENZJUD1Aq5wrjTLZiGPRt710F2y+2EniN
g8pwRyGqT0O++vxEsCYuebCQAoYGPCy/AN7Y4CchYHqkj5al52mH2IIB52PM6luK
YVUxd3tMD53V+KOGLFCZauRuPhkzmKAcOfoOmWN9pFhsu9v/oxFb/CybJTyLm5v+
K330HNMDKDSwZ4ZrT+BGA0FWgxhkDx8tRvJBJxwEqBz+iLHvUj58fd8uHGBmZVF7
3pdUaXCmXFhjGpHOBivEt2iO1F3MxWTFoJMH1K/Rcy5ZeB8n/YiSxTt2J9tcRCvb
hXDuUEZOeOi7HqeWpNY/q3TJznDlCVXmOqO+FzsJ8Ei8g1Otk0yLaQMOf24cNAH8
ZwGj8TVKOE3kX+9XIex/vv0NWhtH+uPx+8SyLPjYFpwEjHtyHVRmbnNxBT1L/tD/
oKUUGItCkj7zUobVgK6kUU6D/WWmdh5nOehn2BDdzMQb2hgkLF21N83OdFaM5eqq
4hBa2P9k96vLvAhK3/8uHsJr3UNN//dntFBLQucKUpWb//RrsyhbS9itCc9LqE5D
+GM1RAwHs/xuL/qNPPYng8wog3XYdnJKdwjZvAjTH11LFv63p5Ck3p3rHHI5lrga
05iOrn7iAeH/eDjqFhc1Dx5waqr0FNGQWa/QERTYbwb94L6L9HtVGggAtFUJo9oq
Jelj+RLR3BUtHlErmuyjFGHDQNocZT4AismS55WFRJ98RLck4DMq9XmNtX4y8pjN
Gx4kGpWchT8KjHl8JM9pb3hD6LzlzCAKgF/cPkcqynyNi/V481hO9F6rWBtkVQnG
4RNgWybhL+qTegh2ugDlk47K7R0+/F4fgOdiK1I5nnwBQyB7EsmMw+eASsI0wExA
xDYaaKuBGmKjtH04IMFzso46xrjP1n5e3JMLDHs06FQCzttbI8qZHu6H+uKTApDS
Cn4Wl8Rk/LyYnLsOFvLRngJ6nIUKwQIQo4mEYQraDj5rtnKf1iZ9c0XEqKtTOln9
MGmwgldAzc6B5DKyIMYnZLRWmUV2QEgnS8pOSxVgJs9DZtskL6uXqK4v5lBq51e8
vtyU2nOzRG2u2+ejZMrvjxHW3YZL8GZ5FWzGAPQybIBiWOlahF6RVAkdxrpbPSQN
H3smVGe1mw8YGPnPVEhd5yc/HkoCUe3RV6zMybA5cNwZBgAkdEMb8JFLA9Q54rNY
CLVF55c803gadpqr2fwUHJbi9lqrxLC0lExN6z9XllDYRJM4JBd0KCxmUkLVFRXb
Q76qRikuOyd2I8X7+DUmwl/Nd9+VKHHkgoLeheW49NHQ1SrAC9szA9bmzK79wuW/
optmZXRA5MeFukxxtNDC1iQUfEt4LPZd4V48CJMeWXBckSJ3+0WvrfC0KtLFSr3r
9DZsSJZVW8pAprlJ2tqaCcomi90Ou4xVxFIlKXOEyf3rhsrlIKbT/V0DcKc2ZCYU
9XRbvNq6ToA5XtNfzRSDoLWIo748mXhTmcmwMY3uckS8aWWlN9jQEfZxrapYuDex
Scjg+pxOS2PUsNdMSXnje4V97dVrRGPy6LPTaqp4ti8fOu20duGO+ZkSQavkT96I
fsfPQhjT49UIfaF0TiJbWL2l+7eNXpQlEZrr/cXf54STvjljxyrMyvas8g1rylOs
8dpEwt7xxEFsgGx9FxWdUq+g9kdjzS+bD5f0A6S0l+hTaMHRCwEZfPdo7J6R893r
OfiTGauYh0fNvSMXVjgeqp0lapMKcS1Ec+mL5mQY+XoAPzWtoLmGhYkRhA+qt7Fh
2kRu06wxs+iCSZsCi5gjw8kpVJuuyT9rYuxJWefYwKRzjUEBILKLJMEPQuLDrpUm
furIJZZYAu04CU99WHM8SLmFAMBFqCPJxk3rjGcpnF9FFBYmWxIcmNWaaTNeLZtM
3k/2cjLP9JdwtCHoV+lprtuW/689SlSWC8pbg6sqvkAV58EP44P7/aLAtyfSpLMR
O8RtxzMJCO1HcY1qXLHPGy8WqDM3hq6oo1FwGTZxSE5c1Yqo83jrojOqqynbgP1o
nHxcs/qBCe9AjCdVwJnLCCISHmG1CtrYsOnD8i9JsVCAIXSKfqlKB9eCLbxVeXWn
XO2B3kJsRsuo5h+9uxwag0ptocESFajrA8q4KUw7g0VWhVoFbMdOJtU0Kk3ymKZ9
m66PT/i+b8Bca9+SznUpcuYp9fCB20Dj0rsY0Dkqoh+JrUWkVBD4QaxfBT655I/u
60ts5LuRmZk7/Xdguxdl4APsYKjYi4v3EmMMA+YesidiLqayUfRa65v7MCf1/g5i
3D3AgZKL4QY9XsdNwSE1hkSkD55WBBQb08563Swckwp2VbdMTdzsUnXLtPZLNage
/xARx4csUiWtG40UnPa/kq/z49kKWECm73m1sgEalwmKve0dUcx5+vBz28bTeZS5
C/wyGm++1Hc4RA9edHAdNz/FBz6ckzKPAde+IC2lUE0Yb5YSJjfPTnZgCTBR+a+8
j6+VAvB2EksYuFWUmir28CxIaivKL5CSid3PjlhdeJu0pWrQaR52LhAOOn6rBeDF
2Iu/DfZ4I3Kgg68tDpZq6+UJKxe26FB/1oEwdDpAkfR9yqjcMm5YGAIfMS5ShFX1
h+UFijRMr32T0RF1jQkGvgtXeStCQL16i2Di6NAgI10E0cfwtmXnNdLGSjGcnzHJ
51nJPw8ZGmj13Vejx6SJMmd/KMTOaldekb/kOnIBK9ob494y9R4iU64SFXOGfAHF
bDjN2NhxPlfqEWTOKjGTUj1WC2nVH6q1HdU/+jxx28yv5YQqosFqSyUNSZjpXEUl
IcWenZjdkOFgtn5EilJOruUkCy19Toiknl96xGUH+jEITrHCvt9uf2ZcKZkecJaZ
rSEpzQjw0z0mWpBTZH2amHYdOVrWF3sGl5LCu0YUw8rEApZ0yU5q+D+qgLJ/EGPR
k2bjaZn6zlPqGqR2Ib4OVOUPwmUAnHOeFC70ob30w7SuozyiT1Z+swfCYszD3kFD
HY0u0ukTCrY6fDl0rZgQhFbMAqelojrITo4O1aRp2hYtKJaNXCmUmH5bsLLeZTC7
mI1ZxxSb189LKax/IvtuRvFYG5F2wdSOpaDs99QX2hOSGgaTztitEI2HkaAzwmJw
D+T6ONbovEm8NBJVcPKaZWHfhO3SK1kTN3RCE/BscBJHNegxYozBMS07liWpekuK
gxT9nj4u6nWjiUZDV7EuVM4G5iKYmLs5aux88BIZUMux0c2ZPPbLQFxr5LLHODID
F9JbVJvZyn/nFynZ+zbchBcpubnxzHff5BaxQaQefPH6Yu5Y7TtoEQhP/JZ5WXjW
U0pHYmN0nqttto7kowc5PWF8Eezt7Q9IGQaVzCYNG5P9J2ubOh2VuqQl8HOVrw5A
66ZrBmXT1qxdF1Wc1D/ltTg67fDXh5EBm6nai6zZ+X3+41uoNL/2Hk/C5xCjB23m
XIXEDAogeXrzQ5jidQ16hPSz3hGCyREwJZhXIDa1fesPozpfw0pxeQgpEu/Tg3gy
RohWkOuEECG6srRgRar0E3Cf7wFvN7RITVyJ2xapHGznfeiDIS7H3op9wE2cr/ym
XAhVTUhbElCs+MZRKvr1VfhYd16//Tt27swIB1mnxo5laTEGe/SGL4h3XrSWfeT0
RSIZsHkG5INNio8mrnTRQNExJjx3tpPjW+c9c/C2sEJ5t5Uv8KmcDMjCk5RfKr6D
JvGpRa62LZ8FkTds1ifugfTOACOZSWsgN1CsxcwDHwGQc+cFHDSAvYsG61OlkQGp
jrrJF/jnr0GFZK8GDaDiIm81zvRHvTAkNPzFtSz3aAG9Codmf61drEI422le3MaR
zyxY5sMs+n6munE+vhM+xNdf6RIxxhZ6FIt+wNLOMLNiPhM6YtObgF/Ix9bSlLAU
hpMrEE8kN8YeSlBnCoGsjPws4kru83J9iVD2gSBz8+FG/ANOpMRpYlmsqSdwmwek
L9E+nKwKHBAK8wL0NlcBsqX46lC85EB0jZ6rrGj+DFUscr+4ozUy9z8AzkSi1M8V
J2jzXGJvM3LM7syB19mWWHSk6YaGSPazVZ+LYhLOCMD5ON6aKuDpOtvdQnrsXMEs
2vmWSq5iQ1FanItmiebmW63djOm9QSwZHH8odeQHVilrbxN57S+yGogGHGj0gs67
sxbnxozhnKCLdavqhDoLsWmhXpT814WmmoSPcyGradHWpzEh7mXfBN6YfflIW8j0
oFqlQ4+1wgeXg3gvuai8TNivgGuVqiS5Gci32z33yOwY17FopIXnO1McblfGSzGC
gV3ICdelj9LAinWdPQrAUGSHmbs2tiG6M5dL60/wvG8vSIXoEvhUQsR1o61iW6Ne
ruZa5DaySRLHqJfKiXAYfDt4GK/4yOYgxUZl7fy+t2ST9vjQSGgLhW7uZqHri4hk
BD1lP0ewa0WmkuyLsWDeUNsgi89PvlFCHcK+xC+ZPMP0nnBdXv6gvn9f2bL1BLXA
IvVsE7b5X+dng4G7zACkt4urmS8E0nZbcMB9cQNf0U9UxNIocX8qbjmMqz8jodOT
kHOMJf8ml0KLdS2k4e7wdvOu0+F6vEwnzphK9gNPHcFYgA3OkhJJfpTwwevl7HpV
6EDDU2mRHn9Ae+bAB/ZaUWLqFD/NUuSWBSpz6GW9TCnF4jqJ33yIxhxgF6fGasFa
ZinmhifGdm9/WFivRHW8M3NsIM97gyUmW2cfB6Khr53BjbTMk4voc/+mngO92pxH
7we9bDzqRpr8NUwvIh5O7EZ5jP1TtXdw/5A9AsFR5Wf09Cn7eYc7fHSFfabGelnY
KpvDOKAcIIUzd5mH9s3ubdRZrhlBkxcoP7vJQ8BZD2vaC/IlOmzMHsR1rucZfUsX
EiRWU/vIHkQfnFN5WRDezxSz64wthEXsnGKwbyXY4G25O7D7tvkzfEANhWCD1LDn
yDEjBU0LKwZEwE5+48QyN8z32MHARQa95VskzVIpXKdWGdqiTOaTM7cfJabb2GVL
7LWKQ7hreMcUj8i2/t/4YUFSjBmVnU15+mle3s/X1SZoUSn+IJ1RiIq4kgTALl1B
MMdBDgRP8KNzDkB7lQAo02SGfalQUrQiyVn2aW4UC6OPWapNzec/gguKAGSTa5q9
7syFOQr6DykT4wzitPsatMncIBoMAInbgOjhL6YxZMkSOJfB0eLvULRIliIeqT58
WZ+ZQYSpCJgi/KMNbyOpyLilTEfu05YL68PCM6cDAARxyUbJhGg213Y9OY3lOITA
v+h0D8qZCD3buBccvdjAokpTRh5RHHzvxzh23fzPau5X/vonlN+7+sTL6ETCFOnI
3G73KwTq7z+RTFcebg/gZoAW+gT/t8VHIBqbOnP0Cilx5fXL/7K0/k5YVz1O3AaH
+td24kuqJilWRVOzACLLXcnTGbCxeic2By++jMXXrk3M/D26N2sepQUlCZ7QjI8B
N8fa17hwWGPMs0sL1NMcSu0WQd6G7r6msw4P6Ygvga7xTHnGCqXdxhstaXm2oMe7
24Dg1ObMFGCWo6DfLpf+5TJvYlbnwASaVzDiBg+cOJ+zlOpXMzgFMJYNNCDVFD/y
AHapAj8tLdjpd4C6bihcWgim7MUGJZc5bH7OCLS9ZB5RRRihh8x2lp2nljRt3wMW
SaFqvCtm0RhQNNa/mxK695VYH/E8+TqmelPRaP9tv3oF3XjhXQ6agvwrtZ1GkQMo
emu2G656EIjG3IIwsOFGXcSMXx1srwE8A6kWzmC5LUBr0WZy+OXX481Mqpf5eLDC
mgZDhPFO6jy4Tkfd67wGzQ6bj0wSlnaIf2zH6RsNotwNWY78abDr+YhxNuMp2ebF
zlUkb1MR1LoIWjVKEG3VH3OBflcUcjbVhDi2szNw65mPAb0GW2SYe0cM7bUD+Iul
O14aBOKMj7cUxJ9c/jURSMyWIhh0Ptnstf5vTzNxKAepvdlVxi4lxx6MrvoM4CCb
oaX3outuSZl4YX1sDdx+u1ieybpGrq5XN+zVpq6r/jviA+j8WG8TXRrehyLXryoF
z0cBeBy2CBnqS4gMCO+FnZSexZLSoTRcUCKB/ibFkA8tO86hQIyfeeOt0dkrr9kd
GTdTRqV5ayP5nIG0JIQs34PrursL27ByG6mfp1kWifRoerddjAU7zdn3yJiKts6S
DxrKs0qwZR48IUg1+ZfrOLr/LEWQ63R/BThBfOaXdEsZzYX53KaVCPyfAaoG5+wa
YrpydRmY+S4fWuvqEwpP1ZnRAG3pAc9IvnM747yhszF9dj+PHvs2cJiYJHoMB/5K
3HBlWFQL4iYrd2TzOU0IMWSeeilD0P/GrYHXcpl/OscRCEotI2P6shk3W5k17+tW
iCwhZW9xD1hQB3OISaXP1sfJ8F1cYn8F0CyTnYStrtp2i53f5mSEX7haOQM8B8T7
9BI1o+D+mllufejj7kpw+1YUbcNeOBBYbYr5XnvuNkdxCMWebABXR5aHX4oG8Lbr
QNOKBl7ILUlORp4IFWeChiMPP61fuHg0Cp9dNxNQtXu2YUWs1uwjPD47dqjI9C2t
9NczRELoNaVFMtIAVJPgYFtXW7OVhlseqHdmQKS4hRCGchxkAkh1XTN1XaLUbFAQ
KRbNjAS2wE0w3k0kE8I4irTVBOpmeLJjmDKfaZDCrdAs/Q6+hMey2I/uahuSNc7s
HAp5g89bG0DgeEji2HGeTD+J5V8GGEDOz6+iazVUKYo7VCzIsuk1IVXiDvVdy/mx
GrdRJqpLGY327b070roP8fg8qMruYkZ3e8vdWoGdV/3wegLAOCXNkySgiEoSsvSJ
XcGSAQ+qzl2rxZu4JbACFnN++5tCUOYt+oMUKJR0beTrsI+XZ48ZhaFB+MfQWiea
tMjowt0XlmAgajm0ed+X8vBagBGu57s+FgmmhIm6veXCekKfdA9qH6zMYGoV97O9
4rxkTfbuT5xLZVDt7lfcQ7tkjPgRqI3IKXhTmHnCo5mqMPA/6VYa1f/ypreH1opH
EIhPiSI6WXfHnkQryMFXoT+lL4hqFtQqqxA7X2JE4YuieOC2SLDkCFWRZ0DtESSj
0T2Gppb6eQPriQBcOOZ+f7sn70zWY2U2v28gLot5NFQ+dZ+pWhKojJhcyiTkwCt+
7lfhMlmrA3P9VUglOb2nMfSuyqNv8W2VWrAJUShf55i7gC93AtR4ZL7JjO72Z4/G
yXpxutXq5c6Yla0IGxQ+O0k0tGKU9uvB6NatLExXfQv1mBli1QT0kxkH2HBOVhSG
kG7kKBBsoHsqFHJyL9qSeWYyF7tCO1+qd+CM8MJOcDRwatYsORH4YIFJVgMOcrQi
KGGn9TIUkSdCfoFTnTtVXcnJ1BYb4b44K3yvN66lqWL0YlHycRjNgPxmy2lHy4TV
1dQC34KW63QgA98o6o7YoAKh9qM+MtAbXoxBgH36x/4O+BsW1GpxUOgWGtCD1yIF
3PWNYV2TEJNVrmb70lIQbqwmXn/Q45P9HCK1CMcxmUoT+Mq6njeYQm1+mIrsGdQ9
UjwOX8idjG0RY1ZwbqRQ7Jk6BTnW6Y9s71ZazmTcZyw13Y+mNsw3WgoJP6qE5DTF
Uy4dKMEnW/nQFgLUydpmJKCsxL+dwBfJTba0lp35p1yU/oxIJv1KjCr/Xhh8/HuS
l7k2ua/q5L/38DVE002Bye9iyijn6p5jTqDpdfW/uRl9zq4XtgfyMmc376Y8goIN
DdmzCIZeGYFlrBzaQYhDz8NxaGX+OOUUpu//zR3SkQrgKVtPZSD/LElTosSG1oXS
gTura/+x5aq6nwd3dM7vzPx3AP1ei3yQlUlS1Vig1xepkWOMfZEeg34sKFcsrxDC
aZa7ByQYBmmgiCvNe72MiW8EUvPKo/hJtlOpOZMOo8pLoO6BM55UQ9VBB7A4Ws3i
epBVzGBMr+veRRgCIN44RR75K7R8BGO1Q6uu4veZFBbsdtfh7CtP0NNDVtzCMrXA
sQVfTYbkQmPipvqNxKkIVOnZb9tdaCrSjAa+y2C3zTb9nk+J3IOaZJ4qu4YJi4ak
MmkZOzImeSor1ph+HnRyzDmB6uzIpYMkU336OtVzh6F1nOQfB/LKkIiQ6lQZocCK
EhZKIMLrVl0mlN/1jKpZpazGcO+dfV7CxSLlmD0VBz5FbaaqW4vBAvyHwPOR1ZKG
8x4MKDwWml1lVCCYH6GTaPjrY9wB0rrM1AngU0PFLHGmYcW/Mk5EKwK4VABHGbvd
fdL9MpCpQ+tIrH945x66PnvPmeBbsygZg9emHkTr4i5DRdJoOXVSeSaEWtFyYtYq
jj0pCmYRSVlUQ51RCBvpUd2/qL/7NlNG0CDRxdaSK9PsbSJ6Wm3/iFj0VYeRh+0h
SFOEdpKeAf2/YZkqjGVUilLSZe9anFMoIr16xNNmCu8LS1/5jQDRZi0vFVgtWGc5
lkf7xSD8QU8/ngBXReDa7flqfx0aC//aUEyLzL8RuhxpO54IxW+RhtMs1CDj3UKa
gr9zrrJqUmcSYsT/kmWHj9pgur8Ct2+OCuCEI3Ud4TVnqqi0SQuPU5AI7ln7KT9A
hiT4KSpLvgpJR8JzQ9m8fT484AnyCVS/di9EO2hX9cysQdcVA//0+GnYXjzMpjdg
3KHpVAjJhdutmRFfo1xbZ/H9E+6YJNXh0z41IAsnI2CZkcNE6bzKQD2Y0hRB3l1c
m6wF3+I3+9+zvuYhXk49ETNerJZivRgBEc0mYg7DEQvFWQxyHoBSeUIIGljo7W6+
oAiP873CkiWlDeVrGGFv7+4K7BGHP0vtgUC2j4ABzpjciKXc8P/C9H8ZAGwfN2xm
HjTCwMcOb6grMfU5F0aGu4S08FTdtSkL7C7VAUDoGkoWkDScib0UQsNFEYxmZhvU
ztMZ+L4IxXmeZBbOAOnW8ELC+TGKxSO8bs0lmIT059bWG5tEXsgeFi/ugroH2MtA
rS8ZlL+kdJEms0upkQVPtTBOjbhzOwswC1CdBvZIl06ZCqybXNt8XgcQKa7FMnKg
GdZP8EMmeZ3QSnOz6dfTPmIbSmjYSbPuncTKadF0Ptsxt0bsTsTyAcux/f5G3+OP
eRy6TQd/lFBtA1xjQw+AMykLrH5PTbKhRVRGIx7C+JzQFDcOu9nwKP33nwiAwPz7
gndedWS9FQtnLULceRGKtI9NsUa07JfXe+Rtau32ILfwLbUfbmSCYhUo/LuG+hGx
5vrjDgIEDYihzSksmni9hpM7j+y5X1Tf7M1YddFGcGhHsIESJ3+3ts5ZXQfIVBBu
dNeKF6Al+uCH+cDXTxoqO3BHB0qAt1UQ3EHvuqG+mDJelhpIDRZrNgOrJmczIbqB
NhqVQZIC8GD7AeB2fKb6yGSDk62hBmum+KDXbTFo7b1yEHa/cIlziPSoN7nt818d
uQ//rgX3jSq/SNPVhCjT1pZzANy0ThNhxDuAdaOWvy92FlNtzbPjcmv8TKkbZeq9
zAkXXpdfi/Tc73tYqh4KVyYPSGSyN7bzCOr5LVBzD+Ij0UpQNIOvZXBpRE0wBrjO
KOAFmgioNtG4JoEn33bIR0+jt+veZrbTM4AWt8UZw+iUWi0x/eF5fqaY+oKprDwH
K8mYqoukBOAAv+BK+lozsFkHrGtQKXDSj97vk8RAaXWrs83NS6RP+/2FlziNu8ZX
X8P7VzPeQwCZ/9V/30sHltfRCc0h0fo6I86sxMGS19W8i6sFrjY/6SHiMfTICRwi
BgjwR7MzV42bPsyl9FSHBh9C8xFAkusymtzY+64QoHOFVmGdWERvOq+6eBPcXzw1
qKRCHvoN9Q/mGD3WWlRMWhY9ytfzhRryx+QXwuBL/4A9h/qhIa7xPgRD2k+/mdQ7
hAmexUpAlMG2Wa8RI+3Jek3zLa2US14qJTgpDdBdeWRiGG8snpR3AmB5pC7JsJBC
onUVjsHg7tCFshG1M7jk2CFDvknjSe7gRS2qZgp5fpqJphckdJfnvk7ZkUQ+Y67+
1G+7dsu51QnekFDxaMhIK8oUlxLJ7GCk+yazEdTN9Dnf7h7r2jjUUEaLzslRgMfV
Dg48tPTrZakDJ0vGhhgMP33Dbe51y4jgpFo/HvJG50PpgDJkii2/FpOIa3qTmJpw
dy9VIDyjqbigz3NvZOW2Fkau9x/OMpMORruPX+oB004ekGUFqD/N8BnjIm+oB66u
cLwqmCPoqiopJyeaecHu+Sb5mLeAlZ/jkFq8HcP5LLPylfjjJbdIDLFshZ8/vHbo
rdqWV8AS529o2OcKgrARw+7fnSgFpTU8QKVEABzlIL89QyrAthY3N2G+3srGM0E3
unVYpPzfPUkmovoaWINn+axwEDRHrc8wRUqeQSiioWHNTDzNFVLL9lAnjrFaXO/o
Nb4K1Xn5F+sjEeYGArK0dfMsv6tLWRigUTkwOXVxjOAtCcu5KMJAnUZupUAxVuLt
l+hiUEIX7CSNMhp8aC/8FPs0N1A6CdCT6GIJsk5ixJLcV+A8R4H3VqCrXAgYUFQg
ZyJaQmczNKkQehklmk8hxuE6alQiN5J+yQjLQwH4WtD6t7xOzZjJZ1lpEZpTgHzw
ng90/Y/5f9JniFQwtBmwDlosaNenlezFfO9aXEOjOGp8JHphP0YF3soajgIbNSp7
reii89+NUMRM3LDt1WBtFQhjqwCLDsxcyaLCWCWd9DuCZ+XWog0wnXvNqO1S9thi
fpam6xNlAzgNjtr+1QNUBj9Wm0GUSMtS7TFm5nARvB8f1vEPuM/bkeJYMrDz9TBc
L7EgsV/40WL8ilNMTwbNObBgy+pjZ4TSZ5CXFa5z158q8SlRqLmXo3b0sYncecho
0dMAKEtC+K7NRFfY33Guisym9Ye44K1KnfzNyeLxm7Xhf9VEIGd2NgwXMUcqTG4R
PZDB7lpG8J+2zg0iRY2iHdzBdzL0v1RaSUsWISbRVZsnxSMnosAVXAkzH8qDetoD
3lLQC9eYUu5MlEAziNT8Dk8NHmYfrfPBT0XFtBcKdh9TrRsG/KEzL2b4uaUkHmqK
UMtXNddurtsV9CPq3X5gddfTDsJ6WjmX3UHw4/CteP60d5olTJ/fE4NkmXQp+sF6
bReV/dA5p09E4GSKdJ76/asv8/r5AvgPMhG0/rQZbqF4qP8FqI3IeWfKRs5pSTT4
ky12mkBJhip7uV5obrnpS8uPVWMSbQnDsorn03xHy32/eB/caH8+s7FQ9JCFuu6V
7xZt675QY8YJDgmgAuFhtXqUCrQzGG8YerOzCBYouIPX7422snFYqKb2hZQ1AMJH
ElXEiulVlpuzfpB+OPAqcWq/nfozr1GBIOh4GV7czmilaZxFJ0meCx+CwhdRh8I+
/fb/B5t2KNiTAAZ7Dn5rPOGTfeyqzmz930sHoYTPYZiH++cNzy/gIdFBhHjuLvMP
wDIlux/mzCQS/YMn54fR1oAV/uRqX/kBZNofYb1GHQpAU9Sh7I85SqGh8yTf9V7M
D5elsmyqrUbl5QcLQxNvm7W2HQKASgYkAKdo/94Tl7Y6qNXE6zhkzzXIXeZQjPib
KgDtsvc1pTYnNrn5NBUcoQ0v/x7HZzBGNmuIJCKwaS29Y2VTktuXX9wXsSMH9lLH
SkvGhDhhPl0FGOgpuK8wkMvICEYR9TSFz9ZPqDaojmexClA0l4ujruW+/PyCnlHg
CgPabE1AZyayFNaA5hskZlcWAcEuMQbysICcOcTYTipsvVNyaW4lz7q7t8tRDs9w
cq7Ls2ea0sGqDV0XMr9z6gr++bVPVhXiamIIIP9xgTSj+F9+rZMVU4p2NxoAafJV
Y5zutfCqfqE1WmknNq0or+tnCTdwKKe/ofi13dSBaeetzWIUmy7H1L/E2y1sEQ81
HoAyeJSHmIRtsUfA1J7Ci3AlTsZVGacEkoc5CmvsMefvxHcjOs1S6yH14lxbiDVw
j9u6jZDlaKxsDKWub2nBap92/rB0Np/XQ+ShfaSCL3ogFzrBS8GcgNzw9V5NH8kH
5FC82a6s1pZH+9+Fb6APWJwRFn2XpNBBOgnYJKQOd/rdbwBYN5r+9gpb6ey8Jwg1
YkJU/DyUOhcQsbFRPXofKobZ1odI0cn9M1C/lrVjt8sU206bsqoocQKiNWH1VaL4
0UvjLq9+KPB/15kJ3U5cmDWX4+y+BYDDYJLOfIBneDxqTCb9XhPcany0f5/E702E
6wb59FeRvo60GQrpdy0qZsliKRwGH2+Tht7difZCOaChy4M1u2R4JePIC/IBJupV
/D2nqlAEtfXMs/PpFo//UhQLlKJjR6r8wmlg5nkcR1jIX9lTbKDQC/09v1+vw4AA
veQImbSkYP0XH7Lm6U7BYRH1o97I/Mhsy/DnfqJblp1s118XgSld5Gjj55ib+p6/
6b+F4zdvTiYUeKuBWwxnCD/lyu4T8SNW1Oh5RNeh/ruJsGu0rmMvmYPCUTfo77Ml
dFuU7Y0azXBY3Wul9Cdz0xA8/77DBFnXcUtw62w2vjtLgCPEpQZM4vJTncsOo5H4
p9kEI0XUuOcD3zBrwyCdBEj24CHMlDjc5nqeX1FWSVJ4LWSotRn9yk4iAGgyXbVG
B7mMaFQl+ckO8imlm4Kz6rpXKiT7V62JaIBedFu+ib7lYyijSjBzKHVVgV8BRSuG
oE+Fu12qT0FqIOs0mBOOz8ghvO8r2Z4NAZFQkck8QOFlvRRjlhOkYGUfhwph4UW0
xCr86oezhnbN7R3pHzAjwagD1T3HtQhgy5KIfGvXRBHDYBvoxoCW3AZng8yl5vjO
kWsh0Ou0qFvqfKoM16F6sBhYi3S6Z7zB+oeWfIs9yAgzDbLUuek9s3qMxnD24KIF
ZDG1VJbJ7D2TfdCvsLWhIjJO2wvApgIq4TJ8ZZfRV9RVUg16WJYG3dv103z+Ed51
VHHqQKF/ngP2adLtRUq9J0YwXmCt3rzuS4ft8iX0938F1Bq1/qkRKn3F/1vGuB/I
wqXROiADEJpJRJ1srZfxMo02Ro5TeCInl3gUkxW+rPSU2BmxXnVhGKohbc9q6Xmd
ZksByN20z0CoSt9VaGC+i05IeRzrOGw58d26FR6KLFY+28ZsVa5giZCiUci7ciBq
MM6Enmq72NLAYH7rHRQ8yrDJN5xqqk6sf1sFaWy80zpx62E0o5cOqO/JgEWf8XyW
xDxxAWzBC/5eOF94rR2rX6+i+DPhjonrVDYdm0VTo7gh6UA92mC6OTZmf4rNaBNC
nHuSYor+tILunsXyMF5Ny6nXg7rGz3Kfvn3vEEYmp8+pPMbco+tmUQQ9DRCrg5ht
CKMHdSnRaKpG8mDJvSIhde2m9VyzdC6oiqojnqaKDRFY3EacysOvBpFxOY6hTjOF
6eRDjzpzYqJ5J8DXXOt6vRSOh0HK8KKUJ+i+RDVDzkUcRKDfqtGkv1t2M82Enb0Q
WR4a1d+GEY68snT1ZoIkGxbN9U9ZVhrm+hegPBWydVT8A7St2NZvjL8u4PveiUpA
kRettTDWmq0JGbpldigZpZevbCFacFg+AEYhfvzt4zpuMEKZ41Hfsvy4fVQ1p9KE
b67gveJpVi/C0h1h1SkPrmwqwML+WNII7BzXEkpY1GicTL+vrcBeivddunqq+XmB
4qYtINIkp/9s0M86PrPExSrW/iFzCBaRxmmd37wNuDMLapXdMR/fhnM+bIqUN5cw
l1SedlKP8WpBzp/3sOOnVsFDA/Zt/5Sw7wFc+kor9KsSLBr/aJ8FCSx665dLlIjo
OhQrlTnhj02hlGX5NQISbZU004etNH6pL8jG8F2NgQxAGzzeYkJk5FWcy3VmVyj6
0JjUpVbup1+WRL5hoq7FhISjzYmTaKVFBdHNb5wSaoNeYFCyo9eKv/jzar7SiHUL
xo+9VpLyRydKEQUYg/jQ9T84nxHXbwMHjArDQDt2Z7MbRaGRW0xDHGeeu+6MWHlz
aQqbzweNj26/lfbCkdLMhQYx9il13/rfu45B3Uw9FtYfbgPdg7RWCo7B1TqUEqUZ
DaHnATNQuJeC5DqJPl2vsp+tkooc3Ty3zpo17UhchyADoE/Xv8RXbjFwkVxUZO9R
/ssVSl9WMcdHr2X+l3ttyf2vyzmHI8KER/6hWrVmVN2EZvS2pI7eXkhWGOgZiisz
VYbVfOaMWoxga/WWJi8hMBAFeHiszjGnIhVvvgsy435K+u+YvjQ8gn5Or5tTiF/O
HjcG2Ww8zF+YBlNON/dNn73hFO2XNK+AsfAk481DoHyZPMfZLbgbO7UQ+DavKuVq
ng7Qdo0rkw/lLajRDiuCzw8DwxwumwmoVtMEk/dh5bZekiIW1M+DIjBgexOgrsho
AmiqmIX60qozrFEZP6TIjVTM2bQrNNOXfyCLR7c5TremY8gOao74GJ3ZUGmVTmOB
l49W/Ku0E9eWa8CuUrSbwLQo2n9lsQ0at6PUESjygjQvftfwCMP1ZUNLNFAJTms9
TTPbmIPs0f4iaupz4rReQoQGPpeWKkuS9qmrUtYNtcmQjP+PQm20y39D75R68vAT
SeUNLZsbfePSlF8poPOtQB+f+Njq4ezDwXTYlXUBkiwLcBsgwWSjl11e18+07Bi8
6HAvrDZSRE3VUewhp/qNs+wdJTVOjyzAnueYGfpe3gC/EZ3/x59CcOyp9JvoCuZy
PCObn6dwc9dg+w8fpZZhc3XrvCnsJI5Gu9y0ANmWFfiTOKyKWzHEoVHLAIShSexP
rXHbJ/VIjZllozIFIQWg7fx2UuJ1oUtoxvEaPSLdaBWDOTsETxYKbO/3Sk4xI6rI
ko8jAOLFeJDBeASFvz5MAMNiViIYq+3xkA4jD3K61adU9Lj+Q1/A1ku8I8kb9jnk
xg9Y9P4slcI0Zf986mwIaifGj8CYkMGfVwc/qLZ35b54L/raucG3zU19RFvKe+MT
PznSgLtkgtGZ7qpxTTZfG5IBUzNFlx1KDAnjEfpuxVsC21jfAmhq2ZNgAd9OLdBd
MhBNG8uBjKW/hkItq6QVLQAtbuB49il7qFYY5BAKVHI2bjpRBzuHSApNJ5264mgj
3O3SOZCUvqcE7GOuQ/3EHf/5i8mM7rw1hTZd2GkTs2o31+iUp5lnlk0UvtMJD4BA
kLwWh6SecPFNfT1ru66FBtA+r9CkonlOkpEKx2ubLUGEzr5G7Y2Tosrt5M72UzQ/
BufONZSE8NMLtD8BIt59l5PPNzoozHg1c6sa4+DQ3DrRrRvejdN9sG0joJLpxyJi
/1GbQSvSBh/gDrotWBhd+sPFY3f6iAlSwVSv2CA2VYsFkHjvZUlpeqFzbOo9Rrsq
RRa3eGCcqp+xLgKp/hrwTFKSVJWb8dgekylvK+v7MNn8G44BPoXB18W163V7MJ2+
XNy9dWTcPVm0g7kPtJQrYmMqvACQzMAOA6ZWmb9d2jcINZYQzG+fi1Jqw2LerxJo
HZjJtZJARjvWc9XaKUqLa25m20dZ9KJVl9shUrxacU0GINl0xOZCJwYfygp39KVD
XcOpyNRXYp+5nc7R3BhL6gM0M6QvErPU+PUIOtKuV1gu9wJVx0XqDEq3J67noHYu
uw0X3WM2+LV/bxebJRGYjTPOj4gGL9jdDgPdKvQX5WevQXgwMbO6OS1CHuxOxo0h
ZPKUkascCXbOv9KajZZRbD8+Iyj6wcOy5Cqh2Kt56uF8pjL+cs33kLPiicvDNZTS
6Kv+YPKPWykf59zrx3w6bkhYxM5azLiF5c9yf+BkjEVD1L9tnPC62LpStSKsenYC
fraRjIEaLZr/YMF0wCuj5ai9+842uuv0bok3lGAZOD3ld8q2mBrjY2aY34qjse1d
kQ5AHuUbnAFlSc+nzIF2zakVQxITkcG1tqUYvKFBl536GSQEOLZtZ0Asg0DkLBGQ
sLVxzTGlT1qPYCjHfbwBYKhXK7hTpzzKUBhUokn0SEBaaK8k/hiWpmK/dePbwPce
g+7qm3NzHQNS0ouOfI0qx+sYIddKNKO044JfTQVx4utocSphc6FKFPR/1lKIj1lc
PYpG/26IEqz/ShYQJ10YzK+yd1tVIQQzDB2wISln5bRUoliGWBUxO2Og9IKWj1v7
GiazBjOxkjznScdifaN789SmLlNlgxcKIpDpkMzPMaP70PiBY8di8immV4vKQIA6
vfPV0s1bom38gj1DsRA8wlnTCqQGQ21TG5v4WNnWjiwkQnF2pjKcYWFrJhHjVkR4
y06nI+Uokqsi76o02kSFnY63K1FlbLbh026E9aUDoJbkjBYyFqTjQh/SxaQhNvvZ
FCbUsUQLpfN+yXBJISXUNQgqIOmT0XvTf4bF8a2N0TTxDumsHgzIE8cGcDh3wfkK
W3CmITUrIU3K1G2XzaUMRsZkJHyY3T89+jVY/5rP3vzIaYj72PKql+l5ley7LwyV
Tazs4WJayTRAKQm3zOIRw7tHsbyYWSyBRTKOofNVk+XpgDa2fn3EA6HnBOvFl+6X
aY/sGrGjHItYTnVbialsOnZWdUw/FH6mbJvLR3hL8i9fgAuvmWfMyUUuTx0AhCjL
mJRIb6fGrfQiRPZX2cVuZDS47X7FfZ/RcwR35B+mnqLTYaNPNqG0oyDYUY0ivzVB
wP+byzbaF8OxEQI0J4xzjP9WpWU0mO1VHpK0r8J1nZD57lVfi3NehrjYlV1WqbyU
VjOxksJ7c4YnXiyT1dBcz9A72ybV4DMD1RWSCeXM0g6a9AX7Ixzb2TQVBGjE0baw
SWqZNi4WDuqFckeIKhdb4WDZT7SrB4dE1zCbKxySBDrz6ofCTK4Yk4UMxiAB2RR2
p21a6hjjhtntdGhzpU2jWDMbwnwQCHRmvky6NotvMTmaMD58zEGAiE1fQsO+OXxw
kaQK10PttSEB6Kk+Bc0bXWjEmk1mNDPYum4ygmINVE6sMCt+d6zNwokOGDFBGiC8
EJCvoycA4opUZsBHQIYBDaRehmd5OMm8/8IcL5sCQK3wFqK7Imq00ImJhYVuuHMR
hzWpmjh72+4eGN+yVhdKCXd9FCKWlS8wiTgFNCIJyR9Zg3c9gpl3Q84t2ktwYRcr
He+URFkWjscoLyqwK1jUwwOpon67OeMlGkg+k4IU19n3v7j7qaDriTLY6P2fj59F
3bZVBvGPxT9P7ZnKbyBAbDXINBG8XJolbwhCTn2vWaKwQ78FdrkXmVUHj3pIfZgL
r9EhBL3rEYEydw2ii3bOEPgf1HPdIMuIYDelsCD3v71z/eYxGn9x7CNE7MBNbbz7
soGyl2hpMU/2UXeMXAQon/gwWxptzX+/T/NYEhwdbaCi2lI4jSY7aZyc3ZpnGhiU
jffqx/G2Gga4Fgj47D020qjea5XPBIZQkk1F4MOPYm7vS/Gm328SopjI6GrEnGxh
l+tqnSHRJtH5OYubTM1/TSa9jQjd38SuMYttOjTcILx/jLEfZNgtbw0mF+ZfTpZ1
I9tYClfT29cerNkUlSbJ4SnpOfTQRYsQ24onNYrnRiQlzmIG8kCung+bmIn4xbAO
UI8SgA7NDDwmml9PNUfAYab7ImJkDYAJmBFc0IhAwtCasn+lteNyIQMbA6L43qJO
JAxduTLdh+9Lk5flCUys0JAqMKDFUj1nJVbWQ6nzwHbbP34cLk2e/vBaI3Gv/DU1
jFXADkFKRpGpwUQ58+iBGieRW1pQ9dJVB3bAL+XDR8oExRISZZjp0ivdABtH3UIi
x9r8Ho2WkKwNA2r2NierS8T6yYwJ1Rkiykd1zCuK1SymU4TRiZkQ7osHth1zFJMd
QRRnc5QPgnFqaEycaeCM1p2IOZ+a2o1hpzk/oMOvuc8mmpVRhhOxh8fYoqar83cq
CF+luaUEofGKcwSl9P28fq+O9fjEJ+xXP5GAIpHuqrGtHblr/zHRbcSkQ4pcyAJr
FkbKvdsR0pBhxI9euvZUuOjm8BoUjfXYdDd6vg7HB6iONUdDTtcTqEJLnZcPX4C2
g88e2jSzk9WCiiYpCzPm/5GDlWha+3oCDeHcJ/CRK/HcrByTNlRNXM1PJ6c2rKbl
oV9K8wIQrohl/T9rAMqBfvorIj4zaIXt+Yph1emPMGPQiwXIsln8s3oMv/PPhoNH
5u7LqnjN/f0yhhBmmDf6c1/9EM2g6ODInsOlEtwCWSZTAK1ML/bvK6q5Iu/wkBq1
xXnm1jMsLbTUrIAU7RmTD61bDdcZgD/KJgTKD00XQf9Jvr8Zu8h6JEIrJNSIK/9e
hoeTlejbbnYM0Ei5UmevmbkDMh4vd2Qx1/h0NwH0OjaeZvvN1Zz9laGSqkmNCrjw
ACjbAY+624eRdIm1ILa1+31Iv82ueXDJrQqqhwJvvTzLylJO4j9t9Wqub8N7wX2m
uXPz480vM7NYNrjbszYG5MUsPxJWmOpOU92UaCUTLtNISt8+mtuLIJpYm0q43lqn
mdJv+GlcRF9vRi7YCKahRG6gC5D6/KmlhNExQPCAYZChGH+0mQOZeWTCPOB6t1bw
QCw/APm4xsmBAf7YsQNpoXtNoGGM0i6uGXrrRdgqSGLPWWsoQtpnWi+JUGQipQN1
T29/pONFgYMn5CRo5OsKU75C/1sQewbCyiCLKlv/2NTKZb+oWlm+pwsbfBz81t3U
Dxz/4VzWMZHvsEAHSyE2uOBnMzxhRLTNBdNBXlNWbcFJXOT3mQqpw1ZkIqq9lu5x
DvqriqfTA8dYiNgti3ht5ml6nygZvEoJD8R8a90DjeTezYsEUFJqG9spOgEO2YU7
ug3aPy3K5kETmsJ3aQlpYiDKHbPhoP3o5IzewyG2H4qAs3cnlIJoipQBafT8UYmN
+dozrX3jQ19wTCn1fXSgwk9hKwn5tvd+FutgpWXInoWYsuwrd08dKAGfhTmRAmiW
VTcaA5GIiE3lNu2exzJYD3E7lZqgGXcDtEqX/hUP9D/5OK+aL3bEOLwoe0SbO9yq
7mgmF3l/g5o65rjq8UBuNKQq5RvGoHV+plo/gDE2RY6fP14wtRI9HNFVvDxMcwwy
3hu2MRqxW0DkDDPNVrIpTGqFp8LCKI3XzM+QDoP+WSLoynHml9iKsYmsWml4Tho0
JE1dvTWU436265aJK/5V6OK73+XSes+svD0Zvv72VbfQt6dyb6edsEbm01oObrZi
M9o//cCwGNHWvjn0ALv35EWRJpAfiJUU2ephDB8K0chqWRK6KasP01WegumJsxfR
Ia1u0Hqrs8xOjpjaRI7gkKbdNPcbW//5u9obp2bCLYl9CdAy3vcGhvjZSYBfpPAN
YEbX47NZx83e6lEQ+gqobXtqxL3O7V5lrM6OC2WQwiwvC6MGgsr8t9/mpECsy8ZZ
0cPwjZJrXmWe6v7i0Avu68jKvnI0fO76B18LIyUsbJUcOKinCdJ63LW4mYreR7Fe
VL93RV4P7uBWYtAW9itKSEx8jdrbCRkf/2/qvMatN5nU6d63YSG46UXJXjLyVntX
8M1x4irTSH41FwqHIezI5pow+ITSbyJe6dMuf39ZkwJoWKnHM+jkl11FZbenTR3K
ybB7L6Wf4lGqCJxALXOdo/U6MZ/M8ld3E0yAE9rA6ycWR4HzxyKiyWegfuDFk0gk
d4M5UJgkUV6YxE/vlPlQBOg0JityN9kpdXkO8BHCjqdaUAVw3793AHQNs3ohLJqy
e2k6/4DkFjinrxPq5IWTwle+xMHgPRCEktIiVhWLXI2PW4T1MRYIA2ZpcvnId9JW
MsTXX/I8D1Ih/KtuahV+Z7uPWoKIR3zbC8cNGXMLQzHwkNfNyIV3Cja29ToOe0pL
GvYqhWYuszjeMW75F+epOLmUBPX0wALB1hl6YGHZzxDcbE7obI4HAn+Oq6zKqI9n
cfZz4WUO6JP6BNuHadPv20h0Yz4bmBk1aUUvodHY8mtqKCzWszhsOPmqDJ74YVPf
kV/sVz6vhDuiwioopfoAL861BH0yTSfGlxkV+/Sl1nyrBI/oy/XzuTDtjxMsP9lO
tMEGkmimlHNLkb3NrDW2T+gSGidsqaEWwfAaVM+bqknxo0ZDYVnIIGZf6Jr9oUUK
VwW8RaU8W2Tw/qL1m/r8CXImn+/CJWQG9eJdKmZr3pj2l+qf3pkJXr5rG+pwUydP
vxwo19yKaLXqTWH5U0g87R+0D6tMi2FaDYMWC/oLMKLauVBOcM8mHpKNdgoWhWxB
Q+dxxwYW6JJvvXCxSIMYwOnLan9DefM5godfSuCUytIk5PASi92H+zs4NsMKL6py
SJRV/mqKTSCWcRRo2egdm3LyDuV2lze0eq724QRMySTEA44DN8BIHYir+1Gomcze
CyzdFxW580TcaqGJBXhiQGX5Kevjg4Jcs0jYxQveMsZaouyUHrHEJOawnt2xR6ir
efDrmZYEEvlrmhE8bIxTEBzwYS/3fVN/noFnHPWTJmpi1uFO5/j1D+BKOy3IObDH
2lRjQlo6T9Dfsd82Wpkt9rnCDNOPOrIqH4IcforOOELmdKu7LCPkutn3Rin5cNRH
2aVDbURV0AjbrXvOMT8ar5xtwVF6/nq9R9RgfcYDWOyefqfb3PMeWmMTMpYQ3tfZ
ZG2kU6S56TKHSGUtjnV1jE05BbTfbPlFzQvlr5v9GLpFU211+SVJagVtGAe88PjX
b7PyLaLL0fD2iIKivPorv98dF1neU5zHexWs+C96BEbIztM9mPbQAg+kOuTpgD6v
wNVxvfu0HwaXuyH+czmoEshsezM9OQ02JtMj4vMbGp5CDq5HD5DWdhcAL5G73POm
sz6nLIH5mgGYtD6sXcxZ/LE6OwA4kUR8qUmPvnzoLpgFnyRbq844eU2cJKVjBJvw
T7UP7zm1NS6KxOOdWiEXiKS/93HjYiXi8QUBHyy9f0JFs1sKNoywWwSoyywBE9Ep
sLp5/z9qacqjKadKZvzWGDTI9d3iTL1r8h32NPEyILl+amwmze1cvQjU2tgB5FFD
HiASVvQAj5jp256M4LNvh2z0Y7RY0qhnAZhQW1otwAar+s+2zlNVtkaDzbMN+Nn8
SuUFLgz0ggADWjT93UdiBsa5ZmYrloE/c9u8ZHR3OXA48xm+g63Y9YuzhPz+PB6g
dTJHk+rtemJo3uMBZBW7f92bNIm0tzIGcmBxUJgE6t8P4jdRJoI3vUtUy+PUEVbz
EDRihoyAQsitsAdpAZK0PmGutfM9jmua9d+jDgEOmI3PfYrNLt7a35p0CHwAObSt
DyQAl8r7rH5U/5LfQFmtJFzaSpNqO90XRnMu0XeTK30YXE66C82oRp+/oHJGdg6K
pjJ9I9XV3o6oIwtnildEDn8z30q6fEcV7TWPYNe9ukzpbqmcY9Ws6x1GBksE9bYx
2LRvNNj0em0eazSNETahIp73v0NpEv9O1ddHZVFUQveMZw7lzA/c5dzc5Qz8Kz5z
Bs8BpJU/vjemG2VDUzSKRZWnU8uKArw7oEpnXLdf+X0ug6ZJfTtd7gVfLGCU6ZPT
G91YKZRYrkXNpVqG4T5sPrbCUaRo+z4nEMerkwQM4OPO2crc+VPtTyHIj0e0cfG3
QVW2RsqBR6KlH1D1gOwkHtxgF03wC38Pfvyio+r78Np/daWib/F/WPHt83MpFBPp
+o6wWLZBD8qehoegPlZUi3oWq12UU3wv6QPRZ92xEEAJ+oYVtSpRyeivn1VrduUH
gp1G7mqostSKKV3QC8cyQ0OJx2QD//oytxWdiprv1pzZiVcpUtocq9WteFehc/AU
EA4v1c1o/5j+MZ5IXaUzLCaxyp/bZfNZE2TXXoNN5z2JzZJrXHFIqjd9i1ujp84b
fgaH6y9OIFlwuSA7QaiO0QEbl5LTGoqhPaVuAx6rvRoM1SkxQTu2GjPRqLxg8uLx
WHJqfLrngaMl+D0FGWtblsg7TAN2f7zI5tQzXtHIdhYNvCce3kljxuERlT/5sK8M
ogr0mA/rVFqUlNQSZrJkuBy8uFDpdpehnfCZEwK38qnC2UJ0gM4h0ySUNdr2L+cf
WGXbEj/j3cGrGeXFbzsAvbOYesclADeNtD7P03YzkF9Qzg0bCE3r9vYELj2V8iRI
w2FHsGm+EKzTBb0owN3Z0xOpsO5EZ1vtWxn/Y/BTUdV/RmC1t/jd20TpnEI55S+N
FOCrMGjheLM8jnjn275Q1drNNHUFgrh7cHtvI0Dslmtdokhfp8e3dOFQfnqXBzdc
9QnwfJey4xXTS9zjVYsl3tOEeaRc0/Y5tLy83/a91SkMuZZAqPiXuW2KT8y7l67d
Xv/pW5JhvQCS4qgPNfT4lM48YqBVsaclpa0VQu92IVtoAFc9VJ/if+0qEK0kdhXK
SpamuugtlOLZ1NqVoHls4p7j2teCj1B/z5qlx8yYQlWQ1iV/BMBf1z9nRm9BTJp4
clvdXoEZQPOmczqCXk+CMFdOEy8CSMa3ovwRNOVeXiaRlAdsGclWfGaqI21i0fwa
28KbVcNelNvTJYtmuEJRLMpYX3drMV4HwtQw8GZXLXMPG6R0aftT47+rEwAuGYp+
/0qvxPiuLG7ujzV3mVpwOxVAGf/2BURHfaielELDt1uvV3MvJvKQF7wMowUFFR/H
+UUJtJtRTE7o2cuZHA9Z+MC/MqiCJardbJCi+nYOLCTVFyaGCtv0N20JMXFP5P+d
m+7ysjFNsApm3f8pPHeW+GcyW0DXauGcGeXwmu7BBYrK0l0yabLIGBFRRt940KwS
2VunTabBElnUg4eI8p6CSJCb9j8lijhtI1P7Jm9KXPO+L+nVVgj4vopZzdArX74p
u4MDEzETnWNtakT5e2JT5BweTFRlhtrMRYnfY4zzGRlX7UdnbCPaACbrhnphYSaK
1UWeOm3kwQjJeBeOln+yrv8O4g9oKl5YE77hJvSmoeoOIBSwhu/m3OdzKtH7cVJX
hQIfqpakkTqSq7Lsyf1qMVyuc/fdnQWi9HtOQtLk16xSnzY0hSJA35Gt2DdyxK6t
1og6Wq4lxiwRUIYpQ+NLmUuqd1waaHHJWvibZ1nd6jnHWRyzaYAl76YXRsP51pUy
sQOEXI/HN3WHDKU4I3i5o5oKBNyjiXyBDGVedv0N6TpvqfiYvqqhlHs9oA6h39hB
lRBybWImBQR/vhe5zxtJXMWxKkngUNRW1zPIKiNiG+Jrv5yJTZwp23PDfolgY5uc
JNBkzXbbiTULOJhyPPMyTEusGfdK7r3rRlN+Dfo5nGcwygsnVj0RGEmi1gPgt3fJ
QgIyp/wO/VzsRkTHEbZXqAuf5tGY9YDMnD9P72zGmDrTfNSg7vF3J9OSIIdAShWJ
x5U96oLV7fUGHRi5q2UQqwgRVrt7lEpuUoy0VhpKb3yud96m1w2xRl6IHF6o1p5b
LK2h4UH1rqg0cK5yfhtNQHTfHsfXJGQZ1XT8iUt5XndC7uec9VhWmo4c8n8fpruD
bBBnlHe7GEx4dABm+pVfOjcq2tc1QrnJ2B7Uhz9TFtTLqOGfR9G/2zd8WxQInTm6
Gty4CCvGs7H+7Q7GMCoNQWn6UbQo0m3zuJZXaFc9PAwiv5Mz5GTngefaDOLHAC6X
rPR1kgR2b527wnXzfIFhXmZ0X473FPXWS6Bd6cWfBSqqdIp2OGkpyklamc43yQOL
2tyi4Jj8/SAj85+m02xFzMohTS8F1QU7aEkGgXBhhM3RhPG6TnjyzFKNteHYAVg1
Ho+ijw70jQ22UAoxKinP+3gVCoZK860oiDiZschRDCdOnknUz1+l73f8YmRIx6cy
LNRGfoa+uiK/WhBSZKTWFQIbU0g3e/KPxQ0EsaUI7rCUhxpOSW7lNV4G3D8w8AJq
FhDWXsZ0t9EcXOAI5jP9fYF15/i+nY4umOl26vmAXU6A0vXNMqevNdNgELjz3ryB
zFSkIGkNOmYFyHwysrcoDbrtAXE/6r4ZX5dOnkBZvkmUwpfjgcuRJy9c1P/jKPed
vphRb+DlfgrRuQDUTpE0OIKiyF5iFPPHsZwNHJxM2gYZ+pFEkimMQsatX5UbcFQ2
HMq8a7pqpkbfUi2btUJlDF7FaEdXYZIqiqS0rGcBDDYk3wEHEAqI315Jyil7tDs/
WTvyhvVkkBTXnX+7gfMhmnivDS6arYrTUbRnaAy5LtoOXKGQEjRznTPAAJLdN2dj
cw+p9QBgNI+45Bpdxr1hUMsPNR9Ie9Ck8VnnrYoKjn2ybSxKQMxvxTonDKz8Qy6X
6FbOL1paFxMbb7+ca0jBjBmDQKIQNFiBpgeKgC7jc4nR518FxbxJKJGsf1ZxongW
g/vWjzLnrLboxKRoVzULOsWk8tVn6zoAL1ihBTRT/gflLG4UvUTL/iB6azhAdwYT
ZlgdEWu/UvLGMG2fG9EV95ernylmms9cQZorSeQ6QeDOX6+kumX5TqxDQwWB73af
Fva7Q7dWPJScFNg5hUEA4KDgbgZ+AZiFoc8lheWviiye/PgjKuLJAei63X/ScDXk
TzgZmHuOgXbqsF+7Ih69BAY+2KG/CHkY1NIEVFP05E09yWL5CnRyOtqETFasv9Z2
JFF/RuEXrrblSbWGwww3UsEN8/DsVjEDyNG594MbniLAYcjwPk7pg4iLpgCUMood
qqmaZLrz8zg5t8h2wAk/mEH/A+KsSVdyI7X8BaxapNWsgBYa/at+BiPb4TKPT0ni
hQsNhPcVo1g3Peq4vo5OWFgd9LQZ8Ki419Ef2E9BftL2yamGO9rVUCmdUcBX6d/s
DAPg7YSYj2W1wabJ5rsusARlEWZOtDFOCuaVIT2uASeOjxGQeoQcwyMU3A9yfn0v
JIJQx97toJ8MBc0gxxEucxsqKvKd/ZxyjinyDAnCzPbIfY4slheQl1PRrf91pwVp
UvAKrNSERsCAA8XAhynQ41lrIONlzLkGvAUCdz+JA0hZkyHfov3qvwmkvSSR6cEB
IXrD4a42HTQ3shorMEfDxKgA1pTEnY/7JcUtzzMpDDm/BHGN43EWcdBktAdJ8dsd
f47BiL5kgwNlTDX+PQvgVNZ6nvjKoFZZOV8VPx7aeWUl8aNFSQUapHz1U6XyiFIR
29GdfcLUOis0Knp8WgqWriDolkxEmIcxafSrreBdFdzfZk7ipuoB6/3DM5vUkc3I
n1P1EA2HfPRcpenuCQFk8dFnAt/rpQSsbLEezBhMlaZpBrQDDTnbLnRjUL69Uluk
WgC5mP7zOKVbA6/Qif75sluYeIpjQ58CMP+vgFk8g7ALK+PB9S/vlkoLQPXYykxq
MsfRn4KPZ16srmTNYZUZ3KVHiq/6Tdbm/sTRYgXBq8K5BWvoCgEA1wh1cEz8RulW
6bVSYL9Ha3pzGZ1wN9kLSCbrFsKiYoTCWDBjA8mh77bt38BqYPq5zvA/k32s2WV+
xjxdh4GvNGdXegqI1M+FAQ+Zq4riFmEH4bi1moNxBBnv98J4k6I011Llla6A5cFM
weVl5qpj+B7L39jOzDH84RzuzMoOHSmUV/m7TLKgEBHG/e2XYAJn4JLyeierAHE/
Ln+17JT/UMlrlgeX/Fi2RoUopmo39cj7+PPIqsx4+ydLzdlhUwxJ1GoOWt3GRC/g
TGTlx5KlojCmM9z/8dd53LgU1HZiqTT7K9Y4O0EP9ArpQcWni59pshGBr8FJ+tBP
Y6Rpk4Vgv6x/wAlRHgVTBD6wZNGtDuD6dTelGff2SqcbGEcHj5KQFsBqLYo53gQS
iW3xfR2S9UoUpmcz2S7CY84t5RKlbzzSeC3e5ksdRKwWThXzi/XkDFIH+LJDOk1d
X1EoFnv/pC0okItoBBfK9HUt4HPEA6nwCxfy+iuKQBwEU8VLLfaB2cx7ycAl+PMp
sqZyZF0nfWrbUib6/nSdLoxLy/am8DtLeTlX4YZfOKwsLKZNFrOH4Nau7JwqC2ZX
W0Dptaiu2dcqv5Q/KtFUUzDC4ytWRh1swjqBI9cbjzQ7XnoWSFAzzht158Ox6y9S
EuJWCeOZsxDRSufxfKlOdHelflM91KoIu8szCHnQyRVqQYAoHJ5hd+ySPpy6x8pJ
EQpA2IUQPC1pJHQFq6X0/Fpf66Ms+mRRY9IvyGdJnGXiQ54v9/kwi/+ex7i1E+4D
LihU3MqzM10fDo7ajiFfm5P2IAqJMi4mX0jQGKC4JJZwqwUzEK4TMll0eqdd4V+C
gUUH/yTjhiIN0JWu38HiX+U+UFEpA6njItiJHSk2P9VemhDM5xKhdHTbhIElQ6uN
atju6VlSpWjVphAIzKWjDsGimRp6cs1ym2W1jdwecEcIv0HfQFFhJM1TXWWdqUYM
TDkJnvqjsa8+BFvkOnRteH/Ja/4rmB08ui7uDNCmKgY5CuV0ZY141Sdl9ExGon2g
8FBOtgWnOwZiSSIwtJRUNkf0QJD14im+sewoESA4XCYC3Z5p3+nz0A75HgYLpB/x
i1kvtloVgM7d49EK+gbo5DqZtp36LXpp7n/wkiFbvPrTnA7+nGs4cQrrefzmlRG7
p1uIORYDNtfYzmQrAjiiUR155VMpkWXz4mdjx91OUJh/hnyg9gRsYZn6PG5ZFbEX
W+N6ZQARquP+68RafvCNVEmJvNJBp2hti1PEm46W9AnG904MoHV8VOe+kmSNC1MI
LB9BJWtAoqAMlGXBza6428gYhZZmfR5zCtU+xEpM6a9ZC6FNZ8LwpluM2Ujq3AM9
UDkNedi7gZNFbNuUlIVacw0uRr4LP3c6p2H2gsvGfWImsKt4YEta+M4n6BEFwlyt
Z3XsV7brpZykvrsOSK28sbf0iJyk+DMxY4zTc1nFvt8T7LYXXE9fODsGc+jq/xjx
DoVz7C+VnWtZULdivxqvvu5xyUJVs/uz1zTsC2Htbdd6hddHJXAFVbL1OrX+ZTU3
/tD8f4AaIWJ//ZaUEe3s49B3Jgpfl4JxhbXrfB5azfz50mKvlm+ChvJxC8mK+r0T
IjhfZV8zN+6GW99UPFnjpsi5MMXRxMfNKyHD1PakvO6LxjclGhbr/x13PbrK6l+e
C53jjGfxRhujTlqlidGNB8L+aoFYXjpaE0ftIgsZB04KALn16oCRDJgtshla1aa/
zn42nQmC/IONvPMy12Xr6JFo3Dkqje9rtAa/WaJ92RABHxlG49G6Lfw02BcA0pqa
HMIVLWIC4os2Bhxa+xuBuPyEoZ7G4UWCu9vPbCfn0mSUKNm+01+lh+8Jhdhr6EPE
cHOpN5b/FDixqs+39C0kak5P07GQiyhlI5u2pPwretVjomqn/na07TsjrIqDWzEU
d+VBkdichvyOnvDUKRajIvKuQtbXfh3RIw4X23qeLX1mztS+FCfBHZ9R3BsTXq0K
JJaGf4FncuzYL0tzsOy8A63HT5a176yfdcvLTl6jyymd8ktKFmdyUh7x5KroT1Oh
YrRtahsEHX/pc1SeqfWG6itsZsUPn0UCxWqhz274N3vCsMhPFm1r35cr5LG7GIdD
jGXxZ2Hsr7eJRHGqw4pkOrOmKFrEgl3cUv5XFsMFDISDKoyLgWVt0UIQR+zQuC5K
avE3b034WE538Msm7JxFv3dPWi56yNBM2QdDW8OD2Sg9HKyFAmjF3GPNLUk7Oytb
n4Ckh6CUC3VCwqMKhaA5zlPKYpTxhghsTE2gFIgxo76LWV5JVl7nEBpfPeFMX0VX
Vjt0FDjrLYmlOLIK6yZioCf7/XLyWjpR4xSdSYWkEuH3+PdD9zVqIbOdfy3Zsy7T
BWbkJU+VJnSrDmrJlIaIR6x5tCnaUQ6paht/yDAw+YiDEdxzE2MzqSSJkiEtBkjL
9MDspsuKVesvHR7LeIl3IBnPDnP42V+n3e15gyULlvBI9q5nX2753N5O9foOHmhC
w5LskT7da+D4My2OBcAC6mdo9CmjY+Y/2kcJGXQcGc9WWQhrjgV9f/Fdp+Xbk2SO
6gICQfGAsWsklTjf+uT3QUMfWY4DNttEj/TrQrIpCi+KN9cbUdLXXujFC5yJNeVK
xnPKoiU3xSmy7oRrl1P4tGYHgp9zWq8O1XpUO2WuRL+aHJwcYmzqfr2JwJhHoyDI
h+er3HHj5HOBh4BXnl9hlLs3KVq5udfAVGSQKly8lOhZj7i0TReAQ61KtTMtEHxS
kYcwC5lrYL7qfcB5SD1qe43vx+rBmB8FS4zCYzVzrkw0AN4wK/b3uy9wj7x1vqJa
BnTuRrDodNy15Kj8QFvMz3xrD9Dy2eWgijSVxtU1tqtJ4bHKEcLJwsJwyd3KCzYA
dhvhrk6BlqvmXnGGuyqQehS/sOimH1t9KOcta+Rpnb+FozgYQ/NdWz4DjSs9BmTm
+bDt7mq6trUT1CBI/KG7ajpuhwMNEIVJklN4ZTXZt2z5jha07NyYxUpxtwtnOqPI
dUaQ3yvpwPAB6ZakrAL+nuUTNJwLhCkRcc9xJesyCwzSSjCdiLL36yyjEq3WEcbu
Qhl1HfxcNkbSBIEMcojcw8pjo4/ozhH2OCTJHXG5Krkzh8BdwS4AhJXpA0PXqLva
yPJylKE2YsdAy2ccUOen9rofJZaqHoS+2qIwRZT4rX7w7J/h27JsRH70MZnnmB1r
pxN4vuQFocX1WzoLA5Qxb8WEQximvprervzeqGmI4jMyfRJo32CPb4jnP8e15g5z
sVs/ocG/qguLZjcsoIcp/2TG6HNF9DFQ6P+eqlEpMcTwX6XwiWropWUgd42pmCfu
fAg+wJRFzDLqWHIT7iZfZYF3CJ3iIpqgIbs0IRmUSWXNAcQbBYOWLsCg4WgXNTG7
aFj92O/bWwLfgsVZhAJBpxO05O9MQHF8gldynjr7PU9d/OAP6Mbr+IEqv3iDAor6
FT0V5ibLtSVxqNaBvGZ9vnUZbqMwFPN2cg335vOIZJkmDQ+ngji1leNgEQk9wNGH
yPSIhrrncSHO4s8dUDWNqwgxBxWoMbxc1tVd1VOMti3uZR1DtmEno/SIk+tEUWAr
xCsoQa01FVBUZlw7R+b5QsPdUZWaSi5nGJHKrUWkLfT1xxsYfVIWfxzcMDbDt08K
YDuOs7m2LKeaWYs+TaQxAo46O5Ay2DVIpDiAucuIb/7FQwajdu/VQncfAgKQoXqW
Ilea6MsAZdKybrNCxnbbK1JW3GX2BRsU7xqa3Vc2Ok+WOaBIWnPycryiX06/z5Qv
5n1Pk5zny1xWAtEDt9w/siC00xsWJRAUIx5BD8L4lRDn0p5gdkoSP3L4FWLLRhpS
dmTZ77n/ReF82argDBt5147lGQyXjJXvyHjrtL6t+Agmcm2eTETvpi3xukAY5Zv5
cXkWvp7mI7umnXXsRfs1yl/QtZPQGSaykqdACuNFy6A4qDFmLU7gqeFAMXeLhulZ
8HhRiaXM6V+vXLGSkEkc2Ta8wLM4PBN6ULbGhH1etBW8KM+53q0yBzL+xPWbiisU
PiWKWzD9IhCwFS2f6js7mVNrHiQmJ8fh0ACLnLWvXCkc3lfi12SiS8DbOr1sHjPb
w/JiPnY9yCCCqf6f4CJLUx1EcTPjfLVjL/xnVX+3FBiulBznOYMoGcNhS6XFGM8e
JXIMD1c7H/T7ym+oiK4MCOTZNGN0Xw4TZwgCDR40/lu9bH5vqOXC/9oGIV50xlLg
tvlYR0dYz7bLLprDhuKaLE6uvoaPo2wC60P65d/nK1eFKnvrNggZr+XuOmW1625A
sXSp9ENorx5L5kMSEog9XyklNzfnENGFBQqKczTz8ToJsAk8WlqfUfNI4R0dlGZ7
JnvrjGxEWOjvxjBi4v+6OGXXCCGFGKz+GKW+X9rLO7K2t1HdNnHR6BvWjYaLexNn
vu8fGIahm/F/Ji52kLoZYn0VZcZ3Qqwg9q//lWNWwFPtdPLTbolq87OekeL408my
ng6e068qalcDO/yHudsn/IeTct+p18ql/wvnT+TZA6cDo/qcIRgqpG8+eSjt2e5L
7j0gtrGcQyPIzi7uowkVGPLAfSF//gSwc/P+Db+hhG+Tirznx1Qzxym3aHihQVZy
z1Jsg89ppyO4pPJZOP24B4OkxzA9QEI+zW5D+e5FwRdNtTjokGqvEXJYxxaSpFDh
brk33vBhB3jd3x5iLuRk5arNt8XfuCbreQHg/bje+hIYmiV7U3rIiR0kI1GzJe+C
LRPoA3OFsCxnkQ3c2CjgbjLBYyY0UzkVH020TkvX/1duJsaO14Hx6gHdiupyW0ip
ht9FEW0ChnNaQwfdevCZIvoh5bXDNsTB23qZHet2AVJBQ/7CAxZoNm9rn/+Qu4k4
/JMcksSj8Mqc8UHRahpw4VWLx4F6bt/90ug0gdPifE7UqD6l+ha30C+3pkhs3AHJ
EdWNm8FlMqhcY730Bvw3eNQlV1lcdN8Y2tma9k76OC2cVP5ZBWIZfYnBoXceQZG+
wazoFMmTFHl21zLJoj7pmln32TGy8dEbwLiir3R1VSeze8/x6LWHcdw/9n/V4ZWg
0cEJukb8Wrv9FuxI6eVYm/SbVTmuIIVz35dz6fT4Kpsir9WgI8d+Zeb6GCyANUlf
GBTRPG26qaX5GaVaeYU8bJUYRIYAIDIeALRwZXrJbutKGbFRsnKHU/ybTRo5a1O5
vH9k9HDywcFpzPDqBf3J1Kbzxpb2fAi5vB3D6pNToYzoa47B6SeKaejYFG4y2XZs
OO0fGMu/gOHg/CNQvPxcj/v00L9uqRqA3EN7vGPrpaAyMW6PRiuhRjiGKxi7AEJk
JxHbpX8DZG0Ksbr+pJMDTX5OcU1JznuEgDUyHi2qpkjGZEuxFGeClmjPlIiVc4SJ
D2mi6ltaeWTwaEmX82D+EzMx+ZWGJtJ2HepCwR/xAxqxfnJH+TzqnrqyFQzZokl2
zzxd3kG5szCb43efmXsYsjogqA1b66Pcuuq+0ON6/4s3LZg0nwsvATKFJHjRF9+o
BVDSwa9TJ5Lw+6fJq9I+y9J2d2iCNG/KbsTfp1GXG8XK1VAf9Qm+kfD2oS/vaCHB
cQB4Cbh9PDKbxvtzkl1cNThuf8RimoTpej0vvvrODzEtljWuPklfFSG5JrtDjNc3
YoFz84aBfDYhQH/DPNfmVOfR51DgXY+zwrGzxc0m/2JPcPa6oEDaOL6Twythe3lo
YGXfEGD3GC/rRWIxk37BuLZlnEzpdhELSJFwyNAfcc9TQfc8hjbUq9m+6X0TN344
LCZII52wMPUig1bkZM57noyjsWMYXkJdj6ptDqwKWn0C6M+LxrnXGAbF9TgLxjbI
wr8fVapWHPQO305CH8COAd+RnA+dhmgKTrZyeJIF+/4yD8LjrQvTt6oXBUBkVPHx
tafJ3nLU5HFM5Xw97vO7RvbVYnFP7OreyRrBs4u0WJ80PfvDmsm61tWpMEoCS9EW
dGpJpnKh4BuN9WygVptZaTIv/RNyam9+aLHtWmTp6ZZ1g+ZwUTRv7k5JNh7OrYXE
Vxs2E7tnsIAzSFirndEePZOlAByNW7a2xClmPrFEFW8kwQU7xRo33xytJxhZbsYe
EJIQhf1Y8pUQ8l3sEnyPq107syXqEnRj2TD8IJRrm+FNx5SkYq0yh+C3LMSJFdoV
Fl1fQUKiI9z2uyxRKdX/U9v4+6mXRZb53TAHggJjlqw87vcAXxs8gPg2OLhoDNND
FEKuKcmFOphT7r5SLnhFBu7vEezxi4jbrhSKf9iAFGCSDBIFHQ1TP0wDuYJH6A+0
/rH33sD2RNTnxUTzHL/qzvFx7n6+Nbhaa7G8SbLXVnIUkWy7cIwJ/fA2COmM4n7Q
Bqp1KAnjZoD+J0BE8+MI7FHOrjgQZYHACMpU8GlvezYuy48Pl1lsvklDiVULU2sZ
1Wy6T5Gy4gzeathwoYDoc2zbhe0ZK3V/Tlkf5891RXm+Q3rFobSqgH+eqVKdQFTp
xUKQdAD6kct0/34RnWoRFLXtv7rHVNFm1lHeHvtrL5AsKR84jbkZvjkgw+nchSjb
QkfZn6q1SV9Ek0WIhl3baYgGmUirZbhqkVAa4UxLMMjITufrz5p4olLWHXYLGnH8
NJCaJPcEnmSlkKb7jUifi3kPvmkkqrzmCnejz8iwt6YUXU6bLc9ew2xugVsCKRax
GggcAam+3fl7ekcaL8lWHHF77NBdr+xRrSAwrKIi+Sr5r+O0ZUf7pime9u72SdUV
XwvZM+lAucN2mBZmk+T13wytJ+vXBhjMln92Cxugm7y6jeVe2NlabBJBdxj+B7ZE
QIDTB5qnHg50qUoh/Xr5tO7j6+H2BxgZgRc2HQ6Kh7TETNHgYhH5nJ4UCsxCgPlb
o9/8AjJQbu+doliee33Jpz4AFYxVGQbnrdhoqG4q/k6XtL17ZQzuzZv957TPNGQK
ub3ufii756i6ToIcCdFqrtecSacUMUrr9nnWt9mSfWWNfbQh94bilJwGyRy4aJhd
GRmxbWK0n2K2Hfx1Nf5kjRxctpqhf31rOC1z6w9GVCvrLlwXQAWxef1Fc1OomAuj
fCPwj4dNNpOO7PxWufC74f88EiV3tyu0JRmYz2i8PVSCYE70XThai7SP54MPyQVt
Ta8BHfQ5JPc1V6Qq3v4m38pfjh7N7BnzBzjOh1vBWXc8YYP+RamoUdpVvVXYx9k3
Ki9dhuRTX3OfQ4+41ip6LL2YO5YPDrSycYgKXqjFfTJ2R8vu8co/9qsofXTmSNOT
Relo6hyhjXmwTYTvYKpw63kg9pphVF75vQs4AvG/SXEOXNSuI4TAnTbf739SmPQF
A9zHvmChvosvUbcr+qbYyt2xYnoKMzJfXw+8onFT4tWHgBhxVT7JKdJDGOGcEoOR
GJu4IeUS4k5yCxQ7accIfhdehbExwaJSC7rR2l3mXm7fT5xRyOXV3mKS2h+q+vkM
4CsVg0ujUlY04QiWcp6kO6Dge8+CW9/Ov4v4T9ymmo10Va+76e+IY7yAX/qnaT7Y
nUFFM7bAwXRhYJJJTmwF6gToviqMT4sEKawmgEpMSaFHcXiO1w/EC0WrLyWFSVbr
C0He9ss2LVNLDwD53dKgMkz8EbTeYQr2BSySJNNS3mkJg0DzsDqDWNRgFD29J6VT
oKbxtxPV4zn21hrpgwTfmdm7053swiP8YUScOk9butOXLgbXiuHM1VNsbm38X0mn
moqKsQUcsfXhOuD11Z8bUzb8MhWFre/HvPXbRkg+mrUXaxmO29kjR/p+s/RFMlW/
jv8HSd6gSQyJP6tVzR0As8C/7ojnc4mM5hKsirKjKlFGsDHoyn8atzZLsWCRiq0u
UHt5txmfxciAaY74RWc+/sffhEwCTdwVIQcKVNWhTDD7RSKQzAbGGrSCoERzOW+a
SCmrliWnzaYNnBpLSe/CRkvxE9DJyar99DZ6d60WfHIjed2ztHbD9tooFA9hSj4h
lXsZcuwZlkrsxv/kXOIBNb6Clit0t8waGyh6GTVEONgt5BmHFf/0nMYE0e4kxbAJ
Xb3bultkLhrvtJLS59OtCj5yCXSrRt78F8gI2kvjcnFfPplypdYW0Xsx2sN2HL0l
rqEZRyPLcX3Kl6ncV/x0swkbi16wLROe4Ud3nWp/BgjT7yUsCW1TtMN56wZvXr5s
AzdOuEbviIW0f+VTrVpLEdwWYw3YkaVhVmMOG0CJZl2ltOmH3SlAk5m99o2Vjg3f
aNsI5gwF9aoue/svUkk/6m0BsPh1XL6JTSnvPF/yNsAnL73M0/UKfnysl27l2F3g
9C6oZE806eBTkQWlEmWOkPldeOCdyo7wBeGudJYXmpx0g0ZGu4EP+v5+JQrMibS6
jGFPO56Jk09MIZf/F3Q3JUkUHAFDQA1gWWXxSC79RcS60ShZOIoda/meOJA3Bkc+
SbBsVUbfqOayznlgBaB72QTnA1HMYUEozzCAtj4ubtz9c1pTPTORX+WbBpwMsCI3
1UGJIyyTKVJBq6i5R5DVXB0Ah35UU8BBpKifiXRJRPjmDA4CNuHEP912cH9hCQUA
H7++vTzKiblORlh6RITH+uoWbN2jJlRB65d6AwMKP8S7OOMgH1IRnXpel5rGtjuE
Il8XqFxKb02GwoKJL1nW0D/HYkNx/8QLidAmVtpEje0dmwDd2YpkSDwTwXhv6FMH
eRMLAYAr5omKovlQsJPrEmLU7c/EpNO2WtR7L215G8SXlM5/PzWBX72uaGMpTKkH
pIY68k6+ntmygpqjKJGZ09kPuDjrPDOlDKa0t2WgItRO/5+7ctlLSRff4KJ4flXt
FyQviBiCDx9egJm99O1iRo/iSzYMxfnFy/OyDFutTGFrtIYkhA7kxSa7qnM1odtB
6GwrQbabQq+Juw0RJgWb3h/7tngV64YN73mmgTx1UFejwFP2JHOEUUN0NKoJyj6E
AZvVC2TCkEA48j9zhA8t99Fa0e/myJiWym+SfjDU+J1FT0ABanURVygCuQMMEzUW
rKRkJk8LC90utelzCWMna55BeT4x5YYtd41lLYqZ/uqvtLRMngwpTS4qZQe5o5oP
sdG5AffYx3rG61mnEr8Ra2bnzmDLk6a8mO8ZALh85GxT+s0iws+butzpyR76nq2Y
5S18CNf6QAm1w7X2W0OqYGmDvQhA9kLojTZA016xBCd52CjVXvNL8DtGZKQ5bbg8
pUfgiJ5C7opNsJTpar9+R0ux2fqX0usKl0t9QyuE2Q0N/jT3+HlJlQmI47rBSG86
WgQujhDqTZbtC3Irx1InzAl5u6oKhlRYUYg2OhBf3FBWqNUnEVjrsE7bsMr1h244
PT/kmGjhbNbXbaQlc0YuXLpgHE2BArJnSn9mDzNtquitjdIawFZAASo3FY/O1fhZ
LFFxwFJRQC5+qe+PPCpvYvw9j3zS9/CTI34Qy57rc+/pp2yGpHIoQc0UY/PLBA1B
S/mkzZQRRkwQa138UpIT9qZtvwL7XZFBgzth6FGp8jzo9ttLu00oiIonlk+xD7k4
zc4Dprv59YKSQtt10rug453lq+j4Pi+4sT0+UZaI6D7IdIYzbsbfXZDJzP4az94W
tRj9oLHwdgQbvjEuYleHo0bLsa3hHy757mAFSaWDSZ76KIj7bwAGNPov/n47O24w
v08KB3ul4zpQsUeIR4g7QoR5JexOMyhz3qXPW6ei4qSY7AJqV3jcqN6sr/ohTAEI
+X2myRNQ5LEvJBxM1reX0p0m0OGPge9A/wQM/wOYKs5/ZwdLW9tO/CuUWyEG/iJS
UzXw6bBRudjIL1KUsGpVmPkZCJGDgtBrMPW2nphZOGVW4EsaBAAZw3MR+vagovCM
AmUULYIoGyg0Ppgd6B+TC6M6JDFuv8r1TB83uHZMNZNiIOfvdsrJrt99sdviM7lZ
/WWhU5Tc6SCTbiDVZ5POL3XBBzxzW0+Z2DbSSDy14tstKCv2v7Gz1GVBuiF4qu+V
R9uURpzkHHwwiijgXrpdetuaOqCuXYuyzpPHrZeoK9RWL9IjrVLyfqbyafIcObAK
CjNr+OVZTOc37jt82MVlWRzsb++vDLw7sUFB8zlTADVnTY2xTMsd5xcXFSdtENJr
oFdnWBdmdzdRw8GtQiUHk6mVu5GGbXh3y0SCCARqcsXKSmYkJ7FHQReI9mRJAsj3
E/v8GOh/B+iRA4LpOndkcOGdzQGfPfu02ou4eWKEc537jpNdjUHIYVelFJDeGYK+
oWt1HUTcwSXUrEYZeMjfdSRdzUIBNwbajgm4VuLrZay4PAejNsyhrgiUagwKUTh7
9/X7kFl8JmXCLvSHy7dER+QrbJD1rjxzti39ysVBudl7jHh7TigFQQdZOUiB809d
eLkn5zlGEjAKeNDHB1juyZ1Cik14P0RXthNvB2GIEhCdFP1dQrfzIM0udFq5lV1N
lJzTZTOdlUFN372IToNM41X48khexOeYQLMRnvvaEgWT5fqqNRufgzMAiz4V2Lhw
9flmeVmISobgkzYiM7tlXrsC9EJeH7FLq2/XU0SWQegeX6hdPakXtgRWHbFxCrce
yNDCHdTFzODW6ldazvwgEOwsraP/wXuvv00+G13BCAkZ4enl3Y7g7XMymUrbsCVU
gzR1rqkGzPjF3QUaE8iEC0cCCzdhQnPP4THLZX53X7PPXg14ymSrI8AHOZ2bdmpT
43jexmM9YSXyG/4rD4sBxrJIuB6JV1/7b3ikeTVvFKHseqOQH4Is99LXMwwIaM91
2NolRgAoTuY9Uk0Pr7uozvEFfP7E9qtUS4DuqNTnkyUT9EdmwCoxTr4RQw7PoPch
co33eW4q3GRSB2+iGFQ+S6HvCRjJGGq1Zndx3l/lpCo992QmI7TDBcU+xE+1D7Q1
IckEdr0s7CI68Wp14brqhCARd92rNw4B+Uu9WpcfnJ/vBpBGsKJghKUY2OQMIgLJ
XkBhmTYMKjoFQI0oPX/yB4DdQPKMsjoqc6kxLsVqXt9/upVqL/kWspk6hgd1dcB6
sm6cGNDvvKDjRR7Fuz6m201igXYBq0BTh3qJnlRMwOok2DYvbZmjCx6drUM9R96k
lzEtxjXfAAwk5e0+Hqa8BBnL46nRQPryUp61Drf2c4fNEGuF/FKrpG9BBGreddDk
daMIOg+86L9ysg9yrlbUHpAg6VX9GBXJ3MAWYq6iSEdtShtD+O7ty0XA0CsXx7JJ
dG+WjcwxTM5OzXGbzMmutucsf3pI20bgT2TOUG6NoSmWQ05ojZjNh1VSyCOyo3nA
BcW5f5fO4SKi7aKwMBzcBIXrt5IXyqIBrJ5SqE6sLsamb2ugmcr7zcVfYkruvfxA
KYHxJpcFfx6C9u4b09ymbgFxcq31yvQuQkf7NyGuool1XpUDnq6PJSajyc14mWzt
FKug9Aijruidkr0i30OMgdrtY/0hAN4WmRTOvJ05mTcY8J9kMw9n37oJW2M7ewxa
eZckfbrv7oNeWURZ/8YS3rB7s8hKx0nv/dF6Zd7QrLOjTYuGF+k8P0lLl9faDA1d
0tzvH0UatQTonycZHhQ+s9ZUNuZhz8XCEGlaVpnvpAcHSOlnc45eDVyr5XapsoTl
MxJRkg1wZYw9UGpzxUYDEVmTELjZnyz/3qbjF1UmU2LLLuyzg/Jw/RNp39hzRHAV
OJqa8k8wxNgv8uLDq2rbsvmHlQSDS3RbukiwUGuNSsqWYDkdpks5JPUby33mYI6P
HIeo6ap4P3nhU5wdeKbZPmhWE8Lwg5OOjuE8fCuwQhRf9amC0WbaxZ77MPiDgW5i
HZIUU/dt68yIJdYFNUWOak9KyllzC87fTdlKzWR+DejwYZowJcMariGau+Lmp+Rk
Hub0D9oxP/6aGZsKA+cKbVbm6X+WDvRSx8b+HLFblhUnUaF0AQHnJfcUeOD/RAGP
443kFb1yVORSki5kAhOPqX4AIJwOmBK6U8YE0m/lbSCUJCYgTp2IZ++0oV6Ug3g1
Mw/yeXp4l2IeSn6HVy+q8JhHi2cuCWFqYR9JNWLH9KC3/xHDMKSBHWekAZ9IWjrY
dO+AOMTH4m8YanNRvaoKK6A62N/W2or5jmfM2nHfu4Pp8d6mp/NjysCynXLpFy7z
UmQWWc2Y8s0OOfggcZQVldz+5hlblJ+CJbkELAzeoduHLkonGF6OGDs4yhSC5v1h
jWtz0Bm2In+d2uSXl3hJPuwrJMk3Fya53JLUnqs10TN92qljnl4lE9YkiMrsLfdX
+q4rf698D7VafLfJnrvNMG0j2ummZGHcLnjfWhVtKg+gJahLXwc5D3MAXGmNIJ5K
ut+1IB8wwUU8IvXngQBVr1p4rZwDPia1/317r2kz4gC5v9PFla91V7lhaDF4OGAu
atoryeApWtDAKlyRO0he5b2A4Ey5Gu77ajwzZefQmZb6jgguA2WR7YNuFzIy7gOe
DJMFTxgF+34tGPu/M5W2xr64aPyojeFszB2DuzvbA+k/KhLhc1Zk9D1IPuWfEXjo
GYl9KuYMKXXbyj2i0VjO5gDMfehwX2+2LGCgIf/2oh5cLLvn+SNJC46AwCZCAwp8
qiGVGL8B2VTyLmThOyiU+3L4RxGgJHX+To7dGpl7eknbm6oApVCFyFWNrjZiKoyP
IwO8TwN0kVG9LUm/gPw5B+Vy0OQ6FBk6WgPsW7HNp+nI5fZEE9wwFuqBhnW2qbhD
8nxPs1+wU5ntCIgzB2dq3oIMiLGEvFlJTFSZaEbQX3TS6lECp1JQyloGd7k6qkmE
1KhAx5VeLwUFhmQ+dIwa7jjEfxcyVUQ+n5NZ8qArxCgzGvw2PcvfM4NwQ39+/NrV
8nlDh3uypNlMsxjbR24k5bJSdriIVC6i0HCOoZSBjIiJOLivLV5x2iBwEgyVF1Vi
Fe6bq7TGkwWDI/tE8Zw0LkEFwVravPoCjCWO9/k+cu68j4ON9LYoPcChYsJ6goem
XkkRX+WseubaF22KgbCgEJWN2jhpvFay2s76wlIrVOS6w4AKP8TkSgnK262souGc
VGS3kZSVOirHdZaC8gObDm6yXFYRA7TVfGD3o4SKX/jpduESVwrI6RjIIkUoDr4O
vKI8GswOXZrT1qA4pHNVx/WkmkyJ6PIHSXKIxGQCSTBRSHh1v+yCZqw+ENpaD3PY
6bgFXDgt3joIeGO08gnEat0p1r3JRDxeb//sr3x9q3/x+vRCxi9cgt5sJliNuzu0
C7EqEUjVH/z1s0lgZMbAEkIs5WIAjBvnNswu/JKfRC7dl6uGjegakrC80dZ0gx4P
GAbKed4JhAckbS1+6a2oeUBGPSgiVnu8KLixR4iU8vfHYHgH24X5Uhim/CgQtckh
YNn/Ex0hi6KXaBTFTE5EdA8AUPaAsLaHdO+UMjnNjmGWYtKk+TQdaWyEipKh+Elr
YwR6D6al+l0q+zXHft9+LTKL2BoPa/zAVQ9Ua6TonLHYNwXMuxtUb73jS6j3asvE
QB3o7nOEbs07OzEtpewK7lfSyRhkzSSnG8zZ1eMiFfhZg3JZMOW2YcpneApyD7B/
TKoPBhuUBCbr5qklx1RyVy+mycw9anORb/jJM5CLAdh+/QKF8OrR7cR6HbyQgP0q
A1zdaabt4AJ18CmCJjz4q3n5MYApt+pRE7Nipi7MmO93Jqekwl957DLAZqKCuWhV
0R/BX8uxlBzU0GlHWenBpxfuH2oixsw0hi5npz6yu5xRRNCqlG4LmHsX1QLfpSv6
bdZil9sammiVUcCkOl/yUPZr2MpqUU43/ACW/P+lY59/5NNO7EfvGvStNDllVTqU
zVRf4M1EC0pN6dIkkHoMWju2/kom8du24JTg0HZCLbzvwQYQZjEo1QbdIk2xqp9H
tBcAejZlBi/dv9KvG9LxLLCxfvoZEcAzSrENo1X7621l7HMwK0OqgF8pe0qXZSuU
BsCYtffAUHTtxAYufkLt0DMHSCohxGVZ/ol4UBtMkO5NuZ3S+xw7hVUPTQ0hLOzY
tOMxOBsdiIHIk4IqsK09Lqm30NFu0VeUz0MfI8Z92H4/z6M8QbKdiNTMQeivFYmH
Xsf9iASMJN29RscUeQ248z/M8SumwMBs0o5u+WopJW264z80TpeonmBD6L81xPkg
MG+TGb4WAeJlyp3L7KEJgS86AQE7p2jozc3NsJsQQsM74Zt2JDgLogktGcIoTG31
k20kHkLzciw3EcqfGXUkHrhdlF7TURQ2qM5mgHO3mznJcvXTJhjGlQ8au/qtFdmV
EzOpNwSUgwxo3nFgeRhChyIIL+e+wPPb70au0sN/D7XSxTcpOMzPJkyqUrkw6H1P
jmMV4qGwFqXW0FAeVwY6bW3dubuGLpLCGMVnIPe47qLlwgExI1N538nXTqydSkfi
Zubii58oy4yJWc8xrP0w0x0+Q2kMx6TtZC50T3Nw4p7CO/weRqdrs4lsxz+9DGLy
NHKlL1G/JPSm8eZmLHgrJhTmsvi/etB03OByKQ7VR24V8mHs6/73gMiDpbPUchbz
9KV5YtFjtTsrxMmo5lqgNaTjmZfnghZEBPUhkJhw2ZwutIDed3y9SixeD8wHhOym
RulQ46w/h/VMNNHP9AMBg2QmhXz54x/FjbvrHUSN3y3MCnQvWJz3maOt3AUFj84P
ksBcrkcuvYFHH28ol5MiwEWOhC2DcpVe72jL+UUCeKIMg4yx48qU6t9C+NLVQ5xX
gC/vrxJDOEKU9OciOQrw3dcOpbmzDAnfZw0awMFso+87anTVrgei756WifvlzXbs
QcPJmtPIFMvCOGP8hP46F7prEWNGuiB2Bs2EBvHncq72o9xB7xfixCXLEwIUa79w
nXXZZ6m7POlQ3o1YalIM7LWSyEhAUDr8wZK3v59D0sryOelgtXK3RRkmY98R8Yet
Z+ymPJ+ESsZYc3obB8HdDDfRoJVLsG1DoeAsznatmjuAR6NwTddyPyuZVvhl7rZt
YNeSudieCdWJVzqgeLrG5YLkGDSTKu2jkOUfBDcDkSe7+6n1phAp1/AgOiVlHVos
itHovRHw094radFVwOEEbIcTcPxuGLXBqEIcAnoDK8uZR9xiI2NhV70kqjJDiBxH
52WzruYIjNy2M3JePAh5kgvA2wpdI19fTfChUjtolyhfdsAxfiVY/QamGQG87FBX
E0vuAtxohWzBgZiYQJx9Guf91dY/yLqGP+a5nKPs9f/qFMXb4NqG/ThcGLWK2FSj
JLchPstkVh4EM/6/lEt5xCJd3XzI8JSQkfX+rX50+g+MquXD4+Mx0OyZ7QRgHiP1
Iq3xMFadX6/utlIig1Yx8YgkE9BEVkRLnYkCjg5N06I0yuBumOo0HsRERxnlPzlC
gRS+J0CsXst2zH+Cw/eftVVuVb0ZOGipFiEQXZiaOJNsat//lJgd0DVvfpeqro4R
mJF9/QyncEY4XPicweaClSDKvuTzviQ4/K5WxZ4rw6/akAPuu5X33F5U5fBprUp/
RuyPoXNX1KXTBlmseaXk7UNNEreVAGTmRNZH8R2T8rR9WPuletMry5/T0ABkexEY
Sx0eAjV5/p1SQfxrqt7SOKnG67Rpw1APIJNJaIlHuIOFjugsV0KLlRME67ht2ywn
n42I+2yPHlYmfNfVs6MrRNDVrnpHP0QFdsukC0L80zbVTo2KpzuKYZRXF8TvzFeC
oelynfgVFVbyEQktAzlo8N4cDCaYnRy39/LkfZY01T9geeDJHgtH74/KAalSo68v
+yRZ3I3C+LHLAV/XbOwTm7btDC4brt3i9oXaGpdbOrLB0sMhrF4ULwBENyZ1T0sc
imujrmuxL+zlyNkUu7bPb+4FA+tDURNBfNMBh32e2LRrMlonvx+vyCfws/QwjW3v
w0DE+vqiRFhlUwyJDqD+9BAw+KAkj68zg5k98b+bRhLDhEYlWeoZ1jxWVoLoLDBQ
dgB3QkLLJWwLjT4cD62GwCRZ7sZGco0qDsfj8bAyuIxL7kLaxzGS4fXUzycQfaGG
dlyBur9gOmZOpiYw3AKzByxEN4a7WYW9S62UpxDTtekKktp7nOf2lQWSKgBEr3MI
GggbIpLxGE52639XA2gKsR1IdcQBnGFQ+CMTDxjaUxGfJD2HlsW77gLXwUdE+4lV
vUF5pzwk+T7CYJIz343Q0wuhxyAq60PC+A8a9iXAQvMsKXdZMnLcmC65R1i+9SCm
TTjjE4YKMByQBikt3ncIuXkAvwl7Kng66W+hh+XeuBMLvQ+oMzkzh2KEH0AIhY60
EpUtLaCskTMWOC2E01UZeYvUw9MGmY6KTmPSDHFDP9P8yrmrKE91wS29azeTGKqz
Ca1VPknVVv18HITp0QbkhRvxm0DpoyAY4uYYx2Ina9F51m3kAOci5NevljIOfgzD
hSxo1S+zhzyyfsbJ0Pig5BPMsN4whd12P5/uembdvdUTdQzFOSbfoS1yfdJkevhu
ouK+Vmhk+WBlAvoYAOyAyG5gvQNrzttQF1p3f5oP/HcSdwLoxG8iednLx9mXk1KL
dWdfqWtzWBrpqOHEKLb2R2ja1k5eAVgMK7V0hThh8tuSPFN4jhB4bqKoRpLauVRb
G1wEUoepqfqu9KfUc0MwcOcXhV+VyW6XwRq+/LAiRaC1OGQFJxwFAB3AZvO2aCcj
CkBzaOVfTZaw4u6YhQ/drkJWyE0X7mk/q6LvvCML3xNycXzhkNxq6q3zamiIDcKO
6QPN+pSi1Y2I5pBKv8/FPTqI6DgiEvm9r95P1gqXdxYf3vwNyOt4ck8VXRCwg7oK
oGwTodaUdcr2pM64ymjuyzBs7hrYWfTmKgJeH2EOSXxHdeoX42qv02XvPuCHsj85
hLgZFhxQaBgleyIdR0s0B9Pwmv+w64KBNukLs9VPm4tMHFZJtfDvnWcOn7SCN7Qq
xF3CLG9p4faXlIXDCdtKwMhzxCBb+V266bs3Y+b/kGfkwulul3JHKrDXAa793hKs
tzZ26wtHGsMTZlml8XwVrPdp1dugN42z6G40qthlkFsa1U/bmBIiJsyt7LjOHdU2
BzWpOMnoBWmoyBKAtkQfm8dnTx9uMKx7yLnpnc47RSsY7dYupdeK6bFA0vPHtF8r
jz/yFTWgauWUxrAU3u/KMkQBshRhtzbaFz/iGD+uG6Xa9dO150ek6Hf3CnXbdFXm
NgL9ADV5S7oFNms8uumEOzjqJXl59EAyNFzdH2v+9lcV4i9DvU1frrtqELm2nnjS
wcaZdOBgO+Q4ZSedA9W/PPiNa52ZPgNwBuK61lArD0ZfOujEYmieh0cwsjKZq3kG
fCiMjHLDC+7dNSl5Fbz1kWH5KmVAxE/epnkNDODaLKb1jr/+kSFGIQ+sZvIOO1Nw
Z77xaRxFU08G+V2YYt2AGxv8WmBfPhIXCCr7MI3f8GCKyVQIamINJjPc02r8GM2P
SR5uCNeEnDoI7yH0sIHnz/hWUR/3L5ZlWZ/STKQPr2MQspUOLRV81SVUdfAUQhmL
BJ7nKblCpWdgP1PXT8fmFjx440p9DlBlKd8XVYlfzZg/hHXRIOWeQiqcQtzoqQOb
S/QpRD1+X5rQyPs2jL7sJw==
`pragma protect end_protected
