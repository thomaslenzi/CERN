// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JkaSxfg0CVfyDHXvlwPZ76LQXuZYuXaDHt6LhOK3v08zz/uRHJYB2doFINnwxQvM
VxoTvvHXEbSwlQlLZl2Z/uNpQbMTRWyq4JuA30oG+FDL5Yh7JjfqST/WMZao5Uui
dFcq78ODUkgSpN6Y1taLZzqvNNdUh5G/35X1rQDd4W0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31440)
7a5549kF8iWFNOSYr5KfwXxhkShsk+BdbjveD16yk3YPgwsU+3rEdGjzs75BXqby
qaIqFe+H/EyoKpJK06AJhbAfUY+mLivqVnD4AhyAoHUP0r2XEMJsdVBMJZ6JuXra
M5a35Toh9FVs8UOPzpWkgwk1FcoWTAD7bdgEEaRodsnEsQphysnuXiyb44fLUtBI
1NY8hQistBAPxplDS16+GkUs2cNcYvLfMaxkFcmqbh2BscKfNZD3U4s4LIXMXciJ
wpCquXwkbZ4CEs+9oldDaggFKvpSwRLFNu4GwiFRHGS8MktBRs4k0/endzC3yvER
KX+gCIqH4L5conuE+X/lrFFCxz/zkLBJ0cyguO7f+bed7ODs+xzyG8a7/Nu1NU6M
jC+yP6CUfJdp+vpacYu6Roavas/k+X/tAEP36+XkIFBWobRZdfLeKRGA2Dxg0P1W
S4O6X2W3Wc4jNx5o1rFJRrbpD+hecBXEPjMWWUcVEJJyO0LMdrdK57rFdtzkcpL3
aESJzTmlFcYhjWe8P65RiKvhNrnFapuVvtaspc5dCLEkSTNvyVc990vY98TJNH+a
V2kodRYRvyXokTVRA0zhXknzrBd8ujyqxMb6ozmFnGQH+cjZMI8UqMqJ6nY398d5
qI5KPZ17TYZssKoKWkq07MitnnPIOQUd1TShVDljdhi501/wpNQMGbyU9/tRKSJ6
wOYSfCZtaLv2vZReAhIVzKPUUoLMM8DV3dyZK6xa0cZvPlgyqFraTdebMhUwxwtC
X83cR6iYhNfNsIsyhBTkOLrbd6es1YAQ2JT9jpbT+EFvB0PoixF3VN4Sy2TGRcVS
VMZv3CPS1ib8BFDf+kuXsdqeY15u1Cp9CMMeJycYVug8gJFnBU5rALLbH1urN+5P
jmD+y5i7tIBkPbBHijXaX1OtIiuC01yAufEJX0nPRSAf4qPYFBv5Ealiqq4dxkuw
YP5YUR+xWz8XpuMHipkLGOZqXoSqa9KcDH0pkd33L39yexnR6VKwrZBHFI6NrH/p
kKxCWFvUXh+k1mV/b647klMTt6W1J+KNRcKn75DZfBmN5fgffLj6Mms70r4J17wM
0oEQ3aqBFjo+Ez0FP0W+mi0pVszgHpniAQ4/Izmedwris28oR6aFWymlBNnqEEv/
v5bcGmNq8Cg5Ef7fpb7UKmbOz13OCiH8H/BPPoBXPC3YSHsURfkzZGKTY2ABFiRh
qkvrwHFG/xXoEIkv3pVjD/SUMT48hRfca/ffyTUxhtcUbdcMG9cgBND/aN4zcHB/
TVfZyi969/U7NmBTPIzcLUCTLyuipKda0AnSZqIhdyAz/1hzVMCtIPEM7GR46Mot
311YgOy2vmKwnp59Bhoya6wcfPwIyEsEd9hH9OZCESSRI7Gu7ffOQwMM54sdhoKz
00jPH0bYvoihEAtUvg+FkNro+Ng9iHPF4QE2Vx6gY3glHld0uQTtQKNecKT9O50S
zf2tFzzMXFEfpeN1ZQvUc3rIUtHRYk8ZxE4tHivVc7vxAwQIyNqbMjEFlziQRQgZ
2NaOEWjBN6EkFojS+JL8NoBgtbQzaa4D5MvwpXr6PEHfOjieH1DN7furYb7+C36e
yqGYHyl+rbN1QYvi8ZMtma8UcfwUWXXPLY3FBwY2pKPatNIGjc8niyK+GhVpRo+Y
0RwUtKkc7EOgXMoRKfzybWCfE/j7ORY6+Ympu+RAUoS047mTHbXxW2ubsIkFY4o1
DRv44KOVfw2KED++olGJjlzDsOcbD6nmSHQWyBRFKoPvRxUtOXPCloF2n7arOTC/
112BMMEd16fRMMUN/23FJyB/A916r38pDX4U+5A1jbBHB7cYrezYILIzm8V4HuJJ
SM3jGvrBOY/2e5Sk5d+6I8sOaIyvZ9I1KaguKTzUlPudrPu2v4lbi/MtVI1a37pV
IKVQuZfv+UNBJT5UpyTw4heiKPjb45qlzA4ILapNyAhBK9UdAEFiFX6laDrxA5KJ
hqXe1SvkIAWbA8qhJCv47sKaVZpV5A/AdQbwvzJlz95GdksdLUvF7hvrxTHGGxab
u5InOJq3KdNax4wneBCM/ZhwQJ8Hkut2AjOzSQdQwxQ6CHHAto/HvXCHowpGVDUU
xePU9w/k7mF+4rZ9cQCO4TmOOt8ymEKGnYmb4+G7w5qxsStFj3URx9++zVPlXGGg
jUzYDaTRPy6KBdjFYRy1+Okh7Ns0pdpkewSCa07Ri6zYGg2n2oigV73BMHcZH17x
d8e0JERoFAQptPdh6r5FpQTTXh59xb1KI2sqDCC5vDL3cKmU1rO6e6xYT3K+IAN2
8Wjs55ZZcT9JcSQ7CTWPCKLt1lFUZkkwsN75qyvX5NSbXFYkZapoKFdFpKebnfEg
qO77sD748MvgSKhXP8FZsWq/kRsqKAJ3B60h9Xk9BF/BpWSbAXOQeb81mJX3OC4L
3XtTBXXmX+tDJaL1kVy/bORziVcixtMt0/jW+j91G7EAC8bB7MGaDIDdRtA5kbv1
rjv/rTv6T7/vPadC7P/FCg2RDAR+O3HcBxfF6pgLrxmnAgL+wtO72dkLm8ci/9rv
ufOPyQOWM/HUh34lBviD7hjW0wOpwkIaCtE1UYTaqYq5UBJJ65ZGB5se8164KSp7
lsMBhZrYeFgVc0hxc6IZglt9GnPuBWGj5k4e6X6Jf4p3L6Kzzi9lNU5sdBIT5vEs
2e7JcRFn7OA7jwr+xO85zIg3tvaUqAn9NfQADpaqmTtwJVpcwKQ1bEak687vZ6AP
Y8lY3jzYfO4G299wO27OlnGc0sqp+jR26FEAWUjlqJCnoZ9V+f99afLyLnP4HVHa
rSvTvb9kn+azpQfZJE7HlIZelMxQbDRxON2MGmeHeS2C/ATYxx+maQidnuCZEv02
d5G/yKynuAn9g6/CVfqZwDNX1dYFP3OvzhxhcPwxJv6zFEyIExNWcyR7gLfzrGzu
Uxl/5sElpCHqp8bGBc25pXVcssEOeNKxl+njiYuGYQdD7lHdXv6etomUN9NysImv
g79W8el6ZCUfPM+BoBgRbm6pgF80txsYi7xVZ6Wzu+SCEwDsq09PvX7rH5ke330j
NN5raTyBKBjqux1YmqVz+Sd9U/pkiCZJzzRjO53CpGJ91GbdsfMPV2/zXEszUzfn
TIIEB5sn/RGpTb03C2R1NdIcZ5FtfxBCukv8839Cq2TXFzKbELl6d3U5z7D/tbaK
unPvY2veYlriYfvC2SHaPU2rfHuKIBJT8KIQJxOSulRV0/7gVgqRqdxf+WFgsdc/
g8LmXdp9DZRtTH5BV702CgRCnlQbrMolswCqU87axjPvC3cTz40uD5b+5LQcXSOm
A2562Zesz1AC+4CXXqgl1yWxF0JQL7H0EEZ0E1GCYXVXGp35OBJDRyXwdJe1Lu7C
qe+UNS2x+5xsSc1ixr3ph3GkUDWv9INBqeKh+MQfjiNuzGP2Zg2sAhDz+G6bbcQQ
zvunhNSAPVpxleJ5btQLphk8DDYOiMSC08AY3sBA9tmuOaG1bHI8Ui30CQ8GREAH
OsllvaUIGbb4f8AjniAs2vwx2IFKsK/3hGVajHpYS5CVN+7Kcy5n83g7WD9RMHqz
qd++s6JPK4j3kqPb50rJ79ysNhFldXnHlfyAfmmEInyqxmVkNW6jYl4T1EWmTD4K
2kbD55fC1cIAuOyLlnKabi0WXXfeJU/UWTweHr7Rp0OedQAejI4c65AOvDUFvthO
ZIKtI8WCbJfHoc7zK+pfnm54o+LuQ+QvLWxd07kDp/k5Kq2JkWflu2jSFkJ9SDOh
Tif2yrrGRuABYmPrWt5MseuWHql9/4FfKVxpnAg9JlePCjLw2ogPdol4OJ9gnqc2
qI1VO8JHpfXEFOfHHeM4uWSkcc9F3aYQ7oiY9SelzNIHNG7NTa+NxcnnkfCoAPYZ
c7yBmqvIi369pYsXeNSYwZydKejmyftzR8X+vfJCLMSKPEYnUOobnUjSvcLw96ky
i9TgwjyI0KYkgmJq4g1rdCBP4HGDLaYePOt8CNLBZYAdAstl9a1tDPXkwVd2jtLC
SW62Q6e/Qkkx8ksGbhXGJIuVSfJCHNmmtX/+FkpFZpy0jKY4EJXjwilqbPxu8wRy
RrDYtMs8zFdK1LfeZDt6yJ/dmxT5H4ElC2LxsWRwYAJ4dNQ5XvR1kfWEcoFMsaOW
fi8FMQYwv5qfC0RrTUP0EQhhtF4sahhILn90RSlr27Z/3dlVULbVKIqeSAo8Fmz8
NtlnJKUYw31jtn/Wl2y8EgWO7WGQAteMKI03GQnV+X19oJ9PX4r6FhNoF7Z4BD+L
e0vMF9SO4g/GmBsGrsKIwUf2gibW006AS//n7YGZPijE56slu8qgx31+WzbC0BIr
u2HOZgZM8BYheiIb3fBlgjJSKvLxCYwxH1Ie/1WHlU3/CJZqrMyrl/A2sWfmBVu6
eDfvXEMYxkoECL5ewAzUl9z7mt/dhVbk7XjKXkb8LZwBWFWWo61pT1aZsm8vX965
uZ7CTmKgs2ODO9yxJme7qf/9NlF9EgahGw1HbgtbxAbKQ4CXU0ni0/P9WQVlzV/i
FdNAAt00SYQsgGJ6OWkocIZLUjSYSfTtlvbMh0e8+JQ+eRcocZ58DODZ45H4DBUz
3LjQORaf432QuwuLLJQV3nbF5BLPL1imzUy7S5HGLPRKBqYxCRRYLgBPlmp0ElJM
vp40vvBWzB6egKEinmNONDaJZxa6sa0VPc/Q4D0NqFncB2p8nSgrvwP3GVR7qp1x
/XwDx+ycGQnpYwWx0P74Pgo9/y8BvPGOn3gEFeFPhdaL5lIaA/v7sqOw84UyjC6t
rxBMzTFIzi6pEUqgrnjwzGdh4zk8TArV43N5/ksWRdr1Jhr12ibzQJlMSuOUo5e4
GKW2JgchhEJnWNJLGi8Nc6+l6EcRcbiZ+pD4jUGRLxb6Qy45nZHDciHuPTgk4ZR8
wi7tgj/WLVKjYbzsYp1kQVGuhWpu+Ag8Kv35ER0kK3B7LruGCI7mCqyUXrudrfZ0
8/LeUtgGvJMu2vGgXMZyTBZIG8Z0qgnTtJnoZ9eX98GKruL+Ofg4hzGBmQdKtNsI
J0X/EZoUg02UeYmYBqZtEEgV8OSYZSK7qahWaQ9umc+0iYIIgaLanTIbaBeYvaKI
KNeSokbGvWEN5nhnJqAM2IRula1OQWAZUrXByldZ+e4UAEoPERbtcAVIcj54dlsm
ca9LXmL35heDuacnexqLeJ4282qI/HdsDzD6CVwo4wwhLMRbbgY8ITGVR/A/nDGW
ZdEs60rkWKHK2ZzxHAYE354xj3fT5494pi9/eF4g8Us49xWsgozR3WWIR9ukZzYh
i5HIceWQCVkoAOmQRNgii2+pFbwfQ8aCEt8Ei6mxXQ7qALiFq09Oa90wkLmZmMUv
HoYk4N31mIsQAtZaKXqiLHdNcHEEOYMvW16j1QsoU94HWue39U+V9N5WE3zrtC68
aE/JzhE4gGWEGqSljn5j1UhEHe1K8EgEAsr7poRSZD08POl2br4rpwlLZRbAvBC/
Kods7wsOe6+P75q1p5W5JkbVjlesivU9b7S7POJ4uKaM+OCPz/fldePZvCI2P7uu
8zXG54wryF2zC/ICMc5oQMcHyNL3soZURtwGNgmJ0xd0rg2mvQTaBKuI8fUCiG5S
4VLSOcldarqxg+1TPQ2sAoe1UTrwZv64R4XyycWIY13bX7b7XDukiUQrXscQ9wDQ
d48DXKlohksySE1gIsAe/kUkHe6JBVcCTvkLkV9J4DiODFr+McldKUlpTwNonyil
PQUUQeUZl+uyD06SNDgrDiQ1AVgsrm8OqyJ2xkFb/bcnBtEg1790TFtS7or2tkQl
gYljihPhmco1259G11y/wljV67XbNUFbKVj1pyE/flEReO6scz6NXthhLQZjpvzs
F0HksfqLNh86liRB7DTQA7Y96yREtudVQsACPMQU22+4X6XtLgmjuuH15VFX1Otx
t04hfLeMP8j5AEJ1NRHBBprmDhcyb7kZhC8VBOgNnqh01MDdFWMX+6O6pZZTysZY
eXr+aeD6+viFCT40LMDDnGN7qBN7lAyZDb+SOoicNWFi9nO1Wd1N9yr8rOtAgvXZ
wg8yeGkUJd3tJVpc/Q06rJnfNaH1G7GUtQX86nsX6wE9PvfkjGCIv4SO59heo9rE
NlrMp/xzqseiQhrJ7Y63ejynfyz5/7fxds/0UkUEv7KNtF1JPy5kAff7pQRTKhyG
8KDSIAG09oRRor77po3zE3ImxfX2mesO9YdAgcr8xJS/jOrMnTxATDngNiTpBET2
azRysoKNtSuZ7FUDybpXhfXXiWkuud5I3UOSeZow6n8wFWRn1k1KWntTwYipJ4WI
PN/a7xKjC0OrM7PjHHl0M3s6cjGAldY8X21RthOXsureh3OBSZwy77C0nC4P1NgA
s9iLjmZM9FTNTPL4ZRW8es7/f1oQ5mmkXAG5zGvDBag1NdcOCnyHn83qPEPsB8mK
nDVmPJC+fXMzH0+XtqRmB4DIzQBwgPR5MbwXK9Ri++NVUBXxgWTJfnAY/tnP0U+S
kfeGI87XhXwWeBsa6NPVm7VNxP+koZ7RPJWfefA83ypdgN/FWJnEVwXGY0CG9RT7
Uh+qPJipTUVnkmNFOpulaibHZQrdQuztSe+Al2IG1OykQL6Es6s3IyzeSGg7FgNL
XH7ssnS75SvXwJpK1knZD0u+474wnnNOZrwr5hpUbS2zHP8xvSM3ysDj0ispfb/V
Mql3fcxWQ/RNnuMiGs4ftFAdHJaoqVW4EE+n1Y9VpIzdUx6EBVZHH1UYm9X0PD6D
mkNFActzyNsJIkm3orQZBUVPwpxz7qVvjpgUXxSemEGFwoLwHR8K36MhkUI4CcrW
vECE8n1u1Ky+S1wHsbgoHO56dIYGlIwipi/kwuxoznJu/vR3Lgpk63IuMmlc3nZG
IfvKiXvIcQ+DVgZQkYHvrHXuAUnHIIdtjXcbONAORYB2I42kcTIY3ZU92otwGkP3
X9tJddQ+GBeYfvRefSdehBHcgEwM8yXb/FIG5B06AoHS7Zq/W5+JaAToNVvI5OHa
h0mWvBoLwKo8YJ7DVyEUT9IAoUZEaQAzsN/fuZOwUaO4p6dPh8Uf+Gb5d63k/YKZ
d+6AacDkqUIXqW/lZIqopzAAH1CP4K6zcU/Lnb5yLNK0Pv5cd5fuNZ432WbOGkWQ
Ce4z3GboZ5Fb5Us0oRQvVQzYzjWUEbmPWBTKXHxD8YuiMH3jd8Oht3h27fqKYk0W
cI9iRZRPTuITbk9nIG7l+5y5U0kvAuaggYecoIK3Z/C0DGRVa7N/IeImssHtnaKs
NSIfp5Mpt/LFR9eLMKGjhaS5vnlTeEdPKXtl0/tkO+KRn6ITXSE9eVZljKHJY6eO
JJ35I1dhlT/rWmbxJZ7h13hfDWZjAHFxuenp2JdTeefuRt+vXC+d54QYqJTb6NB6
MZ+ZFwvl6eBr8tJ7eHxrCRlWtCvI5Stv++hAuUoZ+QWaooS6vkFmfLwTRIudy+UC
MZDziqT51EboQc9gOOcVFBKkCU+3vvKjCcB4sMHT8TxMnuxWxnVFSfCBavES1FyG
2CMSHcYZ3eHpnodRLx5sgkDsRy4QuJSAJa6JwvZimMZ44AsH5ta5FMQBobhonbhj
Agl7M1Ubes1m2M4dGaJqDY0E1lvCogI6vmx/ZyVwBomWKRN3C+sSuCFxkK6IcxG7
6DrATuoOdySUMQdG939GVSU+TCV4HZZBAij4l6v3yVarz422AN5Z64QZzS3XwmVC
Fz/rB/vTZsVJGsTr3IMbnhwLhjkWNu14Xo6novXbGQw3zuwb0jXejUiV6uRxQql3
IYU2gVbJJ/ROOd7ZAve+nXYwIMdHTRowHL9FngCsCNeUD5waB2QMbek9ATEDFTIX
vfgskOS0Wfami3jalpaviUfxtvrFlnobI8/mg0rPi62Zgae+LeEsEzibpdyAmiTA
bBkBatYXLYm3kSsFPlGPEWYMq3TAUWo4znAm1vNTgWpP4ED4Xnld8B9cnk415ktP
7+QQqLlPiojnHLa+XDvu/nkIO0CSxMeVi5TW8De0F1PcSYWYgpoqlNZbUupHzL/A
0aWH7fb8spmEiGLGaeeN/6LrZoetemotOy6NvF+InYB60KwA4h+JzdxU2CJr0C8W
3+PQy8ojon3tNtyBuo3fQyvCIdTQkuEXWmqudDThPrvRydS1Ok5MwM1RoY3Q33vw
gLk4kpxCHFz/R21DHz5qJzcJja+WznUOnICCK+CJff/CkZiMUqrTSDLYaGIT67VX
gBFnYioJI18eHTdrZkmIIeAtcVoYLV5QlIGwrU+Oq/a7dMf6VuNaYlAixcxfxfmA
SgqeYdlfPuhrkuSo9LZbAp6kyTEXpzrjxV7DpNO1v74etBMP41uELorUZAXbiUhi
SzJnBMQh3fjs912UMKSn8mFeuJwSkCQTLf9RfzYkWAM2zW+pcwyXtVHlKVk5ZgvJ
fOA6OVOCl36bglMtPIb2FrW5jaTsDO0FKFz90iAnHcXM/shCO8WxvPIlPZ3ApXHJ
TdFTCvaLcpReGP8Jy+ETWlfeArdRZHHkwUzlIrUV4/2A+kotztnbfB0UqqRbjVDY
8NH0DlWKgQr6w3VWucFK+bl0p0DiaXk3HERM4n/hgv5qNOuh3S3xo+aR8Awf3SWf
egB08MBXHZ6LBcisOsddUsaqb1atAlQa2rIuy5qv1HAYQ7IoZPN7bvJGTkS0z5HZ
vl/vkOy30YcakbCvWp61nzpt/6a2fl37SLxEaoWAMqpOB1FbMuZM4lVdM00+fWAO
MHY1atkAvyfvZXDM2xV7QO27+yNj5wjWsO2Wz3QQVZg4DvXgXNsM4zJ7gTxvMk7x
IA2KTWKjEMsANm0FnTB2GLP3lCcIQntRlxLeEi8oP+o1MHRxuCTzfvrheX7TElFr
yFUdVDGbFfnEBruJ1A0VeqyLcHqGK/wlWpqW9mWByIQxMaQL9VmW9c7Ylb2Agpyu
CMy4oTktztfYKsoHmUQO7vC53Jm2bAfAAYyQeUMlBD0WFTIJEZDoT+ubDvfpXwzR
ZzI74s84uyXSIam4idwAqtb5uqs2kXKQ1wqK/gwwg02qzIR58N8TVcz1i1+qw6Wg
IYIGNFk8tUS0JJUiTai7wNZTazldba99pfGO9lRLBf7Y/XXQdNk257iSdEp/ylxZ
B97nsm4jUrYtWV3b0Wd15EgFJJYbru7FwiqP/u2LDmi7LJhsxqjTA69WkikPYk9e
mfxKEeh7V4H9eEWfl8Pepx5Gd7TkUlZWsvkZahRQP5DBd8gEPXkD8kq8u5ItZat9
6M4w4q25n5dKlMSD0WqrK1NwDQzcfy5dQzB/6unnJR+Gl7zQV207R3fEeY9YDbmw
ueE/xgOM0ydYdGSfIZDRFvpBz5/D/acGPeQe2ggWe88BqOywcpcFC4dr/zHPFRrZ
PhoQuADH/o5zXIzGfSMwoox67DPZCGWJ/SI7EK+R6wZb4hUOTutV8DgY16pE7aYf
C7rHfmlQMqGGJ0wxqqeTdZaehuHfuV0SMCjWBECz5W3LnTit9LGiZ26IfTZzPiOI
L0fc+MFvli1ArWIhYYrV7i0mV9Kmm4RQrh6NPL4AGLJPchA3ObFsNuqbIX8XIgWe
+BBVTqEZ1KM1oZ+6pfAXpsyLnunGyYBDPHyDGBmQ2lHCGlfcsH2f5YDvBnAf+Xzf
JIR+Dx06F8spDA1tOUc9cDzIVYt6aCGZqp11LuZ5ivpOq8tdtgmWaxsUDuYGXWM5
PzEfl9yYmgOVA1CefvFebgfCJ7cdX5+isAKGIUYa4B3dNz6vgwpsd/iW/B819UVD
WxQel0beWPMqdEn2DanYiN4bJz7AztdcgKGj3jVOBB2JQnV5e+SKp9wTXFDtzQ8e
/1DYp2pp6v/w1XCfPqoW8r7Bo7bGddseg5t3ReFe094V7YTwv7x+uT8bF6YVJnsZ
LIi++A5GPpqU1iemGWjsIkq+mKN0jf3T0OeAWYEzNAKcMNGksTmfaeJwxnBZNvaC
e6/PNa7UfqYjXotFSGUtfQDHKVhXosW6KUsL/fiv+7eI/KtHv1tsG0WwrJ+Hsy8q
qlsVg5XUPDbC0a7wWkOf9pRndl3xMTsW4zkw7RI6h8K7ghIP0r8J0t7gEXfAZ91A
m5JdIl8JUwP6pTqfmG+7ORz+2NHQCIQvmC82kqjwRw9/60NDL0bKXg+H9dGQX1s+
VzFOai57Yjf9fWx0S5giSeY6/I5zgLjotBh7QG7N116GrQFp84BsWOkpXRgBriZw
RTlFb9xQhyG14mGwX8VUujgcKS64LX1nv/IHTj3kSL5jpqGAUAwh32qRXUaYqDJE
IZaNbGYd660B4f79PQ3IDKi8twqVrzp4H9OkDAXgA6nMqc8WawjV43A110edQCfj
FmMycYA4FqTCIdduatPNpH/L+IXK0q+uZvv9HoRfWUQPnYGsCUP9QHRQ6Uvn7IsE
DJFZrceUO2BdAwhcE65kz0nUfd0n1mC8UWH8PjHXUB/ff3cvN9/wt27qRBylDWvN
47bUkIl5fMVWGb83O8AU+1vnW6fCgZ//Z9Jfh+PzxZxssm/L/ybKU4RLNUo9e/Ur
6u8/ThZ4l4shHejmLtTj/oP9BKrFRIOscQ+V4a0BZZi85dQWU75hklUL9gepZ2l2
eTDiIE3fMxvTWjjUySeFxwVrgHgvPXMaAh+/1H3tf3Y1MygtItRDT1uXGR1DuBFa
uhoRFhfKdkzlkCNO8Cl6NwG/7w6Pn8fyx+UJjNT7AhATR05dQQqNoiHQrBfzP+7z
uMotw6b0XXAU/atkj45QOmD9lv35EBmd0lauChVE5YyWADlGKFo+rVBy7D4ps0HK
fTIsHwhjUta3o20Vcdy+SNal6LzvkqWWvxiYangwPAk04QPvDDQGCG0R7TcQ+Ebh
igbpzhtNipZuwOdqX4o4P5TPu7ZwRSoYPaOlW43XDwIY13Iw1KPQtlZequvpATwM
a9+yRYuO27LTNl/9cLiu99T3dMO1UTwV4TfjruuMgfEVXfEo6YMKKYNh9AOUeLKm
OzgNEyQbXONU73KKS8BbgC6biKB5YX4KLiRUymuNosEVu6FsLDdXtDtCPOK6rnnm
3RWvhF5URQe3FQLWbfS6rZAOVZXZJSdUXLSSbMD0AdwANvLC5QsQgUkpo51akAgv
xyePssWiSeCqfFz+az9jXcCub3/GdmxIQANktaE+L8nDfpTF60ar7q6yILZVq8Dc
SajpX3p2autYcGfP41Bzmg6QF4tPmsHoYnzZTdfJS7N3zWqFNex7VkKLowJTlNgQ
qUwAUcNr4I6nKW2nnFvT7FyNCzQX5UJEtLEuXjRAtBatDC7Cx85ZYYCodgJpaYFW
9JgqVozvqPZ6B1Gdt1ST8FWn37BoQ/WeisL2FQz29CiBtEeC3Au6cZ3swnHMkrXe
ZcG8LRCMin17Fqs01D4gGFhcNj2oEf10aewjuHRD+UHNpeONM7Dd8y5chIoQ6AEF
0g1IT+SPyrBV3YBUiArLTJpBnAXJO8WjkJ0xAqhgiR7Lyk5pcglgau9RTHDir4vD
MMmm7tfLf0yBE46cc+5KmCeH3WdW2O50l0mrSCwPxnT40d+4ktnjTa6BmqPe2HqY
X7IEKjzG03KpmPX3qi2vcwGUPkoxCx9BE9MKD4Y52sw24xu6dDJy+mO9x6BKN10n
e+T5l1kzeUreE+FRTieaZYO4sD/LZq4XGZllnXRS5DGXHm0CxzyZZvCMo2sZqFiJ
PHm9skjSHCzz6bKhZJXkBci7ABqjh55hDf0JyV59N3jVC8Txj5ke8mMT59lD2m1T
HWUNMfBe6OnNpmz94SWcV+NEyzNclBlfRRK1NQC/o7t+Z0Hb+2v4SP5aYfpnLmG/
aFXVQnjqHPK9PEuf9wS9z5t0bhwnht6tQaqFU7lGJMzM1Sgc/vAy2gLnjkT0p0px
yevq55hkF5lRjbuFrVvPq8nO6q88dn9ziNcRQljZT9Vjz6Q6Mmvbj5IQwycDDNYa
dXUvcXI792oFEsFjm46uOjPI0LDSSpnkxpr7jZTTcADdEeZ9tSJ/aTdhYuAVbOhM
mCCQx9Nh+1Mtz11Uj6+WSllunbcv8lYoT4ByQrBS0svylIYNqfcmq14lXB6fS1mv
/+Qixl3W05jmJdHeoGJNOgMvngnw70/5SjqB0+5UCUQcikzopukXwoPzOfjrKJM9
k+9Z5W2qmr+tq4Ka0gY4n8OtIafyNjWmYXTeINmUOTCjdk/CIHmir2lrpi0t0RnE
dY+GwqqkHq7To4DCmmfIqfvwfRjxPt0iF2L68ALcrw7IJy+B5+6WEmNjHILwpKGd
qU/2JI4spmN3+hgHCAxluphfNIFDPKPzo/BuXaehJoLCg/QIpTtf2ElkIESdUyZA
MX0fudteM8mSGHpDJHfKj983+VCM9ElO80wh5nz3xi1OeBxu5/UWDRKKLYvDjhac
+v/MPVJ+XepNZ9xcUsRFtNViRdlf4bpOGjxz3Nz4J0/Pzsrlt2YpZP7y2125X/4A
3/Jk8j9EEU9ViUYabFX9GFToMGJWwNsl5lQ0h+i6jMDNb0/mWOm+RjlnJJmB6QVU
xhzqkA0ZSBq1IUyIu7tY+ELWEuHZFqYPN1nJJKVzkhHfGUnYG57Julom34651xf2
nG2PQv9A+lUgvU5PMic9UPTq3IEt4rz5LA8hIYVe9GXGGAcbLaX1XW6qFmt6g6kc
jSwi2Ip5OJrHb6ltr0BYwbZkZzsPDEzpAwmHx4qe47WIoQOAHhO7FP0tsvyqZao7
iGzocuRLBU1OOPJemPcNchOsfw6xxsp42vovSGIeQTT5JsBxOXuW2Bng0Sq6i+5Z
d83QV9gpsDlZ/cdJ6RiD3XtSH6FjSnvUgnV+6W1xdMCOJz/T8gmSKRCe4QdA2d1o
zywck5KBwMTCa4JjXTT79Bw4fM/c0A8L1qNVooucNUs/ri2qilSxkgO0K9jHPhiL
pW2UTvKhLTi5iV6ZZmSl8nW+t/82p2GwnEHyRw82WxVjPcBpD/D4q3UPhB64K86D
O7HB8VCB5lKv3CyM5bieNeUnZMkI5SmuTXGNuS0HgE5mOh2ebEAl8pZx3u+UTjqo
I61rNsbAhiu2sgfMmH/e+yTvLwwKYtvqOwheXdAlaMcfkItPRHIzOQgzDMh8aw88
KXEbyylh1eS0HgoxtF3+vRkNuWHuuhg3/Dj7UxjgNlfijnwR6XsmjvTY0wptT9p+
J2lnf5P/E7+KgHGaWkyKwHHzBG53Enjswt+WxwBILwso0QxUmaVEy5dE5ODpGW5l
fGYr7K5eXJhU+ExVfpkQ7Nl8JnUGby3l8mdILIStkf7v5B9zxz9n0pP8f0DaIj4Y
aUubxWXshXSYyJT45OzRjooc5Odj3xLOqPGXI1DyxHlGYYgVC2E6IOw1gkybe9c4
Cl1QUB112SJ507jT34+pdlAdhD0eFE4mVcSndex477gmpcsfazaJT5RHBEZloSLu
Y/14Osy8tDs8eB77IEFJgw/co5CmHKLaWXqkml71ypyi7naKPiyMIGG/DQThGZ69
7dbFg7Q7vPSSLKs/YMThbf0WLHMk/HqK6+Oh8P6LV18Q2YjdBjtk8F197g19IOaS
w+IDoupNLSNFNEQ/cxJReXjATSnRn96OKeIWHdjoWAC9OFBt3f5kraHs1udhl1QB
qbG2kl4tCCD98dc4BUW2MYcRDD+wBdMGEWpBLyfeGRgvwp7wZAOeBDgU8B8cSIQf
x9+xC97+i5nwdJ6RXt50zdNaTOxObxTj2vcE+ivl0O0A9Y2xA8qFOFb4DFVZ9DBZ
6wbEcOI9LQJi/bu2IFqvm5j/FWWumUD0i6t1iC6LjgH5M37kGsXw1FVrzHAjula9
y+GdBU87JGFqzajG8shsvHBaySJtr0uw1ZQXKLeDNyURH/Qd3CFQUB2kEohxsTVz
tLfZx4fFPLUwyhVErJgCLEDwx6DQqzOO7jXJXuDpm/ezMxEowfRMVcTpik+tpBrX
K58F9kBDlYMT0G8QpgVQGtQAhlrrL+21Q/b+biCvKWs9PWyweb4Gzf7Vzi8yKcCq
PJPYwkDq1kSEnZjOzoMhHSElOPLv/UAfliJwHTZs4f1IJ+hLRfhkKFfYmpb70emN
e1r2SBfxi+WYaKPrvARczjlifOSNll1TSVhQGA7pydjyXy7JTi0NpjUB8zGuK34/
DOAbbLdh7+4N2M1oZbn90Eq0OAejWLdlX3Jwa1+N9DdtJuFFefKe802EJn1C/KAw
Cxxs7XpWgquta+hS2KPEycZmwIdxDxEqTfJJ4l80JGyzWtQOEWnKKjJ4X35diLuf
72rYGrL1o0wnWTwKTlm5ba12i3bM6ZFciWc4ObvZKmHqTtBpWh146PrW3BfxxXOy
1sK7UH5KpMrgTcbOBMBjlxhFMqmeajW24Gf/cY1CHEvb8rQWKrICKcmjqjx0OE4p
B6f73cOolQbrCiAnUjXQbc/szdZNIyueKrm2zyPmKDEefbEXoCuo3D/yze2bCtxi
6wj+VFgOQPnPC0mJ/zLswVe8eJrJj8X8U75Ans5e4EHyYjaHeN88KsTsfkN+Ojcp
vlfqSP9IdlCfUbKup1/ZcTAD5cxPa43BdO61rOLMWlU5HK005SW+gH9YCNSWjbq5
nIlkBOCRDvKZO5Gk68ffhDZABmUkNBeLu5VtBCn2vGPywYM7gD7QYZSJf0lEUMje
eBiSK0RZaljrc+Dig9/Zdj2MRslYGo6gTY4q4g11WITWPU/w433OFB4dScOmCU3j
RaDjorJRAmV3o7hJZRkjvhcH7bRyEOzjIrL7qcMntsC48LZzfi3gu4zCoZxryBX+
jODReNcLj98+3eKTzMDnFghRVFgQGX0uA8P8UtDv5nJimxs2P43ZkzxO3x587hkj
w56/diLtvhH/qgtEGQE+WdZ//FNODBcH9laIWPo465fo+++yUJ3kO5BW2zrgZVH1
XKYuwu1S75zzmVt3IFQd484LjF0MO1zg/jwsoz1sBD/ZjwihFR67npDLnp4XHGqB
79bY2erauttR3JM6d9BgwsnKzDEzWZ/fgLFRbsMWVaRJsJD9wk2aSf2bx7hYLtgT
FZ/L8yQgzWXtQhrCbt3dXNE2fFU4tlYOxO3N7522MkRJvldbtVpN8GPsNLImFC9q
P7RrYVRjDH8YYZtT2YY+KVJ6/HI6T8Sh5lC4CchnosNhmilyRnFWtpZLnEAkPXMo
YWuJfrBI7mR8zhYx4YC0PoaZeGBSFKyYYKax5YDcr0/+oOFmvMx0lA7v9IJ7r2SI
xyBriXZm0s8HcZoTqxIZIARh5MV5DX8Bl2x+OjoHp+5TDgFgf0xFZr3TB84c8rxt
isOlbSbiXtycoCogGAGqAW7wxr9THGkmGbi1SVIPTum+s0l4ayHgcZKg0RRE+WdZ
Cl1nSRFkH+GYs3rzjB08V1VUKq0OnKa7skWxzpnqF4XFSjG0QSPnOqeDzxfBD1/j
bpifH8E2fc0POnNfq9TnY2WhpXZmxRYEXz7x4P6Eyr4aKer6WPa7xaD0WgBhaJM9
b3r32kW542khUrC1YUao294YrdMn2AvZg4iLAcv4qE44fk5IwJT6CVKeXXuGRzgF
VEeuVMQNIA+ncXnT/8ofoWvLnqkrNc/d3YcAQWI5QHe3T4sX/Lh+JR/2VmFOsraO
OR2FrlbM70m+xKW0pK2v7k8hqVJJM5A1Cngx2/1uFy9w+cSge3uuyPWynA2goKaS
9mTJw2pzIriHprV/k7CW3DcL1szB7ZAUgGc/KZjZ6Z04jkKWcDTBHBy1BLKmO0st
/wBBjRpjNEW1jlAdldoD3rFHJ8lRVdIddihOvLWk/MdEOfS63KifLzzRUGm11Frm
IheNESDAASyPi3Ub+m2vIjn6X+ztMDUrxrVHViUll9vQtUqYHL5c2HaIv4IW6/mA
pvi5g3liQ4svN34XyOExKxjfJqi1kjSmDDu3cLRKtT2dH3ZHCm9LPYuzRdZe1lzI
qeKuq+CECqlpyQrpf/7wYK3kbynYz2tDchN7dPnmNQMRpYD0h4p6ywaFn8KIrf5I
QjdhrBA84NST0KNdNMbayuLtUi2gUMkpnaaSY7ZSgCM4GS92m1/zRFVV5GmgplLS
/yxCB0uO7aGiUr2j0pzOLNwM8RrDi/SdS4KmT0dBHOV+hYqz+wv4pHTMt4pQHNcR
+Zr/X+30/jDQOgGoOlIe6bBrD79jIGuFGI/omqyqpT76QhtX5/d/O7g/eJXrMd45
e3XNQpTkmnlwNxaZSdAVE85iRjJ3cWre4B/ApIynT58BHqhZy70/jtE8rtl4pb0B
NnEvf0WMblxU3HRALYNa/wnPwDjU2Wb+yZure2IpvD1m92MJ86rlHSTwsUoUq3UM
bR0HQbrspgsuw9EePeAkiX0HIAyQkqrG3+olbbSSX6mbpiX+ZU9cRjCb/Sw0pN0H
dzVZheuPloNtNiPMaVDnSqJn83ZEllDCdItNNFVSlA7ORfMYp05ERyHx/36CHa39
x2q26BdpjPBM5Ii3aHS39VhNO64CKJQEBaaZgcZXxdE4eExx2haaimVdofwNAjFv
0Pd/AbsHrjj+/rmdID/8Qf1SUi83QfX3nelY9WI0t4LMUnTatmyURDkTHWLta0Am
LCnEd3ByDicn/ojwQtE+sW6/vgmvr53DBeLbH25BvRuwO+rC7Da20uPVNdyMnruJ
H5OKc5BkQ7YJfkFZ5itqHynlJINSSegucDF8xzAUXV5orKREq2TbasmNUFlvSlDS
QNS5iQLkRhEeXScluDrK2pH4gELWpty4qRRPLXx1nbRZtF7s/Uv502iBM1xnyzaf
5Iy6xOoWy/KbGlAgujuIMABsStA4sXyiCbDmG7ObeY0E16nEOzje9USZ4gH4YO/9
KkRptVGhNhwXvjw7JJ+Up/2nsSrWWwiLTQnpZAzU1Z4sPT/KF1wqVe0TISebqzYK
Lyv8uKDDNXDJ8kMHDhUjwT/PVo4xmMkTLbvvfpTY54tpZF4gSYMqaleufVEyjRea
umkZ6n3yKoq+a+NlNX4Z9186umO6E0oA8WWO5RRwNYujpyWAmI4fTQQ/7emnio+f
06rkj9if/dz8W8lsca2SXXqNQX6eVAtxfz+zQm1/av8jkuZLqZ8Snyc/DHCEligY
ewb1BKGWR0WaTomUr+nXHKF/BwSjwqUohb8lkYcxf23kwvHlhi0lGKTd5sZpRk3c
CCfX/vJs7G+LQdKmtd/S85ClkJEcF0NLuZ7unH+KcsRoMJTWl3vrXrLSoDwV7A/c
XtBEHIPWYAMeTzv/OFztKloB6oVAjXSU6Xuju3I9u2opadborNnlDlYXmZB5aYE0
n5MFFfHAe0x4LfyX/FBeSLkNg/VTnxB53LiIh6WHxe8dfjQx3b21tHVwjbCpfyvt
h1lTKDdKjYCRwmfkwB2pzA8FN/SSKoe+knHPRTJfONpU2co0cbH27MXuhlOLzA5f
d4Kx7LphAKAk2SwYzl5DHMmKKprTOxBlzcD8ROlMGGLkhXsN5C8LUu14LgQL2T7y
9WRFYdMNXSPx21Kw+5P2FrwXhsNRzAgDaB1X0NrA+iNvqg0dFOQVNZx9a3qiOkmx
md0ks1rtflfUfmHHQhF9pGAWzrHpYb3HXITw7prTy5q9w72OXoK+xWbIPdbe88aY
vb/cs/B4/DMzpDAy5J9qqHAfmxnruijrDqef2yLU8U0+Q0H7erlHFQsl9wwwr2B0
HC8EvDV2DseS/kbEIZN8Xs/6lTdpVQ4QXL2XJe3MRrJXNbUUtht+36YCsvJ8Obbb
2KATvXtm87FkLzT3D1MF1eCUu7gm1+wV70J5KWTDDlyQ3o7PnMluaEBbYOoTh8wG
dqKgVJY1bkrCkFkD2ka26eVxmLSjlPYpIoRTPwDQ8/nHCyNXV63YafRFAksEfMHI
abpju3nfDHLHM22pHrLnVktTqDb93mM9g1ip2Z1cQ/aqODidsjvgMfKXqPc4SBJ6
XkMQ2BuaR++jOBtbNbrP/BzsM9D6xKjcBTdKfscH699Q/l0dCtVR80x3PVy7j+IM
/tf643z+k1fQWzkWicreGi1FcKMsouudJnbfSAisBIYROrUjSTBhUCfH4eKpSaUw
wQOtsc9/pcDdcw3iOqtMqxUgyWAbSFpwx/NqksE/NcqNI+kfb22Lg7fYz7bsErT4
IFe0sVjPsEqRPcoN3EUQYXwCrf5Ttb2SZJHhg/XfYEe/yipiUpkTGf/fg6fQugTe
jzk1t7tNDnO+wW0UKJsklbz8J2eaKILWu/qDot5V+99ssTgYRVaUomHxGmA2tf0m
BROpCcOpQv2xt6bj1Z57RugY4i2Pj6iuT/Y9GuCulJDZd7fiMqVbJySwhqXVwrZL
lFu4yzj2WZ/VzvkSoDPa5E8sjHrtUhkIN6rrXRN0wkeOkSXfCER65mxQYSTmcFWS
vaO56zMpozcrktBD/d+IIB6DVii/8qyLRDFNH+FWK47+/O26WnltegnDtiqIivzc
BpJxecTa06660l20NU0Y+a7QVthc0ReetoaQkR+74r93D5IcT62rQnlJOYM8FK/s
sVssh7MrYZ8wabcHvgAEC0gxi6j7x6vxF16viLqle+ZXZc75k9q6x3E+n2lEz02S
gSPEjAzMHquuA9bNBTUeiSVqwMwxgCh8VIhj80Nusj4mdOCQ0jGsmx4uGDZEZ+Iu
q1revRi2XRmXrJQOjRPJky9YXLdaxoed8LXS8irNnUZFQBFCVGg4C/s+BOOa8Gt0
s1QhtoWUEOiamD+7GTTSQN/dB1BJSid+PsAG7iUfIx7WOIYx+3Zl9R0noCvMKp9a
CddlItb8AWQbunw6NPK+Mp1tlmIJ2Bsab/4vGsp4IIfjM82Ndb8Q7upkxkw2Ag79
EqHpJ++56OD6XBWNayKWrFse00qmbylqTSFAp1UzW9Upi++Y9Bg4TTDXywUq3P/D
PVvgHxYXxhKKzyYYf1feCmt5nrqhLsqS4efQRDpl0JGPGo89gOImNeo5JYG208M1
Wfh1tHaoQC1bdKhlu/byE7xKkQBvxRvHWTZvRLRKX98+Opcrh8V6Zl2OgxSwhnvt
HmDRMFIYZtPUCfRUGNpJZY3V7lGxefXbgbMuyxGnsyDWcQG81IwacI7xiviBh5DG
8tqNK3BsNBNAQAgGO8uwQ7fNs32snXD6WxIwggG+KF81/GAp75WGvIelhR4Hpftn
UqkSVHNXBzlSkuoYTHIcN0vVpjWqPswIQidus9zfbG0GW8gE0Ze0fCffqXrdhkbe
3sieOWTHOQCrOkUKitd8QHY2cJdnYGnAsH17oJJvLflMWOAOliEl6lgk4LiygWoA
04XcEjEN8XuiBSHMDyy6Xu5f72snCv7fftIuWQIaXQovMky+TCkTZWzS7OLXYBmS
5LzTHRxdTVRTBTyAyKvdxWn7cTX21WJfDBxygwCa+3pYPNT1TSyANxyaiAmceyg+
UDyHSVklVx6iP4jAV5sCM2FiIQ5pzJR6XWqCz5rezISo1PmkCq78nWckrECEc4g/
JQQvwhF99hnucy4DYA9Bh/NxpF9smcuZPzSusjdCyRs7Tt9NsO+o1Gca1ppDDgmY
8KF8tP+5efyrNKB5VX+J1IrwGMI4TFCFz7vTeSVZj4R8nfupA0yNFzkugSBTslLU
f0F4VGeOnQeacuk7urTHeUR3gS/pqg1Rix8U4QMWuN9I/FVwGWv6Kvpo2gNb74CS
h0XBGx09vfU1eE2V7+QEZgI15CHQxrPJN3CctjrB5DnVViWuGI+RVSmSkkFOWq2M
jw4WbsXsYGwhaibrrI4fvpauBTyaf+C4XQ5nHvZYpmDqCQI1HtjmKXsSY83qSEnU
zwR7oGs7PLOksPDn+5xWLI5PSLi9dZsCBWWhoB98Rkm+jjlcajbk5RZkq53F1YYM
KLjJmt0QaQ71TP8tokEm0GEI4EGu0nT7AwEH7KL24BeE23/YFiYEQnZ4he2U2dio
sCLYGcAT0o5DidnPAPaRxYWoLuskzw8tCIqVaL6wGJuSKgrVwybGR/ZG33Y2z7wb
9gi8FkOVEyc+wPBBZjADoK3io/dfK8V9sCNHAlN9vJEaGWr8bZCN5LxSb5O3nYvc
c8WuX2SSbYcBpi0d1Pogvlw+rt2xPy4R0pwwMLE5LLlYEV7CrEI+EQEURUA/Y+ZJ
4ccLOO8bINjyjynS67Z/D2B6RYGGdw6EJhOy++h1HLZZWUeKDxSZn2qqGyVbWUOS
uRGJBOsHMms7W4GIY/tgNV9W93XMgJ3MEoXqC2jLt4NoGiM4F7aX3evGh7lwem4V
wYDrAf6UOwb7lU5PcNBx6bDCNI6Ov6R7T/Etee3ld70rJIu3kevXdZqolViPwgyR
ajohppQnYV38Kv2Ohy9jyVnAq/p24kSBpzdvufbRrJN7JzxGsx0sVhkrt+a/VUwY
LKJisNTl1xNmF+BtWqMI1nENI3jK27QU2BXRo+W7kcyTD2yOHHzB/fmBIl4v5cGS
RiW7JkNFPtfRwmEEUHwxUrEgVl9se/ZplLscZ5qd8mobgOkiN8s7zMGb/er9U4XE
UIaRMgYQ7fDTqS28SeNGqqJrr2g393MRxGtnTGGsA7h2gW3AKRjUdIV3UgR2DUPb
9u4LeN/Yels/ulCdolXWkQUZyIKIYwtdhpQghimMzjG4dlWJ5VpdCMEtvfI4knC7
Wvqwmavn2DX77OyOAvgNBQrMgeS7gox2sFyjoaVmBL4HW2WQj8W+DDxur7zzUuwu
p8JxCcinjJkTYwmK1xsQDFfh4IHsm6nH9SkXdJJXPFTddOenoRO8cRtx3NKS9Cfz
oQAk5tDClK4/5eFf+Xt4wq27ILm58n7WC6+606UyrYbMnBxq25mVsQgQoqFBNkAO
xTRpj77E2qfbIjWyNC+jvuNxhz2ccKIEc4GYzEkn29nsYd1+EPnTF6k75jZGs1gH
fvQ++cs8h9Yo69Dz2cblxASdRFPLkdhyqSeUgNHXeIsAWgUXc/QeOu8zXTbSrmZO
RNIWrvMCK24tuvdlP7QPUYV0l1MEy6pMAIRkKFN5nnhBY3KzbZDTCid11t68S65y
Em75qTLpDB9BscqQ2y2Xsw5g08jIDzbbnoqjRhZ2fywIfS1wVtrSpF6Ni+77kVkh
osvOCp8TjQaAafDSuK6L9kdJtGK6KN2jNHBWUTNGFQkPPx0iKt56qdf6kZbXKSNz
pyFUnzxi/h3TS7B5uOnNuPAVlkDeeIDwXezgepIHgKTZnACIHAxX5iT4Y08+rsUX
Je1lp9vkBPiUHUL+TngNGcFRZljfSuvpcOB+g1qW1UTqML1lxg00Z4Dj80w0FeXQ
0N3vyHTIRDwyjcf3wOshIVivc/ovj66/t1raj2EYwDOk281WVQIXXEDnyNCHTj55
utZM3i067C6csw7vNXFEQq35zAmg4ifSypSKR/X8teaN6e3A7WMxbLc9jbP+FvoW
9T0Zhdp9L7PYUBE3U9YklNEL0ZY3ZVZLzlrI8Bg/PYhPndtx1p7OmnnCFIBw57WI
lefOIeLgRLFgjkYj6MuTEiNyVimeiignGrgym1zjzj9cPBQIvnjU2uZh5hDLjJhR
NfDutOcW2wAsw2HwtkkEiThlEi67rdCpqiDzOv/InGuIVwPy3iGkkxPjdfVOebMp
4u+FZNLWOT70GUVixrPEQGCqBSEOyN2kGYXDZnrN7jkBt5KEOzi/fxKoCJaCz9Q1
+ggYwS3Ut2AaGmL5TbEHyyp8ZOuP4vkVmrqfTPHsb+bLjCnqJhQvttHzdSHGJMj5
W2tuyoiTC3Pt6mLEaMWm8gQLtXeOK9ztQ7AMSweaM9I7Z6JTB2lPRWKsNSqwiNbF
4wB3W7BsICo+q8UuIL140vj9tfBFckobYgu+JhqfHyTWHvu7uXJ1d18P9nGmc3BT
FYZSkyRdMnaS+ll8Ua9dVwztp1V9DQLp0ZKYiej8zDkelQOAY/xDciDXMVO1J3hd
eL3l7Ws17x5kCSv+7O5xvy81Ut2zTARbf5tfF4dbuBNNLkT2G6AZZLU1XmlPmen1
3fZWulJ6sUD3K1WgXYdQcbtMgBUL95QW5EAoKqfUgsiKGAZ1paScHN7lSwEDbBTD
qEEf6TAtr2VerNcHoAyiBCD1i5ra2s6mYqfVUi/8DFxjI/clCSWcnkJVEDNl1ctM
RgTUDskbwpMLxklzTr+ysqT0xDRGZctYhshBvTwuosKeQOcFeqcA44n5ulWER//f
QuWTUtbYPGbprukxy5ae4AbDgjUTS5/UbWwfl/++M+5108oHEe0H76ILGEHux/Cw
NSlwGEruP+4V60wxYUa9bWXyXV+QG/o03vQwaWUJEUj69l2rjTBUxwJV3zUdbp4R
6213hI8zU2xKBbfFwOusOWbOzAmjLSf01rojKSlRo5SaVhwvTbnIAF2SZUdRdRsg
gCExq4oopxuGFwvvJNhBT1plQxQKIBaWd+fTFyeNVqfXW5f4bwoFiKdPplU/E9Ho
OlRJkM6moZw7594cLrbDqK/8yNurzRo+o1PTZhb9Gw14cZzlswUnSpT7sTIiDBrg
cunYEpvvC92SewwqdSnAXX+MldxW1grmS/RJ8s2vePk7eaJAYCikm6Lv09lKE1oY
MOcX3SK0s0PcAn1+PIjiatdYygcxR3WL9q7/YlkwZ9VmBKHZBtPOirPQdvVRxjJz
fvEOBZOD+Z7liz4n/jLneVi+ruJqH5+YY5+HluqXfS07QxF5RVQjeUN0SH7+H5e+
Gya1J7l7oM7PzZOZTC+dw3crau52lY/+qN5FHFgfh4yR6fsB5rBSy3PhrmvBpbRU
Npe3NCYCUESDeJ+JP0GNPW6E6CVivsBEL3Ap7hZ3DJmD5/Tzby0vqeLZHbjxfZ2P
S9e95GZTFoUqziSmKD8z82SZ+9LnscEmOF6FQWqS/NAgCvzcLvAUPwDsXbE/7TRy
hzLBXYXgk4BGWh8kCvW1pILq1NwfWIC79hRj1OxnFJ1Nw8kC1nRywGBKvTJD/BYa
IKy3ShuMutFdUpfOUv2plZwfV9Y9lAJxtLK9TBCb1Wpn6x77nYF9LnBwBo/03QMX
oiR7lQrs/9N6PGpgCuF1kTSj/vP7JDkd1RF9oRTS54SyAtynrn7mG4w12/yM4PuO
5eOVAEuWWOaeXdUqEhvm/w0hT3tAfP4691hS9exCzx0iBU4dp+R+e0T0gkf2RXEZ
nFbRq0/H1RopeMDTpHvkSLYzHvXredPr6Me7U5D1j5+6+zPlxyPS/DuRq+a+x7TA
/132rM1Aubry+dndlxpOjcDepyTNRIlPrN+DWZnSZ6LbWkAygVSsmxaCXVgdY0dM
UMMj594Gc467AK0xqM/x+EJ+zQwsLDOdXTnx5mNm9HE27zho2KnwgTkzbG/VOWnu
u45Iyi0hTr/MRPB3Xwznu/Wn1dn8rvRhzDffjfhV7hHouw4Wf3L/HqQMcfO4eOaA
hyWIKSshP5C7GF8EQSWJDNOEkYQyGkuzMe5f+Qu8uLgOex5pnllNasYCZJgdnuO7
GAHDTeTGMo2qkVqJ1l6FHpYOk2u4TE9jQd8G0rH5OiXtKCaX8nFRem/Akal3fNJg
lQnbzTSJIRpFYXRUhal4gNm84NuRV3+rcWr+yrZdKMWZYZ6krDYzs1RJHpaBS4EC
bJhkdlgMcVoNb4XArhJWzJLGtb97ppnPbir5o6tVhJnbBkUslA5cpX+6uKvJdPDD
Jrtyq2SqdSuVpggGPtT4wOph11/tDu8Oty4MPwUtr2wddXEd/Meh618HFnHWmRv0
DxoGBq71GLDMrH91HfHqFxvWnaF9macdKg0w8OtFfpvvG9nRt4nc8pGkna7nqmlY
7DH9nnMDRD0rySu9Deg46IRNhyCAs0uY3TQ00O+Xrl9Ghs+YYpJMtT5Y2zoln9rf
g1XvnPEB9T0I2IHxN0dmXwOSfOopYrisXFQ4filQzSuM+R4NQhfQCZ2Qejw/OC4M
zR+s+tak+HrBu37wZiqE3sHajfQq9YtxK32G1jYfmWbPddu6umZwqtqwFT5R2nzL
TF6PdObdMJbX9O+HTJt29Fs8rh1t5NnE4SPigVzd4kvfPDtQ2XmwrmLYRmR7Gc2g
HXFELAHJ5Jh8NcvNNYmmDS1SCZ5WBMpk2HCuq04ZY6LA6Iy6XKEFVCyijLZogepP
+gEcnr5K4w4tfZHL31rxwvW1052gyLBi83/KkgyQsPpoQA4ix3A6c46dVy+VHMLI
FRX0LVPMzuGymFN5yOvq3/DO4QTRkRbcG3smcmV/w6gxAWGmwiHGdKmq9ECuI2M9
reybIASB8p/Ge2H+dI98zLTlRIFNolGqpdfQZrFrx6gNm9TpavuzoNhfiiuK65me
fWyBUojd4w6zYILYKeYdhdQRDv7UDd+jZ9tnqHUKj4J0zimrPSY7tKWheO/Dfejp
GTLO3FHZsGM1S7Cz+1ojC4J3+skYGqPKRi5CWDIDdI++aSa+2u2UaDCSXrU5/Etw
h6o1TlprMYn1dEzbZNtQST0ghfnEGgJW1Up09Zy6bBG3BMalGwlFdqxWSfhw1bLP
sGGluE9HQrwN0R7csVRVcoHnmRoGLfalObLoK465W1Gm5sZ+ku0yvF35ijp9Vraf
nDzc0PzKFzUWV5C9sLFB6E2T6gZg226jEgWxtJkvARdzFFz284y9VymkyFwHUYNc
DjxEAFYtBGPyu2V39sx9B1xrCO3vlhCLX6+SQWPMLzAhiIwOHAfoLwZ3T5YHFKco
sFXd5Nd9RG2m2ajfklHWtr0EqckjvuthR0+g+ax9DM4fNeaqKnmoIxHAg6075CBK
8/U+gS/5yUhI8SmzDLmO8sS0OwPvq3AhbrPrnLwiasesCJ5ZkB+G+9OEk674BPZ6
K7iCFKeXZZEZx/4ZRU935+qBBoGwVRkk0qokmatwDDQj8QAE7/uZ6hvy5kcul1sS
jJlYnIyzZd2uDcqFGmDorKboHXNIdPrh8oziIUbbgUJjty8swgMLRnqQGolffeVh
O/VHDPqZFkHCiTktRhdFmXbZHbFZYIWrLR306bc4Prm1kveb+2r2GsvU4vdR3w3Z
fNJSj7C2vD+7zmRj1mwQxBP5g0UEL1jP21gNrxPYpEV72lMs5fkhZbHo0ZC8vyel
C3Kki1QE6FTNZrwYZnKVebLKA/VN8BDsCOSsfgZzORLyO36dMG8DSC65yaiUcugy
DDCrzokBg2Z1PNClBmYxbYn0cRDH1unpzFKR13j75vCKEG2YrrUsniwGvhEBC2lw
UdOdtM0VRhCsIJaA/tjQOGfdjBjvPonw/abypJkTCWcMwYdOMebUnvs3h1CaW55/
M+Ynz2lc28YlBhRkPMimAE/VZv5Db1xMXxb8sFh0GEDfLvlKXXamP7l+fX6HMBhh
pvuKgHOO2b4L3Uvk5rSwyu0BxqgPmLP74l71T3jrzju7+LGRBru6h/01vSnA3wiS
lvL5vfhEEj0YgCmjh5lCIrOYJTQvmlQjLsf1DJZZ9eYkaVSRRdfQyiD5tVjXHNrR
26FDJt+Zko+3ArnldP3ExFuckTVrniEyQR+RX4/xa4O2K2i+o2AThIrOkp6yPHse
KlCd5k3COMapsykSacTkV8oyItc59L5GElkXLbnAOFcCzQNM2CaSd4IZbLoDnLVX
9u26MwWTaJfIWGxPqYMgB0ewM2tB2a/UB7ZkoKx3wgZ5bsi6Hi1vqFAazIjW51z7
URtfoy7v1dhHW1Ehm/gkMP4ifZmqgZRUIUWvEixvvs/2G4vtAf1qZf5/IrII2V5j
Gy4aIBJYZIa3m+i18sQysJ6FNOGoopvQ87bf/ZYTXUVOmmXyxReFwXFfqkrGgDCw
FD6Y1DJZXzWwvTSYbiFUykNdXBS9vldVHGjFghXkLa23gk+SQo3bQ9w/wNfAR0OI
tVTbXFvFGP/P/W1CgDrg4GT5QmwvC0ncgS9zDBAwRNzHwJ9qvOTGt7v4Ix/TdyQX
FN5XB/LFzrorXVjv5reRUOJpP6Ri2y7TRQGltQPbJJVPogfMtprMJIqX5TqQiu4y
68iQoRPEAAEXpkvilRF5arffEwQXyQPyAClXeY/pBC0TFXGtZLGQJG4VkyvSZWTW
hI0clTLXnELuiMPKP5Z55fBtF8IbcIIetAZPu4kKTwTkQX6MJkqlDVvTeC4jNuJt
hQpNKpWUmWF5O1GoArvqkeCeexs5beeSz5T3ZAanXtTOm4vKTGH4/clE/x+GTGd0
RFuxboKDv6ZxbdviIqoNe5qcOocdCojXl4sqhpA6q7bpp4G/8KqDFpbqBHgUkNuq
jEgPaHfwbl5Kir++hZrkYDgpiIYeWgikfL+sl+0969WzvoJhUOM/kjVYP9YS+MBI
pjShrWVE31ST8TpD8nTK2i1amkXNiVjRsbnYvDlufzR2j1git9sKG8XmWnwAvFRh
OvYp/Kfg+GiZ44u1bOnNY0QpU6QHrrbOOLQ6cVuYNEkoelzd+2jwbr/OuzUmiwZ+
hku4x00DImDIFxM4Yy9e7mO+3FY8NKtlkg0AJtkjKbVbr7J6yJJT+NgGeoJopJEq
tvU563nRDxz7NJPNq5XTIDwlIqw4EtI95pGvz2KARh2TgqD2i6CiB/tT8Mwk4PnO
jl2XMLuVj9GOivO653ATEfWtaHv8InSnbhj6jBhJFfBU/syNjE+jjkcbso8dW8WM
hf7Z2WnSu8ZwBqj2IggJ3CJ25m5DbuX0eW2FIZafM8jDXf3KblFtVT+zdw/RAkPJ
gCuUjORi10h4RL4sQRao4ZiLSzfLZhuJdH95kKQ/8uFcoNeHMvuA49HLRGb49OsB
25dlNGhSaEL2GhSOwTH/9SwRoT2mj1cF9QviOAmh0cHUgRfA5aIPNnrWeCWkQ+XW
V6U7YlnVkkdaHRF9rA1t/Ig8FYwdvz/sH/FwZXN0Etp2mtQfpBqcntBTIllJ2Xli
NuK++wV9Arl+cda2+eQSO212unGArp/Bs4B11jT64WnQmVhMpoXBDmiKJcAxWdUX
4Y1TJZYUf4pHn3Yfh8wud1Cl08PXsKFwQ+dktjqrt1Mboe92OTbYc+XdTWBv0O8d
Czz9rl4FiJFFTp4Ojkax0aLbL9VkYfYwD9BvaekDrOLfEzVfJN0EtwTPBXk0ONXg
r9QHE8QAy0nKjAaaun/BuTwGxSVhnXcs5ky5lnAi/UGLsAGsooR0S2YWVcZvqAcL
Tanujt6qVlD+WtCzQgrt+A8KtFkREYHcklAEfWUan8iArgJ6CybwnuJoPcwCjQB/
IZ1djHoarNQNFtcHVLnVZAeP25LQF9Gph8cBVMfEZ18LrZlzZoJtUHVlBdSH7mMK
k6oElq8Pl8A+BcUve8+sg0FDW4OJ6NgscVGbQ+S7AOLRxOkGEtllgbGcqqLcTZhh
f5FweH2r6Ni3/VfO3SBd6q+8GKOzDmj6tU2UytNSbjWexySAMtnUJ+lTVO6rdDq3
zQT98lqUcEU/6FoPHIkD/l7moH0UiwveYanHm9vNcDgZwyKTyiqVbV8dnhoyNlb2
N0X/TXJnqU7VNKuaSr9y6bpj1c+L9RgM2WuemYzQzKLPiFbYbi4YwYd+6b441rs4
dyI+MSuORQBF9unuusVwQ9MbDDc9b+37wHD5g0UZFD5ktLCe3W/Emwf9g9tnXqYg
jGjqE2x2jdbj7TwWOXvOvVaJSZRRS/rnmELUJkRmKWN0TaGq26SSh4UERowysHum
w3gi803CPefJyXvavsdORVGCMtVeExFo/mUyJQ+APyf0byVIRn+6+GHRp7lK/dB2
QDyMqrcXseA7M1g85dHtDHPxE7PP0xXAclYDb+w32FaZZb8t4VXwZoNxa4srVB9P
6HBmR6BEqDs6LlLZ4TTcH7wfEkiEspTwKugDurDeOkEDe+4++PsSH712lhW+Uk/R
H7vYApkbmSt+duWL4ii2b0n6krnBuTizjDpSNSmDhJkF2343Jeog+mnxkUO0nDL0
n1o1ABO9OqUatwgrcwyXuSsfisf1EXBgBhreDYzNpb49dJhBA5AQNn1jG8JcQ0Rd
nwoob5BVeAFoop0f8ByircZVny8TQEZBiqlE9GmWgjxmvR9uGfzWqw0c0d5lJLh1
8HeSRXX8PIDjD9PhwjxAOw3NMLpnDbnvR3Pe1dLAM6lI0Ynzf5w5+ZsF6zqOgWru
/jZnUv4vKmUnNHtBPWihpUFyyvohvVi1vD0FmHk7gs/G+p8jK9sZAOGgJBavd9OT
55XGuaqwo0KK7vwxKWxe3YXS/ShuyjJKas4FC1Yz3hXc7L9EBCO7yN9k0V8yFBFI
Sbm/qNscVobZwSDJa0LMcoKAbWjiuW2TetnCv8f35vs79CnuNd8JQrikwB1PIgpl
LrjI9KvZ9/p1Gq3h74HtpgP2nUYY9lZjpYL5k99pwxFdcVhLqXbf1gm1qwQqYVmr
SruNFQSEU1MLIHbcuB3vV6cKnVjTKZu6lSksZ8IdwoL38aROHIWqBz86TqeyRhCI
w410htd4dopv1aGNBwrQXvmdIKP9LkZInB9Sx5b/o6C96ELwLMYqfA84F+fDF/7Z
4Jr+YNMTMNezYGYv5As/ovKzHeWaM7036ll62fmirfjqsajj2wRZIykubwcJQ1jP
BwTdDeZ7xIsSX5W7FevY8IB15DRrjMeQMtO5CrRSbAuF36oYFdU6+e0P2TPwA/CS
eJ3KBWtw/LnJlTNCYklQmirP1iztyI1wSStSN5CPXe0Uz2BUyXZrbcB794KKCMgB
OQtjx6bE2GexumCQLk3XVnQfno7uGZtL5OP/wlOoxm57VDyTaPVTDwJxDOThxFAD
MadVJg9bbHKL6gQnXy6JDClcNcHa8scrMv1EruACSLmIiKJfQ5xQbjbLht5CDeXu
BUsNuKJmwYlCzyQ4NuNiyKDmytYPGOV+OpWHyV6u149bCd7qC/nrtByFOm0eAEaq
xuoJzKdNejLk3RsDNmzmDI3NqAJ4+JDhDsjGKxa7LqUB24G6B0qM1n1QHtNy53Yj
dg1wbdHh5NzOc0qKXnrs3a2l13g1DfN/TOuRv0aUc2Gl5MGmo1VxLhy/UCwDpWBH
W2eYXYPadGsvPLVzq7PdQ5YgjIIgjbVO7AytYnKEJVxyM/S8zSdwsfIw7V7Lc1BX
Mhk4njYlatsaxpfcELtc/bgKUW39eOeqjUxGUZzJW108xKorF9G7QZ9GsApkUQqE
OPhTr6d/fJdspJkxSvNXUjGR8LBfxAumrO1ig32B6M1MhYIF+1OOzJ7rVaGJC0dn
RVviOOiXNmp4/ziQXLTga6D/ve28sgJ5DvqVXHRHGDgMkxwfjkGDU6cSusrhmVXT
tmT28sUSm0l8lVGnKXtAxacz8JXn71qUFh9GCpTgK8LrrczXIZgHBuf7yZYtDs2y
hs/GYx3zfU2CEz2FmlDcnxawk4+9inP6H6q/4p2g6padfJeIw6opKEftltBz74qt
iHteAZRCCPhYAgdbSKu1Kkowp9/nFKyzV9wxa68p1hzDsGMpGSIOmI6EzgOonWii
iHkvBeATGNJTAfdTz6N7K40wULOfqpWWMsExwgbKoDeoFgVm6bjlrF2smfMim1NQ
DG1gxEjS6w+3ojvEyxhcBIKeYb9q4gmkS/GnpiQaKeIegQEDcWdjTR8UmtzgH8CM
YUKu1/2bLZSM8jfVPx5mRvNDduxqZ0sNJpLH/2f2APSnhAkq8gwzaVHcPDtddADs
sdWpqv/HY0kpMfjiIJ5hIRHq+rv3UQ4SwWUOMQKitrCrFyVmmAfWFYOE5Gm8jnAW
LjTu04/XiDDIsPAaaviarYlGPLghey1SH7LM/hxYP8eT/bep44883Z5arhh68uD6
DqYRN2UBznGEO7Yqw0eHqHO0dhXFvIaaONd/VzSqphVP6cH2uBVU0+IG1vfqURPm
0Z+Qg5XydtUtH5vZwW1r2liXWTmUgxufiyTL5VdzZTAXlcmokwhRNdn67lHTFNKx
hLQottu81h9bfUI7ISn6p5Yq76a/30Wz2UPDLzCYie4iSUtbdLjosWRfOs2Qh7US
doYQsCH+gBxH+GqPV4JqXAP6rl8kmpxd/rHZhHrFnUtv0JrSYG1FjTNuwchQ/Ksw
nNqIlo0ZsQf/p4BBcjIkFhLNq7UmbydKdETIBp+ycpCIgADAETYsUmzy26l6+DHk
rHmqvxnMS35hLsOjb0XPu0RymH92rZF0Jz83SElajcA3BiC4dZACcuaU0rSwHuuU
msj31AQaawLxL3GdSup6wFxrjEnW5/biN/GkMsGXlajy28dJ793R4eRjpmosig3V
1zcXKUarr2o4bJowq4T3Ko9jMTn15usZdiqxRaTiVecWjVu3Ns7Bk6nwWU9virat
9kCOszXfXr2uICdq6nn1q/aYHuy8zLxMNq+gSsl9ulE+p2SBjfiObRHivhM+zgKz
5tEq19JIgWZtoOLeSLjqWD3wGUtgZIMPrGaj2fDkVqx/uBpUiVUyFwsrbfUsI+3J
WK8H2Ql3fkyPqOfwLZtz2SgRdgBs9cAhKibq4WF3dHbcdOhf3ok0wwGCrHkWu9dW
cYJCEeQcn/yoxSUCShUba0My2oFZUNDVd6+77gAOWZz7RRBGjX3fTEFhm8zpaiRM
WFiDYy0iVUVnKepb1VjNIkYtzGX02GilnYHdfFHnCBptXHRDQG2XmPyYk5Vv19iC
t6niH4OegvvTmZ76C385zYy52UNBgv8jnONRgxe14EL/4iIodMLy7+Y4nMnpiYCF
o4dPSVHTi+8OtXBTgCB6EVST3P0TUoMAAksM7qKCNFXppVHnA5vavFFlcj2r4Nc0
FiER3KoqSHNT2ENbDXYQlZ+n+vVpv7z2/LkSnP6g3fH3PqZqzWXtkS7yAPpft16W
DoNxpS3qBMMnfDXdUzP4m2lMxQ5HyzkHI1ypY0MkBe09PmR+BvpKCuVRMmIZ5LBB
e6nD8aSwqUN9MZ0t63CG3pnx1bv8XJk6CWoKpa/ztPfpPqApNVlNZnR2762a0/OM
02IKLoNEGLWSHijGiumkDNpYaDsTYruDjBvcH791JfOHL3CK6YtcLcth0/4y0HnG
CG+PeBhJZxfi5Hubv4n9cqAl+g5OrOQ1MQCyQfwi1whTf04iBjD3BEMkn/Fp54V7
t4qFDWOsGY3+o7SitssemiEwO3jYUPAZ9VcZFjsgXjz91zJHLdIIr+M3FceUMvs+
ucLueCBcWq5XnsYRk3lacleWJ8+wTQESwvJca9UWMY3MCGqXHqziGqUoscsHiah5
cAE+nhEoZvsE3BI0biRsG1VRbkxq8rWzIFR0RoKgyo8fSkfmUBhFrQY0UzXjkI0j
s0aapnP7OtBHpSDj5sS5Ck3nK+7n7NbjQ2UE3Ty3t+jpFtHSyjjFdQWdfGdkcLge
N0rxikbRKO853hy7YM/hCWQ2O3pTTCFPVoJYIxnwzPL6T/pzTcx4xQ8fWeVnYOHg
dpKiyxOsnfOP4t4vPgaB2W1tDqOlqR4lU4NncZP4RsSTZ3P29Vx2ZWx8F7wUIrzX
b6RI7gp1lZWgn6XWevw9ZcZEkwVxhUXBFNOfaoZT161L7kI7h6S4OEGSs/9IOloP
Jo4HH3IwBjIt9Aq15252qE3kjeaf7w6nsnmz4VBYQkTpPepKF571qGrXM1p4AoIH
8G4995s8Duu7e/mUUiDqoIvG5ylz9ow1tc8cJe1UL8/YqIDv//hMGSst0mN9MXbW
+7DWQQw3voamDZyI6yWM55db3UOLm4pveKzxEtze3ssovB8hXJc4cuZuRiHFctft
fd0upfuLKGV2Ll3vTRk5mRLKtwfsS3/k9QV8UvUA3WATMLRcdQtRj/jUbAMSMK9s
9OueFWiWu811U+vu2g6I7k36ttc9S0SnmclrPDsdINH4Uj2V6xzV90Bstuq86wB2
9x+tMF8IJO+ZSRxzVM7VZfUUZqnTiTRrqCU2ExIiPcmpDk1WCXppnDwSo1KHE5g5
2hlGJx8xX9CHR6JRYijY5qqNJvAfHpxJlnq0ycaaQ4Tc7JZKLhl7iVug+atz8CMy
keeMWkzhtP2e3aptaST/PLzcygxhIpqBYpo1PSeKQyERTIOpnzGVt3fG7XVhh7c3
0zfNkXn0MdUc/UkCRA9iyJJWjJlA80NqTVytN8rCwlJ0Z/zV6eidaJBiOuof+OKY
UP9mI99RYFRGORcs1oTt456D98nBNIUQ2OpAd6W7i3ZwJ/goT4E8kSwieCK3V9HI
EftgrIBvOwyLq639G9iMjGFd/gVeyM1iTOsLcinOil4xUUUoBMqBscBrlZOQLP50
q4c35xrHWMsQJbFoGqw/H9cSz8EBJxlQJUYdzw6U2EeTZfVqRkSs/PZw3DmkNX2s
NKP9zQq9OEcr2B70oeiAbK3xsPVQpqw4Au1b2idTAVxFVI3kr8qoilBztoRd+L9n
k9i3dGyVMbGP1hWBKvXR1qg7f+7WFDtvRbtXI1GbB04rJWw59menBvyLFy0vmA6X
DkfNwIhE/lYh499xHuWKddCs3ghaKRuSLR0Zs1bpEWuf61bVwUQdlhemDD0+NmeU
OFY2yCNtGZyAUTeHseitolPt5Ytei52Quu6u6HORN6uJ+ieWKHAyrJmNUab0Efqr
RNrhxGjeImwVBiRE6iv779IVo+zs0W6Q0KzoRJSJSCGDHSQwzhLIybuaTmh2cQln
nthOg9xebE+9tegR36TaYQLaom3NIH3veBhrb5vahwJ6/FbeKLcSBWoi76nWuJM3
2nLrKkCkOVTE9Zk8XSorcm8wJQ2QgGoGA+WT4+/wvlIDe5Or5Iuhr0UMU+P3ouVR
iW2yP++3sONbtRHi+lr1IFhGZ6NXyLUPsmPeko2r6B+1Xg0g3nlVouQFxlEi6dqC
9egksC+qb9ItA4u+5MndM9Dvr/dvqEedS9b7a1NT5SlsRuHmif41/no/Dj0slI92
mKZF2SmjHXg3Sl4WDFfBweFza+MaWu5Sg8vxWUJ41BJKRhNk1WbUAtUTuFyDxxdK
GnnUSQ0Fs7Hq//ViH3LZJIItyae+3R5DHudbLtJdhArcz/Vf/2j5ZjuzLRa/QAxA
cwg1f6Vnivifo55u7Rjw0FhzlzhWLOyUPz4PEgCvC+8/EipV4BJBQKsIPrM+KsZT
M4Yw7O2ftXRM4yrX3kx50vBK0FpDBRkDRKqzrTXWjDu8QI1UT9sOB1QRcgZCD6GN
VV38luVDewql/y20NkvxDkitoyZbChv1flGdbq2gT30XIMH4WPLUDcyCsSOb7UmW
5eOtoHz5yMETo7XT2R9Fe0jci0zsehZsjYNkyt6ULaEqb17G6za4HuOpEQxx8VOS
3UPXZePnYYFaa4Na3tr2eWqzPXphN+j2TxZC9G7swDdlsCETCiDwlhPmasSJRWDZ
Z52w5JcZURm8GgYvIGrWJCob5dxuraUImZQijohFClIXzFdsBbZxlYXZZuKlyAgc
RuDFAtNsqkxwqQqr7q0oIAThu4iRqZe2Cc8xbu5HhE+JbozhZ/gq/aC/7bwrcHtK
XU2DPuO8MN5xcW1/yh42fp8SqEEAXbXfCHIoXYibOwVSPQ1jISv81uISkpFYmQ7Y
WsbbnXDyvVgrD6XvCsFRVk/J+me8YL6j/1fD+Ney+1NRziYZ0v/uOUcdvJL+3zvf
Y9vaPc5K0l6dX/lBStTSp4t2U7FBy/ShGqbLj7agX8qHUgs3E3FgV7ewC1mKdtYU
QnRwNXSDhJggqFBCBtXBccp3Np9cKI1Ldjz0Sf9RE7bdez1X0FNqnRd0YIghGr6Q
gsS2BtirYP2go7PDXLbJ4O1f0gULpJmCs3R3lhclJ6glE7gx360J2Gd8wAHyF+fv
s+pYc0wNjK+mQZPfsuuOcZ3cgGj0g2boqX3kl/jXBhY4rwDS28gdu4zulQ5KPrFQ
VLw2KHete/zdUAmsr1GysQ7Qp9ItVNn2hkcOg/Egk7EVbjPtz1gV7XfjZP+S7v1V
mFPRUMzzBxACFRsSHrlW5aPLhUQre2vKPPfu/n2FiR012wpoNfRH3PSW3crBH3RM
WELWYfNmLH8GOG0jHWTO8eTk2ZtL5mlB0IDobEY8lfpX6ebqWi9upZ/GA8ltENO/
DjKjiYJorQt11yJnVolyJtd3WBBrPJpHREaDKlYpL+ROUB6cSGfdGbeR9hGCnQDX
DGw1RoybjOn4dktGfxzsJEzq7NhvWQKnEnxIp86EK5yEdqZW9vSh6MW+o3k7oQjB
4oga6AUmfslOJpuWzfXzrXBqgkw0mPhKBkIOa/hyMUb3V2FeTLqvKfAYmOnzsChX
UoEPTQwv9eg4TOzAc9WxUo98mXxBbLbJJzRhHtlDjBqklMrk1GB9rbWIT95NoT27
WxiM2q9cgUJIt59UFKwGIWgjw5WxXphPondXUJ2vrT521ShFolcYTgCAykd2iUif
aEsZ/+weKuBGFplhWrNZwKW21eisZQoEKpblCpW3jWKkljREM9AYknE/jd+hPD7y
SA5/Mav/OGHCDsHiFTp05/yubFWLXG6M3vmMr4/eIPJ1xgA5gJI8FAi4TS61tGkN
BeiAp4it76MAWWE0PHVRAGv1JFlm/xBsc9UHsZCCiLFi4TMCVxBii8BS1XU4QtXJ
yJU1nwO7RfC7ky5GX7aEfbRDh6+/W0FOHEVE9xvBSflorLUDl/1UQC/tnl7jgRT4
pzHfya9Jbb7+xB5FA/518Ecdt6GNguLO0nNtekM908aj13ZDX0T2or3ED+GDHBHt
cIdD5YlnznRUzhC4842Vp8VOBOLBauXZRInai+sTnPvQprxu4XId+MCoP/4mWYBP
Yak8XG0ByO4fVOqvLJuXHa+PKJz5W4gUqV2f20gPrRM/LSYC5hhm+YqkqKcRJlZn
NVrNeHEGF1Kn0DRLD4vjFrTwiHOMmWvIAkH7m3H9iHK5Uqky+zdnf7im+ISyLQax
75w/SqwctfR4rl31k0p3MSlGKJgDEe+n5MO153MRyFV1bgvj89+Wy2kN1Us7Wky4
Hi96Rh0fnA8azb7Jv/E+fuJDTE6hJHucUvW203KLso1riRSuF3ttbw367xkSJcTi
Km3Y5zBunGRHvRCiboVAZT5LCuEJFaRxiyvVmtc3lzcqXB2Ba07WC0MeUXgC6eNf
hxMz+ei8DwjsYLkM31ruZU9ODc1hFc2/DDX5K1Muzgsa6G5GPrtvIeg2WXYJpU0e
3Uxt0Ze6/d920X1PQZsIQo0KoF9uVxelKR/nXVTgQNQp+zTKwJEj6gxZS1SJSXoH
aowNl31xxuOhtW7ZO+pjnmLtlzbfaBu6pUSHtPyd6FbabBz0b/cfAv+frLu2dCQJ
bTEaPcuaYxclihtPHf1I1F5m8zGHmnlCmy1xuuacXHd5T/Ud/7JMMX7Z0n0bXtMt
0HLvrdAmNNKga4dfmi9DNbV3Db61pwF0mYR+wQZoCPycRQ5QlltMWa769hIo/0mU
kp9X1WOsr8v6Wb+8ZO18P856pbS8rGShVmr1Mys7R35Cn6KAIY9rP+Lp9IxEyMvM
gibMTN77P7rr7nE0Y/9+6MV3mkV9FHOkcQxCZMHYzlxw6qi9xmLJqQxUA7n0C8d6
nyUSdwYT/5pBWLlZ6fUUnO5NZJAqx9wu0RyIKpALaBfvPmzPFoBMSMkjtG9VmoYz
mAKYQX7jPGpROo5Qtzs21JO3CCR89Dc6kF4NjQmv3piAzGdUdz9a2BxL2obcwheT
Zzs0WGUJ12W4Lg1iC04Z7FzmBr/dOIy6QzCN30A4mC6JUaab/uhWVwN2PXLrXC+o
BUjw+hIDgKvDka8wmwg6hqgOXgWKGwPYMDPCbETWR9A3uYipkhi5mk4vIqwkNNSi
elXTGBAiYZIFWfgnEnjhZGHD24Brrnx4ZkYMbtgw3Hcm07Hl1QCXYoW+6w9TdJZv
+X92GaqRWzVCYyxwcunocnkSn9UR1dYOVBnsZdGoxySMC4UZK7DLESMHcw85O6FH
aoM9kSL2jR7NHNA58c5D2zlJOPpvdaV9eW+/9FUtuGiVS5M/CPftJSZ+FO9a45ng
6wA54cNvMQcVwb7fQa7N9SGiDiZdjrJ4QAjk9AvhOyQW/ldSlqq2o6rrf4INe5ZY
5lkO7nM1VBORVy4ltcOezVnIIgtHo/OZbDF0eylHDs56StJko/5K3QgRTnfcDKgx
ek4vS9eNRJIHKVibkghNM/WH3AUVgSnI5ivrceS40t3VtWglRcq2/8JVe3/OS9sF
uID/XGys5I+wJcPsAp9yacktclhDVunTcyF5cCoc14o3oBVd/yMz14HUpHBTWPfd
ow5EnKRjSrTDvkeR+07P08BT2TzDaX+6I6u5JD5chWLAp1s8bKsOIGeHkK++PLRc
yluhNSMX3ouOxF2DAPgb/v1CZERtm4aSobnu3XiA+YEZ3+owD2Yggu44swXzcUVp
PehxTWcmM3HWxtJXLemzAR2yZ8Mj99yFU2RUl5ifhXKbs02AtD0QBoK4ZXOCuOSh
AXpnBFhub2uOpWvGHaQ3kIWuZmvNHn2MN/PKKom0ElQ4XZLjXsH+e/OsuDWNO2SQ
IWo0V3t9BTT85reXOhsl+v41hRxqjzAyeXGLY6fhycs9X5Dr2tBcwQLTOdbz9dW9
tmI8wxXPjGmh+yH6ezfWOv1uaWlTpCUfaIsHH/1aEtZjxrvqQu9t22zIQTP3evR3
JylOLU27rQMhgTQsN1NDjZonFCze/CsVRUKlUaUqr7fZPaeqWDQ26ypeQLeJjoMZ
TqokmnMDkrVrRNJna9yQFmYEk/g2y28eGa/iE5cWgoXY34X7dawglxbnM6Cum3vv
nqWyJQMixKOhKtsa4/hf6SG9IzAQ/392d5aTMCc5rCDlgxdeqeNZJGXjqM3bZiKI
w1a5rVe8bo1nDu9zH4tzUwuyC9fm+THxS/ewmkUe1TH9P+kbL8CdpToVEoIR2MOs
dffMBWCApupsN7K42a4tIeGFOcGOlHHCkSwcP1sxfanv/xQ2PQjB+80kqJv5uBQW
umrUoLjFC4shOCdI/9UhTLNMp52ScoSkw8FFINQbHn9lGPPKlTm+9ez2RpntCz9P
N8m6gIDMMTmAZbif7b5obQ9KWKdXcNPG//D7NnknK/pYs0KXOfQ+cBDyZAGGOjZY
9W0w9h5v74ATowc0LI3+8Jiz7DpGvQcU+mKqK2OtVI/Zr6zO4DnoYkgZ0CgsBYEW
ejHeqv9LKVt/FWy9i3zjfde14GIbLk/q8d7kBzWt0AxDXT2zv5olptRaVVu5LfDx
Q8I96lSlaCXg39wMgMQRA3T5B3EmMLJ6Vef2Sf6LmNIeiAHioQG0Se0UZXI1PXGP
6bxfl+PEb0QPE6nktGSEPcQeOXTNNu2Blwbm0khNcMzHoWXRyLfsZ7r8pVVE9Y9Z
XywYS4Jko13Z5fgosC8A0D/Cjvm9BA2QHyI8uA455hfeMPM74oC4NZdboDCMKw+S
AnX/ElPgDOGsWzwFiAb3fXyYk9csMzoiGRpS5/QG3xLlxGZSwWcHNunlyBsDQz83
Sb5QXG6msJISJS8rz4zszo1XLJVj7QJhGnZUvosv5Y/wbmvrO3NUZSbCxMZNbgUO
uedtN7npBwypBQKtIGLSKwj1QP9Q2ymP9EMuNPT/p6DobnWCZVUTyQVXtkNVU7Kw
fpyXHeUjBJ3X2rZrO8rm5a6msMoH7ZB2GDgnvhUouhlFJrpZw7iGWIq2tbJPt5ZE
t9WUErKCS/ZSG/3wyyg7dj+C+RDqPL5UldeOwzvp9pL/FC4eFKJqo+E4bq4lhUKq
HPeFhjSyUDp4AI4mLAmkM8s+n0SX1eBubqZ9AICGvjphXdeHQcbY06G0lkROx6Ad
buCw+4TtVcdcLhFHqT9NZNkcie3esAHv/pJymTtF9MgA1Pikjvm77JCIX/Yd4hpG
fct1lX3xWwbZ0YY8w2KXAvjQXv1brqYt/zOT1v/TApAxkNRY5LylPK0GwIdAJBHQ
va6B6pE33qn5dIOGh87BjEOEg85EFeQ0oPzMkbGWgke2q8atJLcSVguSbhcnD9qL
1G9Cx2wEYF46X5JCP2eTcRp9SJ2xuZ4KNmupXBibz/nUMYrTbSYb6usRnoCEJKG9
YX4pJ+wyzeYMcaW3kz7k6PRa1ZHrvcNxNDl3gYkePc2mhZadhz4ZO2srxMYRlYtJ
YwyDvQaEJ3TQyqoOjEuqBVIOztvxqwa8XkvspkbC3bV2uAGW21zDg8z+N4xeOwI8
QJGk1BPywf2JmlU1AVSkH0X7LOjBMQg+LzWoF5KLn6YhSFdFTVnKX3k1LXYylVIe
p4dl4DjdTsS2nnAVL2w3qJfGxcFEmKEV4y4vE84QlbA5hbhaMX1F8Cs5zJyjKDfh
39V+d8Y/OyrcHHuiwxe6eQ0tWiuUlP639L2n+mE02Vdgmdd0QRTQChp/mVqykSl/
F5u/Gu83rDXqVDGCOz/ycPgqmcV3sABYxM+tiIKtvOsHSGZ7jfiWRC/ygwK3iE6R
YM6jSppxDxXuzK+924hjlGDHCuplOFn8LzbY/blyBAUG/vY0b+J9bb/vT7rsDh3v
CMOU9O/OLxQLOrTGFVVq1PiA3oHfPdWr5NbxvfoVpy/Pw6w3nWUiXC1pyjZxnII7
3tL8yGZQMess2SIrJkzgAeff+lKS3fvA3TcU8sRWwTCBkxBvX0xh6BRKG5P0sq65
TkLYPoKiXBkUbKB8URS69nCWwOPXcVbQ5DAuM3/oX7nvow52HojFHls5hrIVXdKH
uUHeVtP0n81NfKoh1QfY1WQTDgmabNJjc34TstBVk8EMDNPlFUfWGvvtficdnB4q
dKycpXWcJyYgu9BXvLxkNjwdQFkSeHz2vsCr+EbZcFX1e9i14BcWwx+v2sYebKHd
olZI5pzF//eb74flh7veIBvHpWSYHY8/HA8lIBqJBdysUq1QMH49XSocjqSC/xYI
E6i4S1yBF79Ke6plGzCoizK5AQH9dxbEHiYORLT7fINbVmxsTKGN67DxyB2CJV9o
qGuKgeeUmvWQO26W9xo6sy6J5TNu6fNAKxX79UWo43Zysu+rBOhhroGZGjHZswfo
BeQhZVnnEv8e5wGbfOG/Ytdapdygvsz1YUuIZKucWDu6im8R3uEtb/GpcNiyQW8h
m/7Bup8YEVYl2RS88YoFKDJpGP9OeFHLWed4eyo8iyzuoIdcK3ekj+oMvlggIu7A
+nSW7fMrMmDIZ94FcAGqt71k7tJVhf7mGHnIkx1GTY26bC8o64Zpz8x7CpXDo6HX
0qiCQT7N3C4Of2WyNOut04tGmchqCOv6Xevy06lWtsLBkwiKE+F4gS4qrn6kD3Vx
D4Y/bJ6f9my5n0d9M/tohEuwMJZ9uQe8x4kxhdsxRRCIld9wEFsx9ZvQmOoAh6oC
VUWE4KybtRquNw+Vrum0cYVbzhSvKb8LvFG6PymXp3tK+/CPjGFjrGqCLEv2VEXO
QNnr/3AzJhJ4b94khkbDu2xzvcMFgvCes3KhCNXvflj3phL4769pZI0dRUDJQdK/
0v7mAXwQIsagx6fWZGbhzsh/0E4hi6uhO8yDXdp746aLUZQcCl2wFH0aY2szA00Q
Y/3hOkVtlMMlUd21mamhCaKc8zM+g4oyTWaSdaZQO4mtl+3o8w4pr6jWVnbiSQyW
uri7/5CBUYg007mnbUyK/NyDaiBBZExWAfO7o6qhrcOQDfXli4JKqUHEKxpn96XL
6AsUqh1OA8I684vZgerjkmPrPN3c4y03UawIuLNEOcYmdd0yLGR4fuz0VfFHeonf
NkcSNqTzEvh6OP2R30gL0ebhXyJLZ30ciXk7F5Mo9N3IhHysbOxwjOkUKZ+zS1s7
NQt1/vB0Ny4ru35FknAOZlbXCjLF0SCt5JZp62w32kGtu4k4SIctVp84YYHqN5ga
t7xiyT9gs95HdJmUmeWxxAwRnJ2vO7iK4vpwdRsJ1ILQKZIuroVWtoH7oBM7VTw+
7M7aSr5As9SyHhvjbdHqWBpjUraYP3S6wF+bP0ALNGwelBnXpMVqdz+gXFbYMK77
qfiDTY4W+mI5EPKWUu2BgEqQv7m/0GoyeE/y9epW4GDLRlHHx42fhF1CV1+Zmwep
CfdUdwTKU63hE1eC/vbyZJNUt7roTvWoQMgPGD3CgMruhgGgAzRbVCVI1DysQHAz
zn1lc365P9o702kEhWNpAVw7YOv0YlepsQJtWxDk7s3JfWxV40YU5GtazSVHgcNF
yrTqsZi84NKXWZ6xHXv6ccRAv+rDHT9aKmwWiyifCf3/DtMYGVXtgFrxbnxREP2w
ppzAnA9V2ZvCl/azGyu9dwxbkkalluOkllEJhm9xH/SiiOKa6usxAlxi2dGOGxxB
LvR7opvIOp+PLVxE/AACVQ9fmjxFFzuiaSt6oxCszX4MsB3YpF/lE8mtVvbz7L5W
q9W+NpSGM8X/MuhDKotCVrfirSnAssv7bWxEB1GMvOMN+wreVwrGXuo2MGpM1Iiq
MORzAnxl9SrS+AJhKWFKmf9W/qL0htii6lKoeTklB0XdXB5Fl+Xuc/Jot/mYaWfo
Ay7b7be7AfP0eXuk92ZjjmG4qofsUjmtk0My3Xlp7q3ERz/u0eqMWnfuGvEGFqkq
QqZ6/hcyHjfC5bBgVeWxR9ylQDCGR7C+rHh3FIhAc6qvEHgzZTj9gGyPt6ArcJHs
uS57LaofG0Xv7ujOx0Da2Qr3MUa7wYOgAFlYKQG7DpoBLbHxPm055Qnl0JgJGCS7
H9hYh2ROdS+pqYDHZMNloeiHdwDYPN7oETj3HdxgwkBvlQzt7xZKY+FGzWUIEQwP
hEYhX0FyyvZGlI9Lz1fyoa8Q3ijKvEsHwQ/mImCRCm7a69WOfmZG/VQ98RigH6nb
ihMWv5w/hVXA/k2eT7qIqGRrJ3Y+qEWDxEfzSrGbzpHsHWjHIVOk8wbH56inFc+0
ULvpuLVhn9WYd5BXFL8R9RuoGaUtFTxtGMrFk9lhK9zvU6pix5PtbtJKOTk+STFg
qecHxF68+GloBIldwHhRleqQ1TF4HXHjGsR6PrbjlvMk0ovik56XejFqJv/Z98Fy
5N5lNUbvqdydBir3xXG1dV1hAw06P8+GSgW+V0uA46uw2Cw07TguWEdhZCz1UaCb
n+6zYkAo+IGgvLFLmYu0Tjb7pryDdQAhMwUCxxqVhQ2PaGCdal6LQPK6jlileygG
Een09v6yS4LkFssCRWOuic+X2asjNRvmhyXdFcFfPfuBwR1Af6Et5NOz7qMYLywu
zlwpa2zwlU8TAufCpNCrK8k8zwtgHwQw1ugSAfNnsa+5BB0bscgQj51+HFVg1IQO
P8LsjEe8nBrFOZv2ma2qZBrJVBQk1OMoE8bYMfRXGOPJbW6zWe5iGSyiyclYPTJL
pqusWXCmnuNnb7Qvgg4j/lz3/IOL2DMoA+lPkRDRYJZjc9+jCxcNA5g7j0CW86WA
RBCbqJC2MVDxY8AApSrAFSYDP8RJcXD8HsSvmRiC6wXj208YEQtdgUWrZe6WeCvJ
oveNRSXFu4CrlDvtJsRChB+dW1Vfa1ZA+Nlfz3H+7/NWz0ZSFikB8ZtfAM2L/cwx
qRAOflWA7oI+uG2OmOluSU7PMRHh3BNkp6XuU4RzQwFCAdueeK1T4/5qnuO1mxk1
QfZ9rDY6O7xxscFKXsR+oTCJeKcmJgbN3a7moe2I3lqxXYLCyVKxkpa+DSd+Ffen
5jNEysNScuBy00Vbox1XgtXriYS9+o8IjQOrSRQD9LaO/dMe9uGgn63QE7zvI9kb
dizC63pgYIeXfMqI8CpwJARoW4930bqLW1sZKSvblT4aKgJafkmAw1M7hSqiwNeT
U1QqnefJ6IY11qDujnrpF1pCNiCHVq41/xN8KRiWXWwzZMPxY8eEKW/vRW1M5ePe
6PypEM5YwevSz21FLUETBSWjGYtH0ZYislr9+aX1kZlf6N7Vp87QwWGCz0CJL3NW
SjEY5PoMZVyz7oRi9wmLHRGkmxH8kyf5ElcOwLj3juUmgfyBLzmmPErIH/rD6CDE
ulj2Lxrsu2HFhm+ys/Bj9ywWi6kFfhZcxBzU4FQYhekez4CyY4vQe2VUmaoDMPex
07AUrQCvJz7idx36sWBlpSNOVpRQo2a5MrZC3TGLj0UdNwy+syXLDwbjKZ7hdY6X
`pragma protect end_protected
