// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mqP83fmVXaW2rqlJy+1S/vV81RjrVeJiXjMcmCI3aK2zwx1Grex02iyKKMsN/aTp
w6GNeqmkG6Sgslf2l1ANh7rO3VC1YdfnLqaGRqvOo4Ip62KJ0uFUSp67YwghQ6gc
26TgKEOrm3p8d3pUFytCy2z3eF2VIfj2OlcB0hprmm4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8128)
g+iR8YfKSQT0I3SZeGU2b0naxgVfU6v6rsNhE3HvZc1ranMipNf+G1FyrQdCnQDU
a31wuanWPl0y++fN3SODvVZ63XVcdljHRcO3mb7lqDMYdeKTuLzLiLPTm1hOioS5
W7jAStv0LpT3wc9IjmWyvdivWhFvQbdXcJVSQU2WCy/vaRhsxzriQ7P73Ir4Ye+M
ytETrjWX5S6ZqFQsIgjUgI28tv9POEHdwD9DmuHnq9nsHcGXjtVlSPcFuacF9F1C
4YDv2pECSGgnBJdZWggxcO+tq8wvL0tEltTEyM6yiRrwRxKU7SE5r+U8W8Es6pUz
gKMiXqk1d3aGuW5QwlkVZZ3lo0gwTKjw6eA2QVZivi2oceWXNU7nP3Ub6+CpaVZs
msZyuVUfTJ7wCoOGXqgCkv3CCYLbnN8Mfvs/jV7awR35heqb5KzNq53z3LrCvP/y
b9+2fn4GjodCOCJpBAQehY7VqBxZAb4VGUYCJmqO3kwu7QHTAHvAMAGtvmcPsVgG
Qz+h6pkH52skSOc1Wf7SXU5fRuvAJOEfZ8UVkCnp2YNg2rbQgUxqCOTDE1fShtau
6HTcpO+p78wV2/aQkTpioWzrHTWH9wp9D1nTsqbpqfiG/CO8d2EQJdDhD2Bz5ORz
9Vstjil1DKbFrOHIqSkMyh0HgFZaHm1ho43CF4EdZTxgDsniEp87LdgAM/+lH12i
1rKNSDLPlupiyxddIei8QJl+mO/qGkBpsaQGtw4ueuI7wy5pqVORAm2PI6MwFrU8
JUCuSsuywiB8eAgC/9O9X5uNyreDOZK5+Z6GE1buJQTU8rc1x7gqgEW9Qbd607Vi
n+iFY5sZx149joRD92QR+khqe2s0+uwG5K2EILiI0V3YsHqGYgzqzljzMawDpTli
uiD6OM30XMSKACJanHVhcHI3TojIyCHqtJfqz6xctEq0vPKnB79lqH1PQpXXp1Ys
SewQNr5j9WQs763MioAtERoX9+bY9ysKF7xGA7rSHOQ9PHnlyBMjFimXDIswfJyP
/CCfx/VTJfbMBPyIrk+rPqmCcy7fN86/OKWqCk0YVNLKh2vfLXPFlR2MeeVltCPS
gGPyTmbCoM8PzwMu77N4I+czZTPaCHQ3Tap5fYEcAQQA1iQQBGTqJk4Gjg9s1pGg
2YG3ncTqB8Wg0TF/hPniu3SWTuaqx6iZtwktLPHNZwZwcUZ963MPQhObnfwa8JEb
Qu7hpc72o+mF9mGrX6nKpnqcH6qL1lhyHspNaucwKebI1dyFbwlROzShObX1GmRv
ablkGNmEw8av9vR/xV1ThnEbpQYErWJ9INYpT/45di0dq3dXIQytPlXpDrhmphiv
76O/J7zwaXTGoAF6NzyZupKrts+qj3nGpfPP5KeRh1sLObD/+06f6N7OIV1e3wIV
laxn9IUwvbRC50pgc/FqV5PDwaspZys0rbF6z25UEbUZBMflyN+rEpfnzbaVt7WK
Ao1YzqmU1LiHhGzAfZKvyRaH0dRufKrIkNwueMBSbXQCTWHflPsD3rjUf3Dc9jZV
mfW6JpcVoaZ5Z4WNFp98iK/uXa1Km1E/Lz0zMkB8dld7zyXAyn3jxZCEdnPyRhvs
F3frm8mrs4FNVY16AdCS5NpuNkD76t3gVzXCehK+CQlYgPCWfW/2ZFv1lHMVc0s+
0ecSrIkXFgAXbZxNu75f7tLLWVijZjgpIlSNRHO3Ddafv1yml0B4/nYrD9wvH8sH
niT2MI5mqpc1+F/+rZLDz0OofO5zJ225MkJvquLtBxqj9N5d82zkmLxpFei/yeKO
zGubIo8E2HxTp7DEkXmc27RnYU34UZMqTKfhlu4k8kdvcV5mUHVtRMC17ortmGJn
HF5r27RXzqA3RrK/UsTcGKgV5FvuGM5HS5KgGeEqlJak3jFHnWB4djgDI99cVIG2
PjWXowMN/Bft/gZ85VgeZNs49LR1Ier2U4mJsdEBvCo2vIoPqtOcEl5XkTFGyE16
gAXDiulCrPbLSK2LdOzWNml4C3jU+F5bT/YMAqDHnw3ecA+WsplwrIPuE9sgtu6y
CgMNLbDVrrGexiJb1eaypHz2hxYh2+sn7NgaS27gtY7ZljQayJRUzd8QsTre4Q8X
nV8+trSW0lq5k4/W4TqT/NH+9orV7eDbk6V3EKF2BRzI4Ut+24qbq2/0zsJrt9Ex
H6w3+P6GTAMPc7ocrNRfG+dllLWC36LXaTP0vItzNK1pEDmGBMTU2/mqV83EIRP0
Di7rFdyP/2TZRFRmkt7Hhw2PpSOUSrtfgS7E7uYefKO3IAyygCFc4w5PLHJhLdNI
lKUnr6cwvjdHDqIKt+0HvprkTUjzMIgyHPasPb+IVH5vfxy5o1Gd7nE4S+s1KlcT
xP6i+tmtZVpmUJ8/0dvXLr1FFVbvWsbn76GAZoFgZOvOjiJzyfzybeyDzoDjZWFn
1efQ04A6zDxJI17MqfA7wJ4LPZwuDMnFXJAQM3vQ2sSPBDUqy+qMOEtfPMn6hDQg
srJguI9rF5+HgERr1wyi9GIly8rhXIhLtZePEtX3HLVVleNFo3u8punc6FfsjGR0
D6xGO53SeVQ7elb/av+TZPvUpmgZN8jug/XsEy/zUXEoYNqKU96Z/Xs+gMtMIsSc
oW5W6GKyy75XJiPAkISnJAoFHKPO8l3pk+4AvGetYwDpywxl6K/Y8iVnVHl1/ndY
oKpVEwJmkDG+/41P07tm0B1/SsRBiD10oDKLWmP+uiSh03PGN0MVKi3AXRPcN2j/
uwrWrSx7egfcjMDkmDTpxk5aiNMceNNys/WJ5jt5LvC99o3tTsLiBeZE2aL7pfFn
atDGFhdRELZRc/rPu/FDN5J/1SRHCFEWAWcrpJmMiBo+C7o9E0HltJki82/WE8Yb
ERsk9/y54CWmmB5CxSEtiQa70ERlXZ5OiIb6ttOZ8P9qZruY9UfogYCDL+sukYXV
Lfksgft0Kyczbn6Wa5P0ldayqhnVwZHQwEwIzy+4erXRau88ecvwF4NFL/yHMJ6h
m9lXlAivXwxp5sAK08FlaxrZnUeLtNcSnnCrd5ahcHj3hzQiAzWOzy0+pdG1FEjS
N87AWQiSCUc0FPQOJTibItOQ0lNsf7O9t43VB4tXa+AR44JsQkW9LRX2BlRHHxAr
VaZnveel4nC0wojCZRA9V//5mXfUEMdYZR7rFr7ot/oIl+tc4kyn6O2pMMqa/y4o
st+nZYaW+k4wlqljB8hqZI+fTYZ7bud72/vhFw8q1QV11pbZtgOL8xeEBU95HpoX
OFwdletms3kfLpzTOeK3vDm576q0408A9wPoIaQAeOFE12UHY1cY+iSG88sx4QUp
8qaxysdbBKY0XBeyCyN+wAvNRhlloij3wAxejjfQHI49kDzKusxgz8q4ddzGAEH2
90svg8csyRooItTZRXaQAoWe2hJQ/7eVcqW/6MAy6ZlVxDoi25CJB8h0YBj+vC8a
qLZ1ef1Fv/P7cyjJXkNnpM8Ec1wxZV1SAU2dzivXfZH2aVoOABkECyveH5ov/zq8
NueNb+CU7Ni/gcxpBATqZCri2l7b+2kx7NVZJVtqwxXOrcNjTof+cYu8EzWLKcpG
NOw5JFTB3ABSrvuCpcBGf70b1yGtNIbb06gHUleqwO923dG5RM0rmBm4ADmS/O3s
H7CV6SBWyMGD7a8GjpGq4qi8QslAQKZwLQHrnFHv3c9qEkw8zuaT6JhdgOO+1ksv
ioW23zHZDpAFoCI8Ifw3FPKcXjT+5M38HomsjRmwSynWZV1HgWcM6MoOX5lSicQf
t7P1UlJjmgICGEloEMtNbtaBOYffqdzWWoTpuSQOQ7k8alAHqGLVw4ixY8RZ52wn
CTQefkzdjCWojsEpmXy9dZToKu2dn+AYscLTeLnRt4dH+A8NevlxzKgTlHZLBpoa
p4dLOu9s46FIbF176wHB8xyv3Ry4Lb6Fv+ErByTFaOqBQorzmS/R1HPAbYN2o5ma
c8yyRWVZ7bbX2Yxhgt0C9mELCf5bs+bNSSJBmNl/A3qFcVTnR71CErwhfWX7ljIY
pMGffjSO/TUaneU2pPW4XKqrrHOD3VaR4a8NR9cebs9B89b5tt1uLLkCGBsUvYJs
MhQHD7O2a54DtHozd7NqWob7U+Oj9rJZbhyuN6FAhTmpemUeuda6qqtBsiJkcF2w
bAq4k8llaO6DygTgVPqPWJMope2ckGzuAoGXuOLq7Jr25yjVZLdvUJPuYl2q8aHJ
qZiiDcMiAzMmkG71OQFEDFCcYPwz5weGsU0cPZLOZ3Azhts0jtx9O5j+vJv1jVOI
bCNm/NM+47+do5w5Sx60ewuJW+nCP07MAElv5W1NYRTmZxBc1vJ1kNE/FtHnF0TG
RCJDtyh6iT3L9ThXoxsCIhxAJIhPGUiPT+vW1USPvJc9ZiNf84yvwkcgPmxxaLY3
CmgTcyE0/zfrkVk5voA2jWDVqnYbEuavL7ABc3X3kEEI71APUpe7R//ToauKTZw1
EczesHGHoReMONvCcxBvoJSqfrzzdPZZUevzimwVjFIfjwlbl6jLDRCJapSVzePk
67/eVsfu6VxGzXpGMZ+cMc5Z+NIo+oVlTkNioHxJxbM2IFAZYWZv47NGZ/Nisor9
EFwDEPIufm9ZhCPTmFkLZI3Ww6dslRA0MRgjGED5gCOG4DtX188B85VHmqHW/M30
tp2OwzrUpWBE7u4T8zQnBM1zCV4MSzytj+SqAgHCuAwF+la/Wz+BWjsmIahINM29
13+F/eVDfQnju8ZVH4qXw6VMwO+ReUIyGpkZ2GPqzGMeY6FGmHy3ljD+xQcAe8yL
oSvlGxPolRizg3DzWdvxG+Me86o2wTzoqwbUivAEMlAiZ/H9HXOkQzw2FbbA6gAw
YjEBgxsNL0xdo6FCu6xjYcl30nqdL308ZdsO4iEIxqndDo6Cumdtj+/jaD/i+KYW
I8pXSK6JBGEGXMnLufbfUJNnum2oslRrCQRuN1P/o4e2vUdRyGv6LZq3EXLdm0LR
riHk2SJZeHfQVnOXBi72beW+F9CK6a0INl+1KTtoGokB1FL1Z4CTN3tq8sFjRzqQ
kW3ThASg1NBOUKjHJwp1AjjGkLNbPnO538nM/AyY46OqfNyeppHFnwwv0bJTkf8i
58RSf6/LQINfXiBYHT4aMljSzoAmP/B9Kyt9mqdwfpd2HK67VB0mrsCzfnLLKuyH
Vwo3vM6cRPfBjKxv5N1bmhjaJK4HDWSZ/ILccK9yxke8QOy4f9e34bP0MNiVuzjt
7uMx1/vCiUWrd/3KC7SRWd5awxgzIZPVJfIBdiLEh6QGT91bnItrJKUnPXGd8Ejg
vgn/0OFfXHfY52GZy/HfR+xlI0XMrYlkMYadr8w2rzu+kume2ng5VSX+ISRdl6Ev
PjmtqXr8njRbthD8xKD+MbNCyOoY42LamDdEICxypP3xLoPaR/lGvky5HaBOBwCM
SVjwqfFIHogYxl3E6OnbT96vdY2/HbA6ynnynOpfPR2Y5dJUxqgg0VjjzqWRM8dd
sTGtSB3WAUqeF2VCFi+r6UC3uq6GuTy79bdubB8rixv8SYTTccl4IRzQMcmUNCPH
LdCzPgSi3/dhbUQJWvpcwkKMJk6Kcayb6eNK9NLxfBeMJ3RitqVGnnVtDHboXw6t
Qp2UJiC/Ft36dhNQFQVPE+36CrMpk/fv1XQ5+DuP6/5giAzYiycp/4vTR0LBC976
P56Wgw5TUZnUoQYjaezo6n77rDCAWiFsSNNeG913+0JoyaZ99/ogtk4AfLitxHnd
R3ekk4O9PPwZdrNk+y212xRNyPQE+ez1PBnYm56mHtH436nson+hzWiXyXORC6BN
j/EMCQMaTEtBQAsET7O3x8jRtXWfJAAEb7KAy9j2lWzTwfaP/plkYyTn+pt6srU8
VxG4rQJTK+OMjPZ9y360pmHEIVSVeaQoYHP5BHhPdab9CrOOaJPFQK122NFPourd
1Q80b9zZiPb1iQ6N4Mh9dhmeSB7b1rZSkoVkfaLb4K28/3mewBU5FZJzslHIzlD+
VhWr6o4c/bnXzfCBbZiBfbmPD7o3ps/clyr03x7nLjjEZPoL0BKpgxH8gcK+Q6g+
367GaBUFgsSUCNmElO5QDcZee+5dckq6k3mDxpwmfFqzQU+TYoBOMKPqtTcrq6o8
IdIomT4rHOlg0NWU17E/eLsqO9yTBOhiXBSVUbez3j5C1GvuaR6BEHIXMqlVBrTW
cU8CPhRr/cFq8AtsTGDCGA49+I3mdPrqOUDvb+czrW9kaGAk2ROekcx1tT3hOawE
H5RSfTDl59Qi4HbTUq/9l3uK/qBs1USXn/55vj6dzIGAKKfxUPEC8nstNTOwVVUV
WNVvj6949ZvTuUOR4jRISx4l25rLuzL48MTMhWEhnWVBg9enIdwl+VWlIU8px9lt
SLHEZXw8uv41/a2THAFDPh7RbjP+jISAGaDnlegxMAHYRFMS9nsAR+qOAuKuBL2u
WdvZH4u5QiuGHg/scCJRhiw40Ww2nVPV7um40eMQkWJxfsm/yVYWStu55IpW8u92
MbpnT9cibCc6sYIl9iLpWcjpeOmJhpwDFVsZVv0wADw6peUY9eVtyfQ85JqCJQax
tPS8/7c42XyU6jF1aeeGyQFHLZat6dNzIUx/04wg8pXk2jB1tzXwM2WdmA+pnTGC
HiZdED+KcDnHrcU1rqO2fu3nJLNiu6saPlwfJC8rLFrBzYK7f5GP2Nf1qo6WMKB/
ltU4BhdCYKbfSbU0vbwrLj32yITIlGWifZ+aViQBaUzX0pSd/ta/4B5uQ6WcKDB3
ep/OjBRpuirLSbJrMKrXoULpEQgWezXeBQR7JQSiBSGwyZI1HsviPQcRdA6WXpH6
eT6B3/Zs7+fQW6p8XyTeplBbEiljYmpP/m1j5KFeTrh1tQXfnpIXZ7cPB/4EP927
IH53RqC/oRKqnwi53wrdTR4iFCVorpwe65dc/ssq+Vv8Y81wpsaoSlAu9bvP2DkV
tH2LwsjLTqKJ0pl8IAObeyHbD8th/7PB+/RoTegb74FqP8DFprJwf2nVb/b2mBq+
lEq7hh5PUPUsCOED42Ch3I9Nb3UHNAcwEu00WwyMoL3/n04/vYpsYnT6mZfHuZGQ
hrjU3wwQjfBVpJTpzdK91eRLh5SQRpjq3HVZiP64uNXnXucVJm/Zibb05JXw4+VC
XBlKvHvXs4Go8vtKfI5DhYiTsLKdCgsqGmMtE3aLq0RBHbakHRdfGSWb1kjaVBOH
Wb7KHLed1nZtGLg7o4Prqkq5m8U+vtZNReVwTEWjDb29TbY/2DoN/+qq+ajcBbZ1
LimxLOF5WGYDkm2DXwmuLEyAa2BH2PilWdcNFt4Vz2vh/EfNwrvGvWW83jGJ+0ub
S1f3dfVVrbDY2p4muHcODtWmSVioz8DGC0n5hZrbDeCjTCFLWhalo4NcaX8MN/1d
MB/xFGmTR7J0HvrpTNPb4Sj0PHlzcWvus76bqAUGYhW2j9OnBkzMBZgcT7v9lBcY
cmQeJJy+haww53isCCU6IDDWs0y57Mc4JwFYMVMr5c1p4l0gynPPOvaKs2b+OZ2L
GTzPEv+V+vbt1C+qBkFGrO+KN6m8NjP7Gq8ICEOvSLs3+NklF9lJH6FXJ35ycjco
QKCgrxYnIrrcLoa64B9EzhBYe7Gq9VyfVfMiYBJnyfEhrzwzoa35amGkd1fDHxoB
KmjY+z4KNFTdSXlYDEOQT3Zr8AMhGoOSV49gANTme167laNohy94f7kOzSumowFF
wyxIg0+NJI2cCg85ECdeZCYT/XT84WLxZMSggUbYEp/XpnXfBP4mmw/iCH6oIBQr
39K7E/MUjNU2ejj9ryXt/kak495l97cguv2X8ik6ebRA8O0Lim29o4cXDy2Tg5YT
VYw6tdh9gm3x2XH4fOoLDRbhVmKEzd0VU0QHVrIvZjRXHMPS/UnpksZKVwsXm4YQ
DhxgkrqS/um/s+iOvgsPeZrL4gsX54CUSqhWP8wcqUSqPOAQCFcTAmuIEKKBnf5s
FRc/srktoh8YPIyr+6nrRWkhtm96L1rPNsaNE3ANrHnX6fLQD/BVZ27UmK4OQVgu
EFSsfEmlj546cuL5v6Kbwufc0facM1bniCX20JaM6PMoB39Uq9roc/9vvqTzL4m2
J39I/me8ywp18+cuGITjXaIlR49sR4HbUugIG03cahQCTajXodf48Oll1j8AQq63
uSXG9WgCwwmx26r01HWEzLUNx3F1guIU/S2BR4xplvCKM1mLAqJdbqoENejq+mAB
Ls+DjOIKr3HD5NT8O8eXcfVN+wMwIjv7IpMn2tcFMgLq12L3ZCLxiVkCQW/5ok0p
QeTX0+fRVASAvaX581qav5ZBEs8VcDJC5EiJglG5wl0W+Rnpwg4i4/KMoOCMTUY2
/bJLfWbsVyYrtd8rymYnBbgiqrf2E3CAmdYwGulkvFyRho84vroTuMYXADIndn5i
w4PF/jomer/FIPTkrVC2vgKW6y/Osg2JFmLM+xYjOqKagpYzLlTK4kWXnzlIi0uD
XNYtqi0wbKjOIqL27e9hQfrEJVpZ+3DpYPb30IY/LhGZsD+hlnByHH1AO30i+Ba8
OUXAlrnnQ26gWHO7Ea43FFB7yHlotxme6pd99dnC0SvzLAs8FYegSUhMIeTG+E65
tSe9HKQCF/f0Ru/g98+ICkSOczH8r+lT3pjj3R8+hyPurqyklO5pNdtRIADQJhLh
gXwljAOQcvN4g/lg8+Y/jhrJsTpM916wnyjU+03ePhwkDt6E4wCYfBiniaDxLWfx
pqd7P/kVcgxR4tPvSX+9m1Xeu6X3TVp4NKHtQVvyOZFC/CM6/uP3Fz0Nhianlp0z
76YejfRTy9Sk8qntZb5zqlITEq6qIuxIzCUCZSgfAIOiKxv1D+p4PzdCRD9RYzv6
HpNvH5H+/yMxzWYh7o4bgohQ+U1TwqBfPhyY1XoUv1mYxQ79LZWlY0ZEFaull/TU
k4pcMnTiUKFCcbRIaikQM6vYLC+kLjEOHM7Nrtelp8TP9huayeAryfZmDrjRJ9IP
rEVbIfwZzVuqoDHHj0h3R3DqvyLdKJ2Uu5yYAP94odlF8lBEeS9IcJWp+er6DOcY
LIv+1gvtsucuxDfbyzs2K77QROMtwR4MLnw425YVnhSYwIPn2JFUxVmm6uoAbCMj
8zXH5glIzj44+eaKkOYHxx1WWl2gQCVMHsVQTYYEw1gFHIctcj8y3PGB+mdgAwK1
uBFEyaaz+Z9GT4QKSzIF39vrs5CjwJ1gbqgSFaTImNKSg/Kmlo7Y4fCQhlTrAkYs
yKO5WCEprv5n1Wch2DkgoFMDSE5gzs1XCD4mHMXIEmDPT1LttLeXodtCni9YUDaS
PsOxftVlgmrrIVzG/o4+RWejkVWaBL4K1bTYEOGwi2pUQ5Z7KE3dvQBv9WbhTwaq
qXA8xvW2wWzDgD8vimu4l0RAkAkWyFRXjcO1BCcRbkZcpismwBI+XLwj9zHFS344
l7y205v3jy3B0ZLKtwABlXUPUrC7Dg/jCcgYz16Luv5BafKpsY4yF/RhAzNkSL3+
5aGiFQrglQVO95Y5Nk4hODIAKyfYeZIoqGW0EbFwlDGwTzGHRsvHTSF3fC49J2LV
N1X8Iga5OsbW+RTlg8Pw82RU1pCvtbYpJiU+gmpLvA2SAoHLc0x8Vb/jScEFdc6s
Yoa5OTDCLvxY+z5kUst5hqfdDVK7X+gq++s0l/PpDMBlOM1UF+4fOmFwHufzANQ6
FO0pd76XNcmiFmAEr11/wOvo1VElgifBXjKr5JwaptFZHt1Th/CnFjkPl62pWxJh
M5BS3sOPr5Ve82MOtYN1rMdmIe+i2plPAzGjkYLe2MQ6fHBOlxNx41F+/zL+sFbm
dJNkjDXFiCZS5wzeNlyRKNLgeg60LV6vrltNamS6jNdM3oJUkyI96s5m1HPRpqj+
42KhK2ERvuGdyPl9aumxIK0ezIdHQGvg0GFhxwjkZg5g4AP14YfaIfOBaMsCCi4l
ce/o7358brOdR/NgYd+ezpscEZOs65fTY6SJyE6KFJD7ANTAHhZhRo9KT340dK5C
vm6y2zopFWUIr9t1GASS7vsu5qfmlaklq+hqqJq7ozRgKO4ZuOpLU52IFNdS4Utr
pyRCO8JQDtfiowplTlnx4zOpLUEC1wpg31dKVui27n38Mfmirie3RWE1lY4a7L+c
Qa/ykUh5XVO9p7u8iLHjzsw7bIKDrf9cmGfpZgYoC7oiV4nirBv/XVA4vrTniyWK
LMwvpB2JHG6Di8HrJKC8D7KymZ7ImpI9D1+mmEwsraXxEEHgykxtCB21FsNeATrG
goSeJlU+16UNVWl/yDOmDioYU1vAdXthgRnaViSovHqwRw1DrtWclfBMN8L4FXTF
5o8asW0bL6WpsrrWtn3CWM0O8bP3s8pvGxSbvyPpxUuzn5yJr1QEoUpSOz+UXzhN
ljgz9NX1pB0/8sKbs+ft8hzAeboOwoKQMeia5bblUZN+1UTdmgjfp/kt4e/9MF0S
mglJueIBnSK08AbgWzEwlj8xchLutVJd8xf85isCoHPOA0NPHLWohA8adcVuK9Mk
5u7uWtyRqJ73Cm17drNhrEalEdeMyYrGCgEWXgS1MxePP4xwj/WXlqjJeEJ2OUdj
/uyUKrfJsBjOCjL31ApptWDrnk7h0YiGCfEktnS6aagLqvPz6IprLIWGVnwlkcjK
GuDht+eOYrTeWYAlDcmqH6w9j5vwLUG14wRzPph9Lm5opr478PVMIK4U1V460fBK
qUZGjtC6KKj6rtPouQTYeIYd/YCjeNQnL4M1jd40nBrJg2SDv4d+/jB7mG8hbrO0
e6weFC1Kyi+2lGyE5eLAxg==
`pragma protect end_protected
