// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F53Xy/ZQR7xTjHODWgsTgNt/EnveMs6GLKJhbjJY5RT/6hneNg1bmO2mJaf1Bfje
7qccJWkMDMsDtX2QX16z2q0zJK6x52P15J8Ftw2tt1OGTQZKo7dOzUlhH1/4rLfU
08VSGHLgX0QR4idjwBIVixFWdRFNNC2eNrT/aPrJPZY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28208)
ejmrWr+4hdB/YKqUwS9tv15pBXQaQqR9CD8gjlrXf6twNHLle4/Q2Q6xQX6ybEY+
G/ODPZlu34HUoKl1IEeiIRNR7jsIy0xR0L5Q/kZFieT5TxAnR2jI5gNxF0Sj3Eb8
vq2k9JQU6VE2xNUMM2u6uFKMSHItRSRR7d6fRiLKh9F8QjD+1Dn4ZZhOQFsHtREb
8VckQiNrgqVwPAuEVLVu5HbhyF2K12EIe74Ogm1nXQb9TmQwyM1uOMk22HhMhYrz
YDvW+jKO3Fxd4ke4t2udIMtMdk9c/rh62aBOVPMBuTUBEdt6mIumlSeFj8jEmupo
ceZRHaRB1DXAP9fX+udhjN0RRmnZhI+Rfl81vXlrxdVFs6+zafpiId7siShEBEaw
4fxp4jii4+6tNq2F+JUKJ3KRA63KHFXdikPaCM0N8zZTbLxwAnQmgudS+1psTVOv
7eb1NqpkW+ZsH7SFgFgC5c5apUkatL0AKtezV3Xrj+tSEYV2j7b+r35v8UhR9W9P
9PMmXShijZYU5nhYeUbqCl4lNYrFt1WYBmb/yRxHTTz03e0QrSu5URkAtnHn6+od
apoC0PH7s0dfnj7zpC1tn+cAQkyprw5BQgaDoahFJXQZ8CYLrLLvCF0T8cuvvuo9
O0SwVJWnjmG/H6+1dMjXdLQAedDn/3Wc4Vc0LRHQnfoAhauiVolU8uyVj7sqjozJ
LOT+7kgaD6LJ8U0FKjnAV6Opg5TcRBoIkgjp9SbuHO+MNHgJXdhxHUy6L6pKxk2h
kbIMkRG0jTNHzzh2uoTJXL5jwMpKYscY8U1h4BTMC3MopYbBIxFnl7ghbieQoWzC
2CMI0YPYQRVpOz3uJWbgxiMUU2BGIIo1vQRc6NperXwPLZ+JYoUm4HdILDTkv5Lq
lBt1Vq33VFQLRKet/NCeLp506+n0jCIX+k/yhfbDCon4B85blWnERItxJXo2U8WZ
WZojlAySaEEIxNwqj0NhN6r7IPEh/gB4cmujW1daM+MGu8Q48+4jlJ0wbDPy4Kkx
iK6vn/c/EhqEiGNfJHrtAgKR3VgLMf3/xYCxj/nwSrpMTOucOvo7ZUMvlPfIW66s
FDEXxzuLTQKmhVGiyqS/J0kIEwlfT8iNAsGXpCqfopqg2LD3V3wtHSqA3lrHWLT9
lWzn2EH5nAouxmSD78lzLwSfUnQLhuDQPUGovGcxR9Kq93VF8N/S05j94GpGqSAj
TTUD7RVctlpGHZi3Ojwm73Ra47hedWmuV4deqaE3d4WKf9zNLbk/FbyxCHhgAhyT
5k4Hr4rKmkbZYIJoXz8h1TrTkqeCQ8qGuygzr/xkmjAA9NHMtQjETCBpR5irhyyu
r3cHHZJTOgrn3vFH4ial/jBsAy1YRrZWGJo7+lfdJubqi8hAMZIT+hXFiKeH/2We
OF7Hu8Zw6Ux8d+zAoJCFZgAjrUgn8CSQgoMUCj8Eq/FyvcSXOANEabMoqFerNWpQ
DzB/ParCY3lN68uk474n3lkeIQvGkp4zQZJHXJv//42s/TNZzCKsx4nDz/stiegc
m6Xkw1uGZZ8vjv8XZ4XsHCa+fU126t5i21nwafIjctBCZBPm3UmNd25ylK3R1Yfe
P8ahpr9FxfG2xYoCoN6lLMC71loZM+VVMsPDEb6JG6MZfHiONzT+bNIkKUOpLi4i
3atYw2FHq8L7IVrt3MCbhfj7THGahKfSjX4BBx8Ua5pPpu4u2+6oUXsDJY3KLhR/
rhzc/8cSKqrvwi5WcGBY0Oe/Zp3ovHpA2u0xNlIchazPLCQ2Xmd0s7jysTpCteMk
wgmInLzWDjqzL325smN7ibyQGPViXF3JfaT3ywHUfcsCcbMxfZ9s6Thpms9uq3OI
cWq8/FLBXu6v/xa3+iBNr2cLeSBdxl1tyETTEbDRO5hUU+7u1xOVDXJTi4+qjsS0
Qr7gWLr9iVB8b7wk5oYFMrj6HBfxetKjx0rgRXnUjdepf5nHq/xXR2cgBkuhc6H0
cGssB3eHEwyJFDif3Hf07xkKKEnyu5pcg0zuE3QNGK9heHjxTaOf0o8vaPmeS/SR
B7+6YbBCnN/Jr4KYSwcPu4ganB7I2eHTgvfMxp38s7Wh4KS2Xi9Pe4iTG9bdQXFO
AS85iwgcSaUNLYjlhUc55UToTasPcEQddlxAseQGnA9agaHk43c/FyfFNzD3Bwks
OH5aFZd1IY5dxhfhobjKzHMVZQq/NqA0GR8+zUKnULBeDDMcIVHhCmTAmfBxYfmu
/Eqa87JBjMaVDTVO7aUknLjFwpKiwcEk4TJb2xu5tvUVm1S6uLN8A6kwsitLeTDU
495a9kFiWvEt0OulG2hcik33yn4b7StOT9VixS2GLhDGav9qiGH+HLskZC77oqxE
4nfuHv3NqDtsIWbLFhvycBgUDaAVUutUMWoATm5JisV8ADol76hpN0BxBea89JIi
ywb+2w71IbRhUdN+pbfxATlR5Z9cKLghR5uYgiw+mpnKDQ9tnRQP+bEgAzuysCYY
EvT2GTGeAwJ7Vxd9AWLXRGZB1IDsZNpJHsWuq5cuv16G7lrmdaKpuxJPu7ROWKro
X1RCYMA84WF5mrHQ50sTAL0vdiWOs5PNTg93IBn0EZzB+8D9wRT1Htgs9PnQ4VFR
kpdN4RbedCuGl9gXNft1ITDy7vfWBDcaHbfUqcEZsJDvP0Gt7YpoFHfVR5kw+uwe
4F8rI9mRV9NUtTnAH09FUDxCBiuiXiG6uPenakOPM9UdZIcLjhIvpwcq/tSsQEaQ
nxMc67cieGgSDCKFDmWo2GiEuE7Ww5KJilKnSs6eKbgf+JHdoRbDpu8IUII6ON2q
pVvievLXpCgNB9DZL1o2C1vm+6aDMNk+WmyXUmoHEaIWa7ORsVCvcQqVBk1xtFxu
CvPt8fU0Ut2z1hsqc/ltaNLf4xFD264DCUaGoVa08DHukDO3Zf4utA6uNuMetBE7
CbhpJiAjw/KehCGZf7VGdPM2s+SDOIku+uT/dk6x/FgL4DYi9DsnhNdLvLZpkkfJ
z5ecM+f7kMDHwlCubP6eb1ckCd0LaSAHD2ftpMtugUghQLwQZrQ3zgfrqLawOwet
yXE+ug1v4UVLZ85s11hLHFSJR6dLLISyV1S0JUggGT167bnZGXUNwHEIQzDhEaJj
rVABHRWzdiug3nPvNAH2UDOrT2vCwraKEPc4SGJOJB5XJ0bMmIy3hYsRL8VM+pz6
PFwwCSPT1fY5T8u0/T2NmJ0D4te/9RDZq2URTYjslvW8ESnlVUqlS2hIo6j55gYG
HHbMcfXrh9t7QGgh5K8Z/0f4+8HTLsl3zCN/NAXi93XcXDZVXBd4b+kyDPNYwhHH
XW6NJ2jaxLbEg5r6GztlRPHj6QBwc8JVOFsklBLqMp8Ro6t9inbM75lWMywFpAyl
tSW7rrsp/40ySJsTDF6HSpfKQiSlWq1AxRftFuJHJnWnWqWJr646CvikWfNdfOtY
8cI+MHDtrV9PS0AM6o46aCCvvZZboCo/rubDwFqmERHPN2lgKauPRUgzdU3FPEvL
JGqj/FFORpYI9DFgpErYqzrmBAZG9noM7UWfSlZAsgzX9Zm/G/AsL+dBs+sKGnlj
axJwR4Ahk93sh2siivwyIrE1BhDmGGolsjK8QBCWZUWZ3PgXuczvwH2chIyUZrJl
x+OYr1i5KTmhhGLA8MzT78GBdDDZMHJVJEKfSmyRpVnxP6KtEWHXxfQk4a06uDrh
6BbwrGRTTLYzJWKDUHnpQWaZafiucEbw+CIIU75Z2r0BXe6bTyDNiyFAcx+CbO4G
ilWvb+KSTcTrPfv/EaEJL68HPaHMnzyFXa3q/QS6ka/kz632rng7hoQ/e2HB+kbR
H6w085OriKJ73L2U9tD7WlNq17LOTUMqfxMwnO/+H/YD89X6gqZuHlJAsZ70J9MT
3QleTrBuFwB8IlKRetH2ItFFicOGnq4rGuCfX45IAYo1m0yBf9jIQaQ2FiztMVgN
3Z7jOu5QPLh6DFgnQjGLMXMVfM+SBbOzbTiulshF5S8rmmrD9onegDsjgTVrT0Y5
4Kxtc3aeIfhCAEDgFtkBU+hR4vHSwFfDfhFtpHTheLOxjZTpLFri8ljhY/FM/LlR
LK8bqF1zhMBh75IbhqG2W8VWXTHavhqs+tAY4NQ6ikedbdbtArhBt7hsIG5LSxP/
MkJ39vEXPt5C6vRPO6jpd5uuPVxYgiswzAx5DmZHp2lS9ouEXnZOceDE8uTd5j3s
ABxs/F6n1kjh1B+6gH+AbCixBPCoXuWpFMj+iqfqgiQkM3ZjGGNMrtExy+CgCUcm
5xy9Lp/hZKnOceGyjQk1KmGrs5xUytdKq1hPB0V7dTpnhrlqIzQDH6DNf3GGIKRX
j/vXq3sFzRRRJx+2o8/0eyQJnh/sWz/QYHki13SR7OQiWZOpqEwY/5FuabwKpnFd
aBdw0U/EjQSzdE0gfRG82j5kLIJ4JS5XKGeGwyGfmP478F8Y7z0DjalZGmDza1es
+04ON5rBjjNHVGJB4w3lAdEiP7wzWBxQUCE1zputcrjbJ1cM/Av4zjIcnW28h5Wi
kO3sAzdWvS/uin02wvMPlQru8oPfZjUuPlumKOGbumKBUhfMgJvD6wCND3irOeOk
JHwWSmiOtfZNklXBv4igzI3EVNJHfGNQ6pMOJh4ysW03le7dKzfXKYLAmpoWTtcr
pSk3gBXPze0a+0Js9xWvoH8QPtiy4ooYknusX+LGL6oPHZmHG+mFuAOTS7qfWejA
ISv8bCOfRKrHdJUYa/tEdDyB5p4wsPN57JFZz+dMB7uHYUcDwOsHcTTUWgALt6VX
J6Ts00bU4nFs6/QfZp1D6ZWRiuEyaGwwlgz6dQedKB1vPDefG+X+JGQV3Ip9TFT3
NORxXAKQk+hU6nni2aTflCCKoAQQJ6K9Puswa8/ctYBaccsbUgopfwPCI1sXoUqY
ZqJTxBgjfc35xZy9xBggu35sgR2fGYFeSnTN6Cfiq9791mI8GBBvy1HWRLBB1TCr
8waw+d61tJavB93LH0ddCBUTtwtOLgq8jRFrw301y7viGszSDJU6lNo99FnuIxHD
TLmvfpdPPra21NZsM8zO6PDP4KWbfQG6MJjp2LR0EXkebf8frw3LbMbcVDoB6KfQ
DBfe7Ln3kJmXgoJNTavtroUMuPyw4mQqz6ifRiqNW8NZp31P1YjwGBOIeedWIvvE
TEj1vVR7jmKr0lBuPjSe+oS4QTDPBgq6GG/9oO8+5eSPS2dQgN9lF3SEHBPyyWfR
oQbYLMy8t8II8Khvpb10EGBiQDs4ei0dK9gI3jDVKhDBzqPF8Ph5+fgGwbl4deUS
HOcQ3PLL+mMQdWORRWP6wSAV/KeFqLQ8rzpum3a8wCpCnc6pAY1tnUdJ4PEwMLX+
Ifg7BdC24oEboP2n59tJhPvwSPRR86p6wgjoR6nnq5jfepjoOELnSDZYwJK1u2R6
d2uinqoUIrO4A/OtWpb3B2JZlmYe7fW1IrOdef3tOG7Pp5SF+JFiQXRFbWOLSIRD
BeAU7hnHt4XjWHSITs8PsIl7ar9rw5XAZvORszQbwZNUDwux995Mav3MKXjy7kv6
5vZuo/hXBt5UYUEkf0SMp8kWCFAun3DWFa9fJuT5B2YzQQO8994eejyCiVghbyYY
xVNNgcnftCoz5/Z9uiJbvflr/4XLXIQHC3zRmpU8giX+SQFeTu7m09c3/dZhsha1
OwCWR9r/xry0crc094TXxxrxbqzG5RVu5taqoiqzH0po5U3XG0bzQ8/RNrDTKDfe
UG4VFEJdKNPulMNKjTdffGAQmMePvuZYiexd21UzvFwXzxWOqMkkfOp9zo77HC+e
wvRoI2mKWpBI+4/0yYR/C+O7nfE5kUT2PpOgMPpirbVy0PP3t3uP1R31BZ8Zns+3
N5zoYBWK0aCOCQYH8B81qnieB2xTNIC59Yn/cMZ7zNlDHk3fxc/woBA4DX96FXk/
H0OXBs6l0/DjvzVWpxl1uq/OyqzqdcXG+KUtxCAMnVakeN/wL2nevef9dywgrU2d
5iDl2GDKAgoWgM+dWubXXngnnHQKuJO0eBa7mByNusUMAtJbyOCub10QvOwAs1ru
Kkj9HEp4MkJSecP9gZiSWZcWeisiqNwrbBDruGUIIQOKVVPtn9HcobcyxFR6Qvij
yLpJk0nJgozcHtl05LeFRwy2qwpCri5qh+b4rmfu4+XiAUuEnRy9E2DU5Wam4nKC
iXzZfF/a4DFZzcqbPrnrYr6ZOAxE6X5CBYtBtEq8fIXCPdXe1ekE9nn2Xl6T9Wyl
GgbAM3IiGhY1SI2kEYILxEwzu952Dal//QmlI5/TMbFB0P+tYjBgx2hpeRxfGSnW
iQusMvvMOUyf5k9KXRK95O7KWZoaKzt28yzjY/G/JL8L8gM3QTwD8n1N9NcE1jcS
9MfoNjYLOU4AqmRwABQkb8BwGlFYLD9MB3oa6odKhrAwcGii+excQpQYkY6lyxJr
WkuyNjXRH4guh50ORu7DwHn3Fr9UKgDxjQ/rQziV3bHvpMG2J+l/Y3HdVggK/XI5
/MOEQ/Db/vK6iL8AYjX0AYsXXwDGLKYuPEa8+7+iD1saD2An5OOzHWpVlu24eN2a
p7jxZhldwYPeiFQmtPMyDtWTdkJPo/sn/OTvEDZ1RJ/qiGf/liVSIpA732qubRO9
/v+CQnJKip2k6QeeuIuW4KvUF4DyiW3pSRK0gGDXnJMJ8xJmwWdsiKjuHZDwZFCd
h7uaYLGV6FFWomGyRugKcH8sUUyfa/2/vIT5ZqG+l95jMC211PxNiY385sqhcKdB
nsf9PK/JDcCglTFfh4x0hWk5KFM7JmNa4ebH7HXnq3os0gwaiDtiIDq+sFVyrjHK
csOYwrrG69WRFSpB+8pB3L8zsVirdqr9CMz9iSbAEjsdtAY2x3lP55ooRcgnfHuG
wInRT0XcxBohJwTBSkAh8KFUahXvIausiOq+DaYIJLLn8r0pWI+hS9T3RxiPBOud
7tJB6rmiBJDvZDR2j+P2904lVID0FU6xfx9/0c3GMRdKV0Ce1rJ9o+pIw+fO8+dR
iGarxmo1MzOx8G4mdv1yCrWuBiDTdXsu5yo6eOjpXe6IJhUSNE3xQwAW3F3ncQK8
e5x4Mt7EqTknoLmhgD33MIzTaqyRCfRvZbaToSeMHM0IVEKwtiLse6yRb5/DY6L4
2C+bN7u99skX2QcXa07RmEejY5YL7ope7D3Buci3n3J5RmwOzDpbXTy8F67m1Gb9
XdoTqBrY5bm1lxUwsUSLTGjXazrVLMHtVP2pp/Yw6SIQfzBgq1iGmuJdGJpalRzM
ri9Kl3LgSzDWyGPEBZ/bGOg3s9Oa9stij6KwbLo4Ryx2S6WXWLZeRW+EShxtowZm
meBOMfe0Ib16u+8Qa2SARZKkSeTNqsP6WNiSz3QSUiwqBkXfBK8ejk5zTqR+Y6TC
RPu4Qa5TKvlOPTPn0vo95SrhGnA8+9iiya3OOz8hXHx76NaXYrYeerz7umKxZzhv
dRhz1GHpTp5G1JdnD1uL73o5eRL7jUeEjlffMzp8XtU55EgiRKjRz04OhVNBUWEw
w913NHKUNFodizwusErW0zPCljm9FW2ChuFwNF0o5tGUU1oWbODmDMkYoCA1+IwJ
/cpk158H8UNHP2ZKHm2/6d4Rs1vLVY7ZzXzvsuGnHu2r1IZfXy6iGRKRQhtw9nA2
6tHIZNAMFwt/8l9LPIqpb9LpkFGmpJfT+IpSeWVDAbYMxSaMBCCM+vpp7bLmxKi9
2jClETlel56ZQWNoqk467G3ngWmn5lpggtRDZpVJ4NMy6R7om2zG1sVuHnaLOFPM
oxR+goRdADOpFiVRFOrisHbGJM2yWtgcFHK1za8PZ7tzyWKRyz5y2cjDU8+So827
SpVi9v9Exp7Cg9JciJJJrlNy5bKM0jFoe8hlBmC3por0iWH3hJHHi3hzlBh0bNE8
6em6SMT47f7Kzl8d0/I1jlvyJNkPAewqaUolJ6AZll5EXQxbK+Ptsv/t/agNeJ71
NK6chcleb/SeOHJntLYPTWmwLjgif8CpguL514QrNQuEcZs4ItfPyrWgC9IylAHa
c40P9WcfajMJ2Wj4BaGTdjK/RMaKlElQvuhlZBZaw38q9HSer4vVo+psrT/zBsSS
HcIhhnoShdqCnjiZUJqDfGrxAcKPIBmOGwbweBBDHkkczy8aVFDVkpkY7gl/dG0Q
JqkGxXnkYtO6yiE2TnJlM8EpcJmP6efs2UUTK6cLdHi2R9VPqDMRICdnRGRv2cPG
TaZ9CUJadKJoQ0P2Z5LLeqh6gwslkOvi0SjHKlRifu1ABO4iR3AoVXrWx7RaYGSt
Jp0CylP9hznj2St2lwedKym93ftNNWQU7i+OZ40OzIQWWFxFt058YswqJRWAvlVu
MLsVumyc8I2WSAjPUadiy9+HjkyXt69Zvv2yfsd1yEBSb+wEl2rASAmZ9HMFC5KG
t9fCm7Vgtx6PMThLrE8L0ts2LTfjvr7wk9N/chUGVSjkksqOEFgC866afI9rvcgB
ixNcJameaX2NC+oPyUseWLn6bRPb4VKW9yncnGClO16K2KRHsAhlCkUfX9JYSS0u
vMMpqztOjRcHImyTusmTy/RxA713gxS9aIcNezjeGG8qFCCmD5WTewQnqj4mntnA
bJL84WzkiPVUVMxAC9PkuQfmg7hm/cCesFgPnNAH9HNObGlqcNxredJvJjIrvO2X
L+errWfMpqt1l0IGjphd9O8E2uttJFeLx+MarxzJumNWvW9dbf83Rzr8eW7GuyDq
3EDKD8Ir/WBblG62VvfenZiVhI3Yr3vVulv9B2NgzWfofw+lS2bBIAmJeIPHZXar
VOmhtiTspm5OUPFtweutf/XvPwwYo6CeHDATJv6uKXMjgx3a2wfQQpCSwD9MonrZ
3xlgmbaZkcXskMWWuY8nxE+kfHWOjry6PFmRgUwE7p6+0g85CMQaWzcIK+tbQxz7
6w62MrDrIm9T8MUaVLU1aVaHI2vX9MgGQ8XY9zG66lrnFeiZ82O36w58oc9RW1n2
TtZvHjklCu8QHFGeVaJvYlPHD/dg3M+788DJ/scP4bX644vKLF1C9U93uHgXRnpR
3J+SgFJEHKKoZaduF3UR+E7BOYrFNTOEvR2U069faeK4QcftzBVK9hNVmr3P6bfb
APrP8VWXPC/jK5Y4HQmGmWCYSUx0OjHXXC0WwVHBGaFo9WAlTI0XswjYLdfe9Uxf
cWbuIhsyuFl4AdFnfs0XK19Fct3E/IJjRIrlQopMsrYAr0qh4HeKg+2tOtic24qv
x6esFSJflyl4rvYdj1Ex2DYadFCurnsJ0LPNLuhrqH/0jhv3HdfkNIwZdaEEiC/+
rg7g6RGNf/mo6o5eHffw3Dq3XxMDwOVUXKXhnUE9hrKsUrmt6TEuHZoX+n3B4saS
smZmd4Dc2z9G1IFSaTyqCP+vAXtRm3uDUjBxoe9ApZUzBzPoZEg66xtB3qVBvDPE
CXEi/vDNXzUqXVo8xYTNC3iPZy/16wuDCyHVPMYinKbZOea8xj7YD/A3iWahQDpV
g7DGL6bbj+pmvScbaJhPYPt8Cfb1O5SbupZ5U74d/8Ys6rFP0R7jNITTx/NphKAK
uuX4PhbcPKSC9MtgIoTmZwkcnrxcwxu2v3O2VFFg6sduj03GMdWH1XEZCRMr2bAe
ULJzvhYXfe/cILFnMbQ2oFzjjVIgPNsfJOFfKz6K9024FyaTULSKusft1e9IqMFb
3AaeH9F4gRdgGxxRopHGuyYJZV3krts0qpdkHdL6N8FSuWnfyeLDi+ULwXg//In1
+RZBC7eb5ZGtHO9tgc0K0Kz9fpX9IBOdi546xzngVinT24vajLfNaEO+NYACcyQE
CYhnMyfQBcl5P7KUv10rtIHkFOWtgHGxl6fTrVO6SVqNrpbYTOOAlRDANimA6HaF
4Etpji0+qriGEwmCK9boxO23W620/9rFPrunhRDhNO88nrRymOPDV66szyvQ5RrB
e7ZwApV6M6kXKz7fmI7izs1QJ/97cKudl3XEEpPDZyMAtfz5nQmevOUi5kbC4p70
i/MzZQds7zMBk87MAAJpXqHNdhfROxFprC+I8fZJK3jvSkpVM+8QaPYj3JfUpmUA
AFi9Zel0TBAzoCY7AHPv69gkigSdE9ZlFZV+T3XPglmUade4UKTIOCGHW/RkCIu6
Q6+N+Pk5KJeDpBI6UW/xTkp5IBPveBaMGw8UaB+HHFCnsA7z8+FyaKtsMglLbZmt
SV1yx8/pEiqwWFL5kDJ3lRWLoWt21XlmF+e3T/n/cTCARtsAoKs4hazqLK3WIs7o
22AeBlGv2oXHN4ZNzGbdI843HMOTuySqz3Q+02AN58CgcrILXgIh+xwFUMGVZyd6
vXJTNE7ZjS3ctajYse3OUOli5waSu+8pdQBH7kFNgCnFqK5oYhM+EpUw0jV5wIyj
KBm4lFpYnw8Ce8u5a8rdSyjBEZnOPnq+Bm4KaGRBC+NUDljTI/AOC3VEIndlSPh/
o/iyxwyn3hIpr/DTGtd72EHbw25P5/+Efbl7WCVR14+E7guJS3gebXbjKyN5qxva
w3b2MKP3274S5yImve82ICadfJGduw5i/lZCbU/qFaDjObi7BjUVwXnAzfSTsgpi
DvnEA3Dv+5zaViR6UxQZUYL7wCcSEyxwb+yyD7sZ5D0aL34csLfkwMW1vyKmIdXt
mI+losM/fAC4SBGFjlUcRI/df142UvMlxgNxbaCAYNSff5MFVE9NL0vBJXIo94Hk
yga9BU6aJhs6cNbK0GkZet/ZDK9tCgWBQd0Ol5XlpDJDoJYbwI7S2SbiLMytSb1s
iPbY+dREztR8UZ+Dtggg6Ne1v9n6gr0kTrEY5fMsusAsyaWnSGbwP9iPpBA7r6ud
tCB/lBB+kCDoThvRiyX56v9n4EbXbSm1u9mvsEzARtB8pAV4fpz1BJBPOGEwdaNG
tflqHAIS7REzvdPMS2IRZN0p+SlbrZCUBWy5SPhU11oUwir0vm8wzRbZbR+r3QjQ
OPyNMiyN1nDR9tWUt2wAj8QL+4XG+WecYVXpmIb0WSRROK2juoiZ5ta6RqD3nQFc
y98da2m59T5h2kRbkH+19rt04j3yo/0evi8GJpiOkDBvSTzAMfn90gkgnrZRrN1L
+ktqi2rO11bxcFtz7qGLRO/XQe8cdwowcm4eeQPWbbzIrzfAPkLmrDRDbKNJV8qW
3XlCWozJ2AUoCruHu7sLEuCnFyrLisciQpvaFIeffh2cC0uij0cDXH+rwQrB7y7y
iCMKYCyHvjH37DRNq3N0I0dRfbMU4ahbdKJoVqAOdTMvWRsMth9Tx0S/X9oOZKhW
0T+ohZZQWTNAllmrgfF+m8KZ3gQWZOQ9Qe3WE9o4fTv4jUYaFho7hUfBcPW3Mi5u
Eyr+SBMEPJmYgS0CG/EBXXcIkDn5OxrJvA11g2jRZQJBxIJ6a7Rr5C5DepzKCSVv
QucrZp2x1ObSpd4h9plBzRP8IoJfZPLytD2Sh2BhV9uap4bZdO7BKn9YIfaJrDFY
9LZ69rmj+0MaNnDbQ+ERjY0KFxBi3VkfY9xryAs2xuMPLdgDl3AtQnTwT9Gj8LLN
ccGkRDUGWbGtM7o6SMlJxqhKE1ZxW2td1vza6HBOjyB0tLCEsVkX825t8rHHXF2H
sBArEQjPEHfQ0Sz0+wEdM3iGzqGlct3DmDfgZ4V8BGDF7fmBZT5j6nqaOoq146Yr
gRvXoh9Z6w6LNFDGp2jbqwJ2JJvlqYn74yZXm9bCEXt9l57iuP6crA+mjCj9bvVP
0+d6v7bd/jt0Em0vdBorsm14ZK9X1tmRaVwsmQPgmb9ufeKQOMcbgF8hPq6vlgcd
FArawFCTyuJwaDKPiQbivE1jNm7L4d8iN4GNJyVyLzwCang9iKCgPPJoptE4kF83
VDQ4xYU0OFQ+dWguLt35A6oGXebLHfy6guzeuiTdO3GjusnHbOmmvRJXIJwwA6Xg
DoMleAmxN6YD8wVoWUONwbldhYWI/mgQ74WH4T+UrMQ4zGaYPS4sfXbH8ScfKRUJ
YriXm1StGS0hodTWnu6s395XqBK1iWbhnzu9+ScSApA5NKih1pbog8baH4INtkkk
K0Rqy7VvPOK2I/NLCIjIGWOxFjznAuGP7YR1M1tzITpu95BjmHkW3WKnIBPnR0d/
5IXecoA8HkDOn7I51ZB4FH8x30kONyr9NwFuwkpIknJT92M/o54KQjo1txZrDX0V
l0zcBEi1QoCKNsjVKdbk6yxfWUga0nG5bWKhA3f5Na5V7o9n3/8UDCIdIx0yPSpg
drislh/7WNxDTTcldswV9yq8nKeQDR+Jhthd3jGc7hya08L4+lszwrYo5bPpfkon
XP8Xz1DGE403l8ZPBuFFGif1Avzf1SD/fweFHqF4sW3GFt8nlkxHZvqpz0oPOBNn
pYHdLcc9taED5PnrszxZ0vIbJKoCYiEcfgyTowsinPcNcZcDskFW1dCD/d8g82EA
TfSVpzvjyz5pK3C48zWypIE6uk3Iq6aB7/8MvFsIht5tjsJw02a+gwUuSO6yrtoK
tkVGbr0heBl3Trbnrd3cnM829eLniBsq4KxQpUBZe1Do4iyVg3y251WbbCGu6KEI
vrSUKVLlfb6r7SqJoGnq3OrUnj1j5LYlW4fLOTzaKvUPgIl+lhSOO7Itq/fiO1yN
6rsFnLOslFB8pfev19kg3oB5BqgjuroQWtfNa8mV9s5MTsh++KKPpWt4NfF5gDTp
dTlgE831lp4HSCBgtMEgjj3/c++n9a0/Vj+93XGP6FJ8tdu9+XhK2V6zfBDs4dR7
CFUwP/wWSiR0UhSqH0CdXFyTc8gCEXa6KE6QGXMmiG5pNu4p2E9PYvKjYmdWIyt0
ZgdwreA1Y/cgRKMz4eNuYrzPprMzhI/NRrTNepx018aQjtTNznXXQTGQEnnw2W2q
+s9BqeEck96h7eW6QPaNSWArzQ4Guy7oSfM2kgSwxVJNrNCRLv6dUfsPxh6tI9LY
8aX6L1iIsW1QB4zw2GRuDsRMZaxy+U7bjbbZ0Z4D4rlDhxabvzyYH5jD9yd34ids
1KQPF8+8HchH1fOjdGfZ8dcSQOZtBSjTDGUKBw0hD/eZ2TU6zszYoM5dYJCdRq6h
5BlvzEE+cuMdsVD9UayJMyWRJ4QhYz3qHQLUYyaGwWzjzDuxVq2cP6NCsmb1j1t9
mG858pS7ltL3Au52EKy/qgYJ73ZCUV6JGiA1U4Zx9hbV1gHhHE5u2mvQ6ekkM4TF
V1V7MeREcvqevHoqX2YL1ZcfRGIjn2sT0gusCBcTz6AUxdgf13iEsThuN8CxaIPm
2/2AEatbcWZxvZG9sPRDfkxuM27TS2sRGaz37vfXKW/zbu3hUsYtgwRcV/SGvbtp
I7pzSiHfO3+rRXm0Le4eXf04ApuEauFKiQ+gph8Sy81t5MX3VBDYTh1mnIV5o1xT
+Jix7b5JWsW0CNSlg9NE3MGxTeWuPUoBV3dKaIdUowNrU0i0LRoDexIgRi9Kjt5E
ZAYY4l8r1HkplOh56dXWCZiBLBi+pmlmRwu96aruriW16bzZYUUZ1EN4uMnLDqWA
1YksHZmc8wxgPmO1S+Q7mhODEcqJvdsRiT2oFWgfX4rBbCsUWApDaNmkd8m9i66l
4mra7i16dMZO7B4BaT0XGhgq/fJtbQAtNI/MBLuIR30YSpsbt28aAmJhO8iHmSe4
PAkUhG/MF4putbO+VwzPlASHw9sbnLC2yp0Kb1u+ZGYUUrMyCmJtxtlKy3P6X5L8
lcivhffxng50hP9Ln3y2VdA+ttGOQtT8hTPRAa1L4TSs2kBvZG3W2NYz6b16IWKX
jx0tW82SHOiwVTNMgi3ZJpZc5DjdNsEvZxgOljyz+UorFtUDMskK9TrTHkJb0ZJ+
haPZyGiz4cYTbSaUQ3DnUkkm+7Jk2jy9UolgVme7IswARlSZqB1BI71RoiXyS81r
flo9+G/kpSJwO4HlGA+GNVkWKGSKB8LP9DR3kkDl5om9Jkde1cbT7h8PkPDiaHn/
BEJ80E08hcvsNhs2r6gwz8Ya53X4sROMFwz/LDqHYl8tyIMyTgVYCqNHA6XrRMyQ
CuvyuehebyWG7g3BC0K6oD94xPxaA3tOpPVV3N///bzTOxiLXwQBaBiFzr/rq2y0
ALXIBhFebEUOr+YpP2jwJGzwWd2DvH15yiLxaf3aaKpO/fltBxcGdyP8k0pJ4kuE
amx3yxi2f1PPDzz4NLr05zCgPArnm17ePw/qKUIg+oxSIn6gZtrBP6CWltqgQAEw
/6BgTL9WDwn0zxe0bFnB2/zsE0+w4ur9xXeB81Yruj9bzLqfveBv0MEoAlIT8R2w
TSiy9xyub1WWbG+uWjiBRDoGvQsYVqAeapN1g61/ILkU/AxF0PnDuzBmUy9s0m4s
mHncF1CVgLWTIM7jSvI3kFFZix/Vsb5N62hepvOG5zjHhY7z04c2Oe1UO4gnr3Th
HFSP1Z1W+jMKRtNmf1xn1H0G5sVDTbNPMZ1A7An6q/gzPftVsoufhuCUIPi5MXFu
rgnYt7izb00IMY7vxcHPfTUIWzotLiZ2g9ZO9LVuHTudorCvyhC+rkNMMEj+BLyZ
JJjJywquozy1PzJiWXHh8oaUHZbrnu5VY3CToLt+g6snFXQXiaV6Y9hd6JeN0FNU
uX3K/ILnCpcj6pytsAe0A4nvPXCTnWDqKx4EX77fHVEL5vWg3kBJId0cMS0Z+NMC
9rZKqJKYXk5MiKkDCr9JFeZ9zG/vulQKx9QDgbj8bYEImudK3hjchVAknLbI1baw
V6Cat63b6AEGpOKahwEaT4rAl4lFlBcOmCa29OkCvB0wyS2gl+E5nKrkX4Mn4+ej
u8zHW+JDTCbAf/cczS54RpST5odGUHl+GJT+7wLCR6T/sCYjrvzZuE+rSp2TnMq6
YX8/CqRmX68l5h6/XhkGjGvRBmTwh8//cjj4bQBN0CsZKrHY6Em3TQANlvS7wnYW
rPwlWasdnRqE/3JsO9P+q2zyiUVxJSKfquvvQ8WWe3vNFw2cowtwZ4Gm9LNol9zI
mggMOf7GCj8CsRA5tKrpnAn6iLd/RyDgYvrXQy+JKyhMUORVfGSverca9h/jK3+f
DAgJ76UP/bOxYcKq7TxoC0Brj/O5QdpNQ47iIMwsySVWTo+mLfSLbCQUNF942KIW
u/3hnHiZTdcK75qlWDOUz35y3/f1R1lsTaGoEdA4BbvNldd8Jb5gskZigyJ7Cf3N
lXaHgVw6Ve167fB1Wgn28oePGYHPJa3rO1YQtUNMF4SEBKZVjgBwzPVHn4ksxWPz
zygwD0oglRn2WTsKXgG9UYUl7I6hAXfdrt+foVhEca3duhyNjZ0v09V2D2zBTdso
BstXQNPJh8MPkL3CBijA/o/oMwHQxCHbVoJSUuelvFLAWaDhNVhgYVTzotoGxjvt
4OuF0Yp6edSH+YTmMhRvUlTqzWJwn8FdOUCdbNWfDS8g24X7zmwAw6AAEB9O3t0x
7gkuE4KzqSVzevERKe0iDUO8P3D1umV/dtsK6j1K3Pf/x3IJg+e5ypk4aeokUx/x
D4Rt965M4CFY8ZmEs2DtunDcrKAQi1N862Tg/+hZYLpD9K8dpQuoJ8m32qUejUvP
YjGWEuro4hWxJvMNsQcYJK+tno8l20GgODDGBNrFJ/GRINIgY7QAKxwknuSLCQ9D
o12Tf66Rs1MtcnBVbd+FwGaNZqgupl1nSZZYoJDtkRRui/xxxCZgtNYgYNLDqGsV
IwRxs/y1Z3R+uxrNC+e24BgAJHzl3yHse+y8eUT7n57wVbI9f+OWo/6yedDpKvJP
COS65Ks0NFctw+Pez/FdSYZ9/O233mCylOY3FigH5y3fqfsZEY6UWKDHcoWiLQGt
AEskfXw7JDF3vKLgACGXLbtRD81Sqz2hhU9PPe5+KIMgL9Gm38ugDEFTuofDxhmn
8+AVcrFfDF77zfQnRu5si20JlV7qFQAhvpZbQynKYgPN+T9vv3jugjrARRfpQ82a
Qe31Be85gHose55b0fE3CoCVNzrbdGoP4DYPwfg4iT7tZkx8Vz+KZ1Bk8/njxEBm
5Pu1Mqssy4aF3UG0/hH20EFK+QoxEEeFTU6ywf6VapgOZH5UwXIzjlanIGMsWsYw
3NzdFIZmIzuMq28i2iu/VumvenM/f95XIFfSi992+znOLQJI4AhJMXvpKeNRA7mh
UqW27DABOs3IKEZyNx6sa6V8HPPY2jg4VhwXJmE0J/CnZw7NQv9mOYpeH7UgC3An
In00JoezvVCsePJl/60l7goLFK3VYSpDMfEBli9sPNXKK22ju+O3g2rCXrla5DkD
4CDnvmVYT9UAZVjCBsx5U7N8ahnjwegllbhmmSB0tXdOFlEUdt5etJ3wVdXR5sOa
TQnKy72g4tDCUN36savnUpcwiyo6NYxvxmE0CCwPo/j3sFjm2KwJQK+Ogn4DabSd
BI3j4oQLEy4NmNgO+Ku/4wbeRLmHLGwTZcDQJLDFW2wcQxeqcZDGO3EFX1vZtKRn
r6f4eMIg7mKAsOzjLxEZfA8ccN3PZXxaVHkt7+jDNffQpoNXaYb/PkH4RTstfWdB
Us5t1KbpjqGdnUEHjLAGpJDEPrJreq4BnopkUFNdSrAcR24/fNFHFqinkRkzRkHv
bQ0qWm71Q31FG1gD8QZn3gtseRPRD96/CUP7pSmQw/tRyqqyDD7c5iAwqZCrlHSd
PusC3O9poKql4snj563u/9BQN/pICVUKRBr6mxDJBo5dQCO1h78kprCKMEiAdNUe
s9xXq2qd+qUxfZ5ppvaIKc0TQxfU9wHj7tisGCivyKhWBijqLQDpqrScE9K0uqko
mwqbZrHa2AMpkdCQE75Cy9yD907RfXEtV4/sGNWWu4U6EKFcFn780IWe3IsIuBg9
6g9y0Rq4EZJWFJkogzY8m6Wv+qNznDV9g+ZeXl61ldn83pJI4njrkYvOLFm3P0O2
jQRmkx/AX/n8cBUXFfk6LT3Nh7rBSjR99ud+/TlDw9g7ZA+6wJBEAEEHQ34fQ5gA
akyUSzS2sZNQnJ8mE+EelsAu9jD5ebunbqyWOvoCPBiz2qR6j956Ya1qIWnaOKtC
zFIhEc5k39K6WY+WPZx9+nqzd2cj6SAJt+9eikgXdvX9TP4TvFu8ubeUkaxH8g8X
tEXFQwEMQ7i2Xy+GPhdrql3s6OhJTWHerQF5UQI+KHtQb7AIB0KPXWUXS4HtDU0s
eu5Vjj6p0U6B30UaoBr3jDdACrgPd3rt7KrxFfjft8vd4Q5tA0OjXvcmlU0ZVPeH
BSTMQDHWlwtxCEGs0A2hyf6loc27AzKP5nWCN9KwWPcrMDct7RFdSYBZHxqg9kW4
OGZsgcoucB8tQbFXe1eYFt5UFmHWdT+36JL71p/rkopIfxSY6++HKkt715LuhhmQ
a8Vggz1eLjVmitiXNQ0/ppSiE18sW/RuCDXMM/GyGjee+egbqLCl3OnEBYk/vUdE
LroFmFs4PqG9XEWVZh1H2H3LUbQ2pZIFhvyMyemcoQa0dpCwhINOfqIj9STDoGpB
aKKYNhNqKTT4LYMWGgl4TNSmfKw1XpGoRbfTGyGt/SyMQmPXtxjlJhftm1n4ehug
efYhagUJONScgO3xAuLNVUGLyZwdNc3oDyjnNXPSAHuLqK01MZatIs/PCUWakT6M
qO4BLgApU4fe+VBP1R8HABh6qyj7BsYtU8nKiBYm/7oj/chSbH16BqKvtxadPF4C
Kvt0EYqw8dwyz9NQpmsJCO27qYWOzEWYW99VL4y70ao73SilGIpCfhnUUesTxWIv
XbVHasdfENsk5ucTxYWTdm3xxDbEv0H7mhdwselxIkASBlNBe5lRxkWW8YhQ+7QQ
h6FRjBJhOPBxqGlloiR2YdC+qHcoPQY7aI3wGV/jLRnW1Uef+vp+rYZMurch1wPO
Ou6rzMFUKMfGP56MfX3apqQXO56bjAOGqYRAlaxaiy7d2UHYRpznywm3YfpeF8BN
GFKZ1O/pu1qsMpwHxgYMG4Wyf4RcNeYW7fRBI1afc0/+zkVKGQDDKT+nmToz0L+S
mfrCwioQ2ayaYQGTTmpl63Bk8Eyq+TZ0MqmLIZtyl3+9v4gohrqJVSxHM03XdqDC
8jdZCC9cIRHEuOz+P4cJ5otr+X51naEmK1vqFiyX/tPpoAfhPh4uThqHVFQPUQiA
nAKnhWIjjQX/xDIUcI5sAsvL+DbvX9LCs4JMia6jclK7tEIudtjcRGY6UMTmBmJQ
7ahsXQxSs7ntzvK1Ek/kZzAK7pZdgwfoG88iXPWSpZbTl6by2soQTJI0AXIlUL6h
vPtjIa+qwH1kf9jNgFrTAexvhjIXnDKy42yUAYyeFmA+98xdCv5sMQcY0tBZPyar
TvEZXFy2nwYuSaGDiQ7ZAijMXH08x3YSHz8aQFaUG4pQPsE3dIFOPrbeHB7I2Wbw
tRXGvTPXHi1/kQlyFHQZdcNoOl7KL9kpTHOlcxYUGGsjry0X9JjuDbBsNLhkEyu1
8/DS47Py3U/jpGcjLVHfN4g6StTiF86YRTxVrG4TLM1XqxjPdp3ovW95YdRDKY4X
ONDYmX+2ZR+G+uTZmKpUvYdfYJMbusGlbHdeWRwP1jf2D2gKz46zOqDRWGb3+M/v
cmkv++KA3BF0/+I4gmNkag4nsDsRn/lDpBGMCiNfloJzta9PfR/N16cFBQKopEE4
qTIvCkXVdHn/XwQ5BOW2RMI7qUfxgMUnZ0NKhg+KGV7zptJ6S4CA6H4OkQxo2w1h
mUY1uAAaZaDxn7oP2qy0AJddT0ZQgcsy4biAP4h3oo1pAS1wY7ZhGobTndnOMUfC
9tGbyjZkO9RFKKyPhMKpuuji/TtRX3XewixALPhFORYyasUwBPMiP8ELyPViRKGr
JR9v2rX5NjZpkuRSSjnqvsnuds4M/wpXX+v531RqaORNoCtEOZQoedK2pM/Glg/x
giMDXtEK7MKvXisE80SkHVpCBDK8seSDqA5AFdaPIztRA269IMWqrSMDxJ5qdiP3
0dYSTiVxXJJ33WP1MfMC17YBf/dUBRZqLzFjgdc/9jkCxT5sIemLrti9QFRxYyQS
jWeIMrhQhvib5F2neRoVSA1fUTjIKgOfm+LfJ1oSOdjOPsDbxSGzITIVNK1kuo6A
ZnDidmJ9qCBlcN7nmRfDjiL5Q1Yhq74CGuLRFi5eD/ZIvzX3s3I/9ZBS273Ls1I+
VsPkPOnwREPi+7kuU5o1UPmXd+iOJBJDedaP3t47szcve/GvKKiiajrmc/e+oTTL
ijrLF1EhTO4KlJS3739BZrW4vAcl54YTODNwMkIq8yfoDqx2Xx5bczkB1mcEZ1AB
ssuJTL6RClji+3YEfi6MU8fTDRJgwq3/lpiRJBfowzK81IQxRMxHMUvpbhPB1ujK
D4Xotv+FaoZEcjAgiMuCx36g21TsNl8Y8SFUYwOB24PNJeorGBqUv8N2A0c2Ez4r
tXIIrSua6gGrSiG2tgbOLQEzyiUs0LS6kgTuJYNxxkjigrQ/o0TS1qTeIyn/0A3Q
o+Abq4ZEVJz8iaJjW/KCSzMfyoYYrY7nG6hVz7QOY+QBopiqfPFod0F9Q1EDG1BX
ZtK4xdEIman9gSMsfFvrd1LsF5bR+7AmRv0TafZ2SMl75F+Y+8/ONr7ylIlbV7IZ
eTtQ/tSBFOdVOOSeAgKiMtxwUOopCcguF68eI+2ZRHE1heG06/UDGiRs7fPWNzkY
jU/G/KmODbvQmrCshBdFUtTzE/KwjtYXUkwK4clhMb0WnDXElH3G3PCPOkNJeWlr
gqVds5aT5APUcnG9nehN3OBLLqund1WLYOLyIGs1KdZajWFi0zZfr9/s7aT2gpSz
+9uHI5yebGigCrttLMQWZo5d0Y+HMdlTYD8CUldlvQzEdvcMA67ZGEH1A2/v4U5W
owkSM+Q0+/kPO5KfxWfXR3HE4NkfPCHYd72H78Cj72H0lKJRTxK2gstNU811OHxc
X2FMZqFyh4r4pL8oI2tYYjGXbwSg3YcnACyJORgANH1yUctyc/WdSMv8tlk8Pc5x
y6T0qjqm7yXn4Ig83UKirMZhxU80rO8Yvs5D+B3uETSj4Al/PUrHZ4UaMTLY+fua
CuOVvLh2tpG9a4s6l7Xp2Exv8FU0yIxlCLvj4tPwseaOivpKbcZ7yu9II/EHNPL5
lctS+ephagSyahOPVEUCL1l7EgwQqnYUrXEE2MvcxIZpp30vnNh2A+jtNi0xmY74
54NKgFHkOKUzMaxtfjMAZgIlvofb/Xvy8XhYxeeVWUlVViOYux5V4KsZ5uCrRo6x
HvWexYunjixtwwHYGwdvIpzWEWfo5cUqucYwPOJ9NS0zDeYgLovmZ5UlqlJuUD3l
iQbLM9D7SPiNJ894xlKYX/VsBHQdxEy04IxVqs8hRXk+GYkipigdGTGU0hOypini
apuCsnD5p3AGZw4vJ5h7wvyfUsGwV+49nfIcJtqB+AUXiE6JdBtkbfJmDb65ZtNT
dzZl4UTG6bGi2OXMAFSFyUCQR2uJh5PXiyK3zB1JcQhJcOrPTmc5whfbzJTb8pFN
Kterp6g6/pm9nfFaOyPHGvV8gVJaPa2vz0jaAWBQsUgTsptxq9pe4nEophtIiskX
E3vDg8ukuAKHEnnoN94SH24T4R3fKYFhR7WozdiB+YsfHzZnzSxCcDNT04JT3GuY
nU7VH0b6mKxzRxp/E0RnBoQ5HWf3TOz/fDMHrBzpiupdVmgGUVHbUNHwC5cJn07u
3/0s4tYFPij3kMCgnLUPZi8WeXCOnfrevss4F8HHV+LtWW6QAgjlrzixcZtFSRwH
56JUh1+SdedB9Bvcl/mlNvn0k+E9wsLpq8LdLZ/6Le7xO/Ww+77rx2hKuuYp2Gt+
4qx21U8xhf4JguPFyqLbwSvsQMZzEj786AqHdEt6S1cVn6mi7J65DwK9AqmCzr++
7MwIubssdGBXZL8w8VCYVh3mpyBdHR7mjZmw0cqMyetT6BGkD38HSaD4ZTcd1vZv
3wUOJXn/KIbxKh+4Ephpnm5KC42sDTH31L4forlGqzH765QQ14pz0MBHH4Szkyo2
eXp2HMVM0VsG06IodIFDw4AntdlZzCDGfwHPqDEBXV9MQ5uuh54xjmGsKSTpIpZl
r7+SEuXBWxB2aPi1dOGbebpvSukpyVQwkmF3Pqcf4FLSCGvuDD85H5lJ8RI34Ixr
RNKok6fXqZcy/LO4PIgTDldzmwQB/pHSutnvGflXKbJgqSR3vZufKgBcN9UoFM/8
rW+13kX4b1xLGu+GeeJ7HEqkQJkSansnWv8EkGJEnst+BgsZpdHOhwz99bHeRCZg
+hxaOlWK0YlldUS5YbL3jycYlxqz5qu0K0gXGBMExdqCGpckzyYLROoM7jtAZBrP
DQwhw/2Ua1fzSYavh3A2cDn+sxve/EUJ88fzPeWUOMlRizeU59K8ZGyqaDSIwkV1
fb/wBt/nzKddTZtRdlq8C2eL05kuhZ8Prby+GnRRQeCQRgtoNe4yZ2sGq+Z2dy6i
mKPTQxvnPWkXrjmQ4B8wK3tdL13A+dohGJzvLxICYKksWmBA+FZXNenMuom5IpMG
4zf9OHx6j02/yT6yo/gRTy0WxGhRpc6Lvh7KhoJi+H2nqv/3liOJQ0x5Ke+A3wSK
D7wobFUrjvV71mr7vO7SH6qX85gW99JWa+XwPYog32nX7bR12y3qGc7YyFg3ljgU
eq6qhp5iIiVyhIOra2Ysbh2ZIXmL5hU/r2KV5tMl2rl/E2wuaWAzEP/Ss8sWvkBX
8CUgkA2bW8QJDrTWoeOfyJ3FF2zPjj74a5Nr1QNSZPh8PS0KoWbE/iPZeYiOt0GL
bZi5Qoggh3GsrbKAfndwQCWf9zG0Dg5TnpB6iLlG3jB2LZiw+RxvcSFPyvHBqMkK
y48YdUFRTxArxWcVhSxCtOtckQB2N6qRoALSBL+Icwl7hB9KhDr+mcQGWez3G4i0
p3gCC56rwVanReeHxw5+sf+DJNo7tUsL0KFjQ9EU/LcZcxDg9kFbGcwTylW7b+cO
N7OCvGKfbEgBbL9rbH7AtT9VLi10V8NHWaxCcHHfApryEhT+LPZ5tdxQQaH8iY56
Mrzw6f5rYtNWUOdaoWolA53tAMggiAdHOVY/bPI1eKK2wYxIpUfWjVldt5MAyHXn
paGIkceMoVIKKmKhduHyJIDQP7ZRJC50dk4kzd+SiLA1e7dzDsTPVaoyY3Ujwmx2
fKQx86AvQeHqZMTf4l8qvUDgcq1j9+IUN3APRoG/mnMhn9x5kj1l+/68xr5TCpkr
gM505t99up4YZfcVgUbthPsJlimdhJuBWv6Ux1o+dFK3A+StxcsGb7X/08LXm1el
8I33f9TS7jsZgaFBsawKgIcJ20ejsKzp134mtJGb9HMa8kasTFL9ONyfCXpunGjw
jSUh0tjP4evmWu+1pLY83lPcAWH8f3vlB6CvO4FXFdit9dVqupQCD5qQVIecsq83
KUnoClW1UCks4cBoKbsRUIn3jvi1QXTEcxQOK592icqE+r2kusL/8u9X/Qnlku/t
Rei+/4JwEvPH3tQ1Q7Xx5aci05iu0M56gfBgMH0rQa1Hdg62FftjkMtKw/iKAa59
JhbgEEIu6w9Q50hW8KgQs19glcNbMezWvKL1ox7uYwfFoxGbBsni8QV4tHgjfIUS
6QSN3eoDXHNofBF4abCuLYX9ylscB8h5mdLbf0fsqYzRHs4pzzMJFAE0Nfzck1pg
FsaxI49wvt/lADZEvs8v7k9ZnvZBx1JcZhekChrtl9JoSFMqTR7FUTFcIXdAx3qa
mczqVexdxm3X3qjW9xQ5bAa7Crp80swckPWAtv8EvcJsUa0zBe8Nl3fqvwIYsIws
UQr85fBpfvbqyBX8D3+ab4hv/1fm31CyDpql7V2c4Lha8qB94+McpqzO1CwpwYNB
XD9mV3MO1NwFEafytMcFGnaIJHzwmk+VKb7uqSRG+NI5X1HGX6Z08JM09KwOItDZ
vS5TDCM8zNXjaZLEtO+lYNlUjtSvXtUvPSFs6m95ym04HvNZorgzjLCqfqQi2E46
mPiF7hLlLaZrbDU7h3uCWrmB/l5RB5MacHxwLqVsm6HICuPiaoh9TvMJx1grNgJf
nUOK3I4aKiKEQ0hLfhc+FwdH/i1aou+adx6IMn+05wtcSTKX4qIiGqNs7lY+Re7T
864YjEKI9sgwh/v7F+CipDFxmmtjXqgGJ1HnC8NoTYco7MvBNy3AYwKNqFyGUCu2
EVReeRcp0VSRczKO3SLfSgRXUXY/6XfoMd8z6y4FSzUEqyrTfF+yqhAXcG5OtcwY
cDboxcsFTEcfWW+i7aAANF6MwvUjadoXvvNJzVsCfxPJlHTtfSIsarrKshPeAoAw
wwIhpz37FnXmOp5YEs5PdAD8fLG2YTRWmlvCpBaCxHUL7m9Om9mAuHmTBYgELhvg
XbVjm45mOJjYw67b+ux+Szj3NE4sHNrwffmaVVuZ82mhC2bilj9sywHHn+HP4XNZ
iCvK67mwGsZhvu6Yixb63uDdPjecpi7b2uF9DCL4UYt5BgDbrsVYMGXSTvUbrNaZ
oUdZFDKM1m1IbiEfpy601eRVIi1+H/WHsb02cVtuI/Baupz6VYyV/6F2i9pKtX/I
wv0UH/TI2bvSjTE40id6NB9XReGSZYFWNF8ZJZC2eccavs7A8LUU6awOMUlcoZoX
506zxAdB/gVxAhHqNux3jGa4SklV/fOkNmqEr8CqkZv17e4b3W8SsSyO0NHUIRTd
s8Uzvu7sjANNLzTi2ZTpXTEkWoilyLutowbLvp7sTpPUH8JpaEPvsTxxPr+sXrBa
lc4wVxUnfbLQvNPzxs6cVUAoiFdM9ngB8w7MnhIcGci7QMQMyvcEFEcxlyyVEJt0
8KzM6AglnSXoSODWDLWDP/feuZUhIbNsOoSbGgXVzcnLCpN5W9fG/i/JTp3xAPg2
brYrgfM6yVynF55EVYKmb7hGxpw0Z8Dd/AAgpjXqZyVHux+5n1WKD6o4VVLpnLrh
kHzmMrB91IWs1l+WSl2mG5LCiqcpn6aTKALGjuXUQCzVQh+MDK5/1V1R3Cfw4lZo
93Cu+Q6mz5jj1DEmnWgW7P2WvGPI1CQig5FhYstKxmH5khwotJVYesDs38kM0lh/
Xl4D8eQaPukKWzQv0sj46RNNPLwtGEmBGj2py5N4vWGnuqfb8JBn9Mn8F1HUYf4N
jthIHNvhB7PcFRlWgVtcTLGq3GHtUojMTu5bJ8SRGmIHMTSwku0BYyrPl6OQRmy1
GLfChCh4YbHbcnAC59++qVctSRunpdo50jDoT1S8E+mQODo03nyjZ29Sq+KxZbON
J5RtMookOS57zPnTZ1Elw+Ij9OF9RWtDp79M1B5vQpqxD4+DiCA6AjxfAcY5FJHC
jj4TKlQDCqUhUb4VI2YwZRNUi/XeMwZA95ECV2nYeCvvZesdKNPGlyZFpSReqiee
f73lYxm8egQtIoKvqZJRlCuwxhZm4lod+QsLdohdQM3xZvgOZsbOwkWp+edcZc1J
Pzjf7fRaum/8JeqGwBbSiYGfV8hHxqs3FwKhO1quwYyVJbUPjDGjnRoG8MgLxwAQ
YduR13Jxwk4xmY2ai4FXyKrHHz78QA07Fgkm8dJHqZ56u3L6PCBcOxq0Sx8DZTHj
gXjEw464uJTCB6HDpqXIu1GkarKAeHUkYbzsSumdd8F1E2yKOBJDtu73EUd3/wNb
Ari3f+42spLo8Tqrkfnb3e1SOI+usb6Fm5NMmoj7b3sLN3hrfG/K6zK7ZAfghuiB
Swk4FiJl+VeP9fHJ/HqAWfF39FQokbTOVGjcDHoupnvT3BBRdO9nVuaxSdwb5hqz
4MfTT2qmHHWJLelHX4LJPcuBa5RCYT9otDwHJEVsCY3MXJbbHxBeJzdmsRK/9Djs
WUh9mCvQjsR+LxOzSnOsrQTaY3oz2E/Z7YxqupdOUb1jHLx9A/pe/4nlli9MZkT3
DUSMeq5v6YIuX18DU5/fef644gKp3zIsAB/fm7zYdkCKTYJbrNZpsfDSeUjNUAAJ
a8vxUQDp3dyujSf6d0jSybYygtKcTHPBUshxwk1VJo86XsV+euAs/n8aGRL1Y7Lt
5XpmUCs3akxaUe/0uqlzaGQuwfq6UEOqy17g15Zm6m/VSjcmxKsskRPhTVdHx3RZ
HF2QFMRvhq6C806BJFXqJOi96IdEyjRWWA6LC+sH8tIyChGjhY2s7IQtectKrnpp
dc2kNgn0HUcopFDWth2yPaEsRNVQCV0a+4amyplCe7wPQsIUvTm7smKuJ9tXpKbA
JvT9h4fZF/Zhu7V1jqdEKFpSTmAolxhUyKCbCZe6xq+9gHuU2VitZ5eGaz8pcUhN
CnJyHlZFPh6e83srChNtcAfLsrjB+hyyFeBwh8h2+8GAGiV4EafDmo1d1Rrl1AOj
2w4U8WapE98+IRkUeVo5Ky+hNdF/DsvOtXRL7SaQ2mqmzMCEh74idZvjgTL7xSg/
RIepI0IqHR4J+vdK9oecURglTmEFC2VA7rJZbjtPeuPk2lOvKcW//3pjX4wzyqZ+
RUO2Yzkz957Sx88sXXkzEWHuXJWA4dwPSx+Hsu2irTEYLeHJHeH4bmHnNgFdvSQ+
Z8uAI/+CJ8osp8wnlXLS+/C50aVjIfBNVTYzt3s7ZRak7MXDZGLEPQOvWlaFBVxd
PTkkVTW782dSp1XFhwKboBAY6uLGI9qBlxbAdNzptOLM3Fd2nnAkIt5WqhfI4Tl9
+AtaNUFA3FOsWQ9eBn8vcS+yxgBK833volLYFvTLoqv7oqzWIWGUPObsxkuSMc0h
M16YWq92wvVRnmyKm4jT+sPejgW84CPVxyMVmfNvpwmeBaC8aJ1Kz+flhh/EbqaS
HoAU19Pqjr4iqGBYvWUWZAiIs4yjSbU9y4Gov5JyRWn43ZPc4XETgxs4dUkt7ENz
asQvnsT6s5gla874LHyc88iOUNK0s9MxGdXJVpqhVm8Oq8qF9q532iOGo46w+5DF
yZTDdgfAMWIV4eEhYehbFn5bf8PPFFULCjG2XxWJlae6/nd+6usz2gMId0b1E7bn
cfUigKCvdfaMplhDqtGznV+VjLqskaMYExMOw9fTx/QtO9cWHDo+XK7gzBteN4g7
kGphP26kysueRPiD3Zn93HTtURGarRsHVaAgzFyozJFXjGEiMi6tcwRhbszRsTGi
quQSPDoQHazoDxsn7TKcwdLgXav8il2JQ73eGRd8Vo5P9D6CeMT4dKJ6/S5FgX4n
trKrj5VE7P/C84k4bm0b2HgVR7SeyI7EAQo9BSdRswxobTS/bzWqSwgEatyaH4iE
i7kla027VybgnZ7fK2+dvOstgDiPihNpb1l5czvYahyWv/KPdl0x974aTxTshwSf
93ZApAw8lknotoUraK1JVE6dKGMFeVrk9jFYH960rKu7XA+TPFnQshuO0mGbGkeO
IbRXFQyVQGX3Js8vEM9PJ+7nNDQd53pwzgtvCpQc+DrrC7cI3uc3QrLBUPAkja3x
EuJFwNKxFRbRKPMjo7BaubdSlYPBVx1PTNUQfBYET99EeDyKtZg/XXDyEYfGs2e7
ydB/73mVS3VJOv8l4m+OYzKu318nzWkA0WyOyK81XEYQuGwpCVXWW4rcJTUFIY+n
4qG2MzyVKljgc3gMKBko+gwcq1LL+IV4fOi8GxEFRYI+KIE3677hqXDSH7LSXbat
Fb6tM5+BR5/RYPNAvxZyNe8HbnlQBoRBmtjNbFttreTWPlmipbzkMrAq56Nd0z5j
VREyuI0VBJ5Rk6TW8IXgU4qBew+gGSm1t+DgqTbloxvYHHX9YGi42Ob2b6FTVKOA
Jj2VGe6LUOKQEI9oi2v4lNkB2jrIy60pFwoi1YvE640YNM1CVOFnjgn6BNr3wOYA
KXOSnCQIQuh9cwect5QtX0qzTCrkwVi8bdZTuGMWPLGp5lHp9lCqYOwGD8Z/1XBA
fKo0NM7mYLwKW5t6W+c7iUZ5BlcekK8HTX9VbEd5ObNVHRuX4m9tZnkFxa4EH9wZ
y9VOPhPgrPg6cpdFJIEattJWzNmjPx3tOOg3ik3r93GQiQsbXNbfxnIE9vBhWwO2
cJNHmG+mLT069qRTy6wtghLMUxl0J3WzeDySOehFlmHvg0BpqG69Dqs4r20LmKfa
AtcWcMxQpAlx2FDOPC+q4y83ZK8ekbzvzgmRIKy7oEYZaU7s6HM++Ha2eBYs4X6M
y8Fva/vzYYt0JPJQT0Y79nTPjBuJv4RFZ2fS4ujaLIgdLQE2zUNVqJhi1QKiMM4s
VJNXnkhV3Vqfr9sb/wcrDl9YA2NMarmV/GNkRMecGNg6im00w7EmJQH359Q/iL2K
EvimCZXj9K6xYIdOVNirSlPU4qHCBHKYGoFVl6CPdTBBX/G3VJ/veugc4ifOuXEY
HZ7mPhcLnYXDRRcNuobS4AGY84+3CYzX+oDcSWVwkw9tMlaxiXh1OM19TQuL9qbm
VJJe7vuqrXoJa/tq7F32VjAXjW+oDU5DBqpOW/aiQTuSeKVGGieMowEOijwtOisD
70PQUHqRTJv/XCoXGCLvOHYQoLSe3MYUaTINR64nr/rNLJ2ZFoqILNDjoite3+Ku
LpgzEc0fKxXZNoAZ4R2WrqZtDAqBkd3C0SYsKxT5tsigSlGa91bjlqsNjbJtEZPv
bnR6dXINGiXGzRXhMxDXYu1SJ/aahmf+FOM5mjguVvmmUSCdaD2sN0c1ynB6RLE1
XoJ2+myPwxf2x8BGsbsVGe3WF7OSanLhvcXTQZjuv9UpSuF+nAyU/7E4G0mG5WeG
UKtYtXDe4dPTeOn6LaaxBiInenmd8EmABHbz5Dk63XX8zm1ts825W59p8V07nQON
WWKk+uI3+5AyrMEl8jkTULrJgojN0DFx5U/6arAbS2iS3p4/gCbPKYshIF1WLCeM
y0JnmEDFUODoxykDiy08pGzsr+5lULuq7kEFum84aEoxchwSuBXlDbdgWvNeUk+T
NLouHKJleo4XFDV7CW9F/XX7zaQkTjAjE4lNO6FQCQKl1bx04bqMsjD291wgKdKw
ZPwXZwRlqVsfCGDKUKqvv1yNUOZfxf/ZxeqJKuteQds8cuM9ih77/hqAbxY6baTI
f2ZPu4A4QriOkFQ8ZD9hXMuRRxcM1BYBgDS19zDfO+sHwHEwpVr6fcufUbqXrEOj
Sr2/Rz7CCA+86tpyUKgGdDyEylIxWGsa8gIiA6OSavy/YpyTe7yHTtsLngNHFuei
jPyrtKh9Y+zZU37wb9VfMYY95xSVSxR19OYfBKV3SBe+XgLLSX5qfLRmRRW/XqJc
7j4drdCTqYWAXCy5lJlEg8hxo2oOynxtj9QH3W+t5YJo2XFyoAzTytWJL13iy1Tk
4Wjsgrovc8WbEmk6uSCGHai77afUNfToiUJD2TCNq1LEYjswIuxQFPYWjkxs7xip
+cUnxXdeL3RPCyEmx6vTCBspfmus0beIwDW2PnNAhVpon9c08ryr4I3Z2jo5RAhI
pTR99jkzJU29k3AbtIHZS/ngA9tXmlQcfXVA+HSukKEdPz55dYyVmLdtEtyrqaeM
eprBKkogBh1nCQJ7DhjIQp9qLFGbTXpVBbINTmA9/rMk03v8iHCIfHEbibQ0HLaj
HUgnZWGywNQxJpi/4cMjqH9uNhW9u0zyErL8HOvLyknlQDw3GPo56gOxXwGe1ja2
fcyisczm9qvAnSIYVnxy3PzoxRenllLe4h6nlnBx22PMwBUmG3s8pfZDG7Lu7HKv
Ir7DhNRW+PAuq05oD8jjMwjocjJTui5YpuxNlhYdexiDP340rYXICKevumFJMd9m
3MwSwg6ccL2tAZ4ppIoYurYo6vRunwEqwBnD2ekQrVWAfZBxKs+zF/zzcplXM1Je
39HL2sHV2SwNwNRhc3cUUvk/5UtIk7sv0zLZaSdIBSGwmzOn0CIAdBtpJtN0nQos
3tI8lWnV/fgjGMV13vVSWYIj7hzQNKDw3zVsnI3d5HMJglsMUyRAQFe+18wFn/3F
AprElcQ9Pqki7+M1vqd1zp6rygmOq84JZF03YSeb5/4wpiMwo/bzaAypCJqJ3CK9
zxtZlVkoUtIXAOBlySNt0NBSgFnQ/6+AW88HjZafvBrDYCC3+a4N8hb9ukcH+IWs
qvFSVtRlpbIZiytRkF3IzgPrexDNABaUw90noUKjZ7+FGuc3n8H3ww37k4jKwPtJ
EOF8X/v/oV9dS2KT9CEQ+2LndKIsrYfPxAQjQpbxH85elXXUe+nDSp2KauO0F7FZ
gNsEzirAGEDp2cwR/ZdV9tpFiUxtl9AOc4yilonVCFFhgNLSSlVBFLZxHU7oNQu1
jikXPc61j10b3YdDPrsBz/tXgFdz7aL9miDNLSV1F1yEPlirnEBxIywZN6nO7KnM
8OLY/gy7tUbtaGxGf644cU51dfdPkRwBtYymfMdQLT/iUeNXen6dPw6D40lP2IB8
/Lcgra8VppZyzWm+IfSbszFr5PMDec4AtlPBu+6oqLaML5G8Oof385vaTEtMYXs8
yJGs8/o5FECe/qbZX0inhU4IBE1eomIQjI/DwWyRyAJ09044PVf6SosdTgGZIgY6
6t+ZnIEWZdK1JqPbwYSQTc4LpK4ErYncAxiREP9Zvf3y5V1GAP0ILEJkpCJG6lTS
jS0TI6npWr4BSfmHNKWGcX3GraEwaUcK5HkqpX94Di9M5pmrKKhEXHE4qQc6OTaA
VnMHcAp5tN/YEHUui4VO/BfSI5rM+HuRXFCtJWxMcgM7Qs147ND166mWCXLfB+dP
62dhfpwfVPX8CNLDU2JtOdgE6r+an8gmqIB9ItCLSbk7YwfKTGOVUCPq+V52O7Ql
kimNzmfpc57GCNuXNVmx8kbbhxmMJDoNDeQHIj/vnmL6wxGx5nBtfgCwo5fRq4r7
enh72UDoIpOme1hHDwe8eS6QGrpOqddpItmZRKQd1iAsPAmMAunCLKXFKJPljljv
QWEtEey5xaAHE86iSunZm/HZEkznFRmC9eKRxnDYxaymGPvECSJ24gvU2NU4YHNn
pzs9x1ZJnqkE5hev5Mmuqv0xwgIYTah7joY+/ZZ7apj4z1FPEQ50cawJlUtAaeI0
/GWqHxy0U2/nVSurbx1iKlAI6FwTihBcEX0EB1RwwBHZUYD2iKW6tL81jbqhvacg
UBH93LfO+XO3U+6OvlcARak6AeR7xacrqMjWcgRpmz5338va0rjDI7HwD/GM3EFw
H5kJaPVTeEREmwiATBuifZpwl1B0id7+diw95zzlTuvEB0NshCiqrHYXI9fMSLrW
LAdVXOQcgw23p2iBxLycw1muyYOZ4P20zXNok9M5fDIxz3Y5RIsbxWGcuvODtk+T
mRaT6tyU/+NZpkf6urwGmCBUuzBLGyOYoam9MbmLFwi5UkwopTVx81bbYaOOn2Em
Yb0LUoVplzPqFzAxJGYFc9C1smqaHkqPiwuYL7jY8iEuIqf/gzFuR3v6dSrOZdWc
r9R9pVqFwX/1L2Yy5kHWJGgOCrwe5YPLjE4gzcIa1F5klyyjoWoJCalQHb24mbs1
kObvLWGGQQt2cG2brAY/2B3ZdSfPl9UU9SfbgIf2kYLblvx8alebO18zUS8zykiL
pmICV6OKsyT9LtgEY98pSi1opM5HPe2RzC1gg/DW9TLQzlEXr/Wtzvaha+VBexIW
1xq31vKq8705CkdS21PSKXRHK9mbIDNSy4eSuv2XtQZmpEDilep+hSrT24YgnIF8
2YEBmlO8ZIezsYOl4sjh7ekE9DLT3ok4cS5fpfq5NNoGS2h9b86X8eycZYAkSP3D
laeKxre67rAQBRmMmhZ5RwD2PVzijk1ft+/PEHvZLGnAzXSPpdM/d2xdr54IVql4
ZDluaAO1TOz4Xe48ZVRKu4aWG59tybi+vxOd3B5ABFq7RnyJTsiR+q1IvQo6d+H+
QNwsruobv4AgL16xXWdz2+5QmFkLOQbscZ2Y3b9UqrV2m856U3kRasDJAXUl9iyf
VDnZ8at9/IfFt62Eul73SAbWnIw0MMBNY9lSSmfeaOywbuTiWlgA/rocLmmeIIdK
wUDp/cd9luZPdsf7SvKyESfPlYUp2xx6be/qXMrGJlsqPeeHMtGeKFDObH8qlqnS
k+g0x4huIztlMI5pukP+1U6mJAdVR5MobLLm2YDhz9rkpNUojOPYe+j8vxNEcUuU
Ha7EoLOby3ll60dDpW314JqjNSORjXjOWhwGIgDgeoVgxcH4vGuWCQrdRzyf6VTX
khAPGWZeCAVTLvl8msgIHMb6JfM0Mesaj60IJbS7baYDpz9PWNx2FR2qmKxCD/VA
VhsNWb+YxocRAcqQLa7SownQaxLH/fSb7imSa/9OEm1tdqHCUdlzq30eNPS+XUtw
/kmIUkSWenUtq30ClNU4Rw0PA3QGhP+3UTucT823rX4wy9bza5fJjZ57kWJ/uCse
cjtaouqpqnHY5Hzd738pFWQoETQeVaSGDKtZQHePwOYy0rSV3zBkPlKtcqG4l30n
fl5uBpUW7eIy5gXkPXDNl6eZGGS8i5PNs56dNyY8DLKLET7oekQeYGRLBiFmXY5K
E1mfU4wLLV7V6Wxs5jQwNGIl/7lqgNdHNNbz4UfSmixXc93NHXUC8LA9sz2VC0NG
YmiVS4JwdOdgW9yWV/lRQGrNSefTqSx4s8Uc+oMhy3rCr8GBlba6Czkfx7gK4BWu
8H5Q1jC+ov/e2iOQFYEADu0/e4/QGNdC5a68dUIWSEMFP7zJ1cE63jRkdSQzbTWO
mAtsP8KAP9VgtlN+4h2I4s286nB1XkZDUwroI1WT/RjummNd1MEGYaaiol7juuq+
R6ELHI84hyQa1ttW+LfDmQvecVnK0S5gAdY1IQSm+4Y9Ury4OYvr73xnIHkNcgKx
s1ydoq+WSNfdXBfM89P9FdMGIFqRfHKJ4oyNQiYDdLgvULwqAVTUqJVyYwobLmL9
VXrQp+hfnkWMwq1fpJOZiVWv/Y2RSa9qiFvUYkx22EHEmRR2ifRrjAUmLd8keMuN
kB9Rkq7Nlsqp96ffbyXF2HZNQLILQTqGzSPjNXEubypkHTC3l3wHisBt7BKW5t0l
Z0I2A78K9j5zpiroQUOKS79480RBKR3WCM1A/jYZ9ZBhprR+PNb6wx0v7gOJHO9I
BXj5Jj1lK6GbBqLSDRN+gMvKa7D7pCNIh4G4NeqgUA1VgzYRIoCUk/RUTnO/rRCl
oZklpiivWQNeCc/qNafUlHJyqYk5bggREpp7GwFfg5Kxlcuic4XjRyZD7xpKhwMW
7+XE/i45UI1PxCtcglzYsTr49MArxeEVOhjUxIuvIQzxGsuoDawf6eJTTohE5eDh
GBn0C6dPibJDEMaw+lVkhRaJb9pieFiYtUSUzI0KDvHmmRpLyWj4vn2NZRldJQIh
F5BZd8eeu/e9rlDRdEzxrsyjwAJGWDI9MEfKVBoNZ8UGoZE90TuumEZc3A6l7fBR
OU5HnQh8RMpOmTPYfy+hJoVz7ga20wpUNAyFxaxyDyQFOZ7Q8ELsrNyRJzSZw+cb
rl0I7EGU+69Wz8tYZrysVaIPKwYtXuU4/hqdZBCeqFe24zjvow+7KZdQuyHH4qy8
CB960f16xV/B7erUxI4eJBosCbrqahDfxqI0OnE6os7UbwBysiGix4iSn181lwd1
VCYIlHY011cRxb/vuLs7dvoqzjzNvXGEGDwbTDD/5cFfGNrnvxIE25IGS3uc89vu
vNWFRT5qgtWYL39Wtm8oOUhuSGS4ivH7gGN5iSJFup4NVd7oYwWQrDF3qtmH7p03
2CN+4q3BFVYr5nyYPhA7LvSbdgTS6ol+QQpGFbqpix4IbRmc/FRs4oRwEjb1G8L1
Fabycoe7BMXOZKYxH8trGqIIUIcUxreZXT8KwrPxjgudLP1TOiTm7RkQpbx7jrhE
YG6HrKY6/x4zKANPnsFrfWrTV9EC650il5ppsEK3+qkl7sxMAh/M/mG+ID0w9AgS
eirlifnrM/6O4LFTyfnsACu0/vBC6gtudSOoWd1AruP/VpiigTdCAqVQHefH+T1z
qy27Ayfkj+cuss+b7zUPlpBJUcCALWrz1XFs1QOQ8gXSZrFOjwLs6H/vk++5wFl3
U0fz6RVKMTQnErHg6RFpLa2ga04BI3x4i+o125jD7MJcZwDTySrJx3rjxOxBprBm
vUU/NakHvC18fvuELDrjjgkggVzuzCbBbQ4u1z1G0I353cy7nMhn37YC07gAsoX2
z7gGivzzTHrt9HeMMYuIku8mNSobdSC0DHbFJ1ZE4pqaFVNhugkZdlLLRVXW/3gU
AIeGe1xKIkkdKDgPlktjNhdFe7JsIJ0QhY8gdJcU+fj/1HiJg2Pr2IstSrIg29pW
CbC3lhx+CssSVYabhfgcAr3M6kv5oc8HSif5C7arerRElvF3Sy7rMjllJto7YH/Y
EFc1TbhxejyaX1VM0+cU0aCN1tNougVL3Cu5Cy17fMfIIfR6rhVFw4J/0vhuIhrK
ryLb+pOggVXJtXqeBHKDdJ3vbqPre+gwXtgWyAs73AtTbZPRmLWWOXPRzYIGbms+
KyAkAkoVvI9SWQ4dw6pe84XP7mJQTfwjI42Yr922uTkDh2JoN6LD/HMcHv6kt1/k
ybJqsGN5hagE9/Z4PWBLZZkzFSEBIjQ4JbexhhPm6+dNEuB6l2uKgofVhR9m1KBc
tdkdkwxU8uB6njj7G8orRtfxbYOoKflcQ9gnfv7qmHZSrbl+Sk6UiAMKdy2KckZI
fmCgS86DMJNQlPeyfF7M8raNW2w7Ay8Ucx/wsntX9JilYynWFyNOlqnJcjAcCfSu
RAZu0KEBCtOnsaiV7yATQuGXXnEiL6yjGV1+9FTe0q70DAtPvcbs1o2eEEAfTe9a
GpdbW+UZIi8yQWGMVzHMSe7aOjZGgXNGvq0MBPhuF2UIrpN10+9bM1pQFOdXrLeN
bhISceVYMILUUpSHiwpT/Mm2kBUPvecKdnhftTAYkBjI7jETf8kXK+/g2P200W5+
qgybWFKD95M/ezI2PdKFxOb9vnjPWHOcEVkth0RFTo8seywllbdeszeyuYOCxUTb
rfqQNgiE3caTQZ6q9YG7YixIzZPyT9EaWfjROuBRnAaVIqsE+t1JrZtjSCU0XhQh
DoigZDHEn7ggzSyl3Pa+bcmrTFGZGp63sVplgSXDXAvdkBT651RWUdSL4ZMg4eti
qV0p2vAHXcY6V7dpmb2v+LhjUX6j68k+Su7Eo4LKMKO9JS7p7h91ubPKRkoPJkj3
R3A9muzI1Nelai8rJGIUd88FPAkNb6hFB79zXoZCIWassMZZ8zJRGSPHuCHUVD8h
PLNO8TRSdL2ffjWUM0SObYeXk5Q0F/m0ITqunuSl4VQIMpbC1OJcLejp2NXT/xJv
5YSXs8pNEZ1A+ZJUDaN+W7eKqR+3IBPqPU9vewfmMdXjvc8UXAehUFcab4HY2bBy
pCTFFGh2fXUcqcb/Qy6p0HXyKjyRR1KUM3gj3swJDr6MWtITlIC5Z/EfR0DWPj+1
JeSGiIaHW86QwhfJUNMoQOwQHoR43Fnd92KzFDpggqtQKCUbJWkKYuVMJ4XzOS3i
TKBjgbjjVFWpDDrxC3EVH2OgWtiPdYtzL39ieEMvRSTtYCjeNs6lDnvxX4/AcEpD
Ae1+BWrzllInFO5gdKOy+sTQgEqkqFENAiH8bzHOFTKqF2kRkbIU5tpYP0ve0Feg
6ulZJiaLeQv3VK80pvRdHrbienU4Bz/1LfMayROW7Y+MvYgZed8DxgKbhE55GXCc
Mx5WU01IKKYWd1NgYyxhJTrZn7aenUf2GFXfeVESsVt+bLjWMxJNSOQwPBSuwIX8
R2ke8Gcz3aZ6JN9IFTRN+UviNyzBPlKKQRe3o2QunX4CsXRT+BXW+uiV3jGpGyU6
BvcUO+sxDZ718ibyk8FXPre3VWDKqJwXC4MBy+Az9BE05z7T+yTzLs8R3BOcDfvp
M7RiMGIPmgfP07MargSzsIL0XFuoYB5deJH9XeIoRZbV1mBUF5OxitbckvuAsNw5
zBNnz+xTbocGFtLTU/Y+k3SHxRJcY754DiZpaOzguarIlSBi+UEo3tMFR+QNJPbH
dsUpRYsqkD8vCT6BVX9Me4H4YAKkozXb26+/5YT7Pr4FySII0ZOj79UsrbUzEN3y
lrG510DntkqgmEYL+G7knU3mF3/NwdjwLpHfgtfx5w/1xbmFu6rmbclMt1jR7Sm4
RQ0Jb/ouirVJ6dCvE2gaxxu+6hTp1PsSFIzZLz+ePT0z94aUVJouKmMWxZPerO5/
CLuEIacdBqv6YFqSkzONF1uJiRtJuI1Xx5VJtrm4pOLuhpATgEr8ghECjnLkaIR/
P40UWpyv50aWF5fmQJui8EzDAp/BYI38i2DSCPV+waLtgW4m4J5/pnHRGaGBbB0V
DwG8b2gWwLFveoZKS0/ATwl4JDBNkhOTaxvRco+pgSdXuBlzPq0OdnK5OMf0I75u
dRbsGRG0GyWOJi/h+7MkVoqqFvM55snAWIM4XCDm8+UtCoC5CBqKss+wcq6Ki1fI
5QcHSLYLfOpkdm3GYLKsyQUnt+AqHLzJjvnbp5uSLAoePimFJx83Mnu/dUfm7GP8
fXpHnNmfwvAAThjEY87p42GOOwEdrmljChD9WsVXZFLjWEIHhOI3P0b5k4OV4cFN
p9aKKsFySYQWk63CjT4UNoe7KRmGtL6wJgxaKL/nktlWkpD3IrL09kz8V3aU4WVP
S/XlKuSZyugptoEcCkX9qYCr8Kzzcz+UXDSzYcV32vTDX476iV2nwjgrNQGvngft
ZtYsqICtqYOIdPDXdGz+zF0uHg6o6mAlAQap6UeEH8izRG5akE79V7l5ind0wFJs
Sol9TYP8tqYArmDrJ89M0ng39ZHic6Jdw0wJji2ZMXaFAS62emh/eg9hV2MkTFQ7
9TyoIc7RtH5tfR77ISBRg5/rCITlAlwOE8snqEPYjo+BarslRlnoXsgag1uiyf39
deEhUxfBMta1MW1IpJa/is+gHj1l3vGaub42PohsAJx26dc+HDmlgblw/ISh4pUY
kGaQ9jxraD+eoXec+SFOMn4ZZMHste1TIfejY3Zuo+JAvrl9hiyRSO6uQwxxbYhZ
vXhJln2d6HcBnDquvRUo9Xkvs/WEV3XQFU+PR+UDIBnA9uyTpXDtl6WUmrcC98b5
jLMluib5FD2ZOXFDVWB61pS9DZ2vDjGTgwTkyl2JKuTF/9nyvWW5Rkmb9toXYfTt
c/AEl2TXcjyameQTcGTCqxk0YmBDIQx/CEGUntbHfKg7ZzUmCl1L+0F2dfIMxYTj
cpVJ9QgWKAH/B4+puA1tlyjzzHHf2NAmtdNRDWvWj3hyFb47MDiFSDqPKfs6LX3x
ksoJzllslpPESL6WYl+VoyHuyJjwI96Zh5QW6j5pFVzsrFz3LgnwfCGpy8LOercr
jdNtTJWBJe/LYEeHM7kT0UneMumHoEOVaMxfcTFfMt9abvhkttGTXJMH+SiQNjrc
jXELaOsKsV9GeZY7Gk0wr0atU9pQGBkGstYZvfBidqY5N8BQdk6UWzGms0o59ypf
184jPn7aOJPHwcy1b45LWHYlev4pu/LTYnlTyFon0LCAyqNbr5qGpWYDjQBxLc5h
cteo3EQwXJXdR2Hhk5VeZhbgXhTnvzb5NmsaSaCSYF8/q7ENbV36rXY+vzlyIC0O
NWUASQL7b5CEQr5h3e4zM1FnpSzD1frMcVIBKa57KrMP8YkOcgcaHxLI9wnKPJ+B
a9s2jnEU+7m+8aQLk+9+DdyFdwLeeYOrULgnS/xUmgZf9wqUKRHyg5nU5N4BqnDZ
tMhqM463+KdhNlHkWuUiDvzjnsxKEVDpui6Iffqop8UNLsSq8+5lvb8RB3VOxDxQ
Lx8pbQUvFzogJyM2EI9ZpqtEiBrYGOyisDfzHo9AXLdgrLaxTCrm2nDYAq2cA+ut
kYIIFKvyipkYJ9W2jJOehs5apdfkH+/4u7+YB0pbOkdHY2Df4nPGMfIpP6BSCZVV
J8bkXhWlTRSggBQfKRfc2uRWRsW2ForQobk4vygd6ry9SZfPN2PTw2etSz9RwQ+t
sVhecOL3Pt+4wA3P0Ldu24hj1A3NGSVrjVpjmzWLpJ6mgyNF5xXIUQpEIcT/dfrK
p+XL/PL4SQiUcnQWWgFVMFbGzgFNfXMXed6SYfV6afatM/TiBfNJFOJa0qWkkSrn
fwRlRczTqZOTN6eOjcbh/JRfxlId0PluMu7vRy2ZdZAg/CAv29gfsxW3cwrW7qUE
nPbm1jkx3h39U+EPHOMQFpq1HKVr7kkW7Sd6jZxJFflmhviSYyhVModvdywiUjjS
r1K11whcgMPdVQrGkmBM6veAXn23J+wwP18VJq7PaopnbRtEKcih/dxS12GlAqWW
3NtJ44CIMY/gKO/OagixZ3v9RoledzrylufDLot0nrzQYBF6evC0FNQJvDvxqD8F
R5wQHXsp8/wNZdqlGB+dmEE1gUFv8PbJdxxvynX0dSoHZs2Mchtw/P3gkmrOhGMr
h3Ea1h7iUAa3fphANX+vDryNUmPfWdg1A8OdeIWLgN1dki26pQXizYG436tcj6si
I653jSjmxIDxZ5wafq7/rs5lI/A0BnDf/WrD7e+/AyU=
`pragma protect end_protected
