// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IaDPjSwCpjjiUZR3IblrcM21/W/LUP9THeFFzo9BSo/7PxKm9Q/70mXaWk/6dKFV
uX5vZQDclCoZbG/7pNkCbVqvMyeXN/xexJsZOzMtnqaGGnptKrILaxEF1JbIaxL4
YnyyuSs8XtZmz6fbJLycFcuPRkbtq2YQQCz5XPe4MkA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 177200)
xhetgxZzRzb0QhittowslMORKfrLgxEVRmwn0wEQwdYOLeOogRkSuA89SaOn2X/t
VUWdYfsaZbI2cqZGqGdmnXgfYhd0hP0+K+DncXSsmeXvv/0LUd9hZ04q0M8vbALP
tmix+vVz44/73ULmG7rpkhqoQXN+tp/hgIgNzSq8AdaByRyU/Z6b5LpIrJAtoQoL
Ttmy0UuwNbbuJU26fYJL3t1RYtMh8eVs2QZu3nXU3h1nIo51D6Uw9rbXDY7Scs2o
SvgC6HjQjySpyRRp3eqsBsDQR0wBTw20rTQtPSe5EdG5GKiabFgHc9iH0qtqavKV
sjQrK2L4KKCww9nl2DhIimzsPMiOEWJe777BXijIbVyTuj80VLl70ykPkd7Gw1hM
Lv9mq5MR7sPdqHTQQzwTCLu0mwa5bTP9lmu7tLOWnXhN782++d3n3OhDaS/BNLDb
PvjJJyiub0DSz3J79zbMgmFxf4acVKcSUATQHACgNDKki4iOAPodPHsRuB8j2BEy
cv7DqvVmMS+B3w09pdTvMpch4+nEB/FHTyYopnfGObr6/NGLCuoVdEZM111Knwtv
Zv08qTcJkAf0jSWEQ6hoFfqZVJuhrSo1jCeS+mcfPdL15TKsEAkyauaUOby+ypyp
0HaJycgdtCnm2zMJYwD9hj5ddAFZzTCJfhuwkokYcou0Def5mohZpZs6019+pEln
Yb/EBUiHI2U3ySBnwC3k+ZifevrxxWtnLEk8iEOwaBaYWYYyj8bwiEQa7QJd1HZS
RZCtrw4fAoNx6keH6o8/etwUTGJY7w4fA7TM5IRAalsa2fWJhPMnpxnm8VEv9zOo
3gCf8p9ptYt4wqHCn89DUSSCa0WNfVZd9I9u1ZUDepnyNFcXz6k4Jpf0rEnJvIPH
83hmNYnCi0jtfg6ZIeYal47uasefnRHrtHS7NqFftG8WtcHzfswA283BP4dmUAYF
LfxYbV7YwNmSfGx4klZxSLUsHlFvauzv19D3f4ztxU7y4hTd/DPuKRP0/ha0XJji
BPqxMARnwIBM5SrhtqO1YGxRgNPl//32zYcxVc8aUPDQ0ilxe1SregAnsSnipOEB
9WaMYr1mo/ZlkE4UISSU57NWWpXLZvTGbeeS5xRERxLp3uM1S+iavkWJT1v9TxV3
7FkDPHO5/G0MLZtMp0A9S0ytTXYiQcN9ABnYTaRL0zpj3Ejtnq6PBZ2k4Pq7IjRP
1ZaQEcka3sS49FxLRb97TR/mUyFPTv1yFTBo8Jl32Z3bqQG6NjE/y8Kc/n8UbxEE
8E5H2rP1Jwg4H3E9PVUllU+RmpciDPA8wg/Mt8mExm+jOKjg4GAL84hXjuWGUSw/
WJXTpeHrZWlKA73rD/U/eWcZjm/4WW8pPP1c7YGaX2rDr2bMliG3baQJ22PKcpzM
mDt4J9jC9ioJUT2N9UlqO1qxYQ5xytmFzkaoIf2cYHoU8xIxEe5f6OgDaFQeYxqr
MGB18UD3ho1PndDp5U2/7XyCEwC8P7r0QsPFxMlojDo7TDcqSGsMRCoZ610klZgL
3QXeT9R+chcaiay7KZ7M2x3T+MCVkXeFwJ3yXEo3jUL2jba6T/UpJkeSgpkpXM1t
w6rv1MBoOkUsIpVF2lTyqPsH0OWArkpTUI8ghMOEdGEq2eavOY5GxCAztUCJTIcQ
uUiDCgsmw4WjTqnEG3drJjxkXT1N6fIJn8pqmr8ruSIS407XH8UUSneLccpZeuxG
MY308aPUdchfd6EaKMJVCKEgO7QXOQDpwgCYyIRoiMXD6wdpDzUkCe1DNQt+cPiX
O01dtUYxrUI2Tz8lMcvyDAC9Obj/nqcF4afbL14sLjfLaBoOKB7oYi8v06JlM2lP
PkyiZ7q6oXJDot9lBcHmlb0VPvBATnhLvMC3gEUDK0H98HKXgVatdR+k36h2vYVJ
bPoITkF6kXx2Y5974SF7VlaQi7dDsE9za153rw53UTw6QzbVRhpaquwy1BCTsl9E
PrNNiQainIGvQBa+hhmhe1fs091dgKu5A9Kxl9rYQAoHu2dGkdfvimpKJofaNp4o
t9wpssPVCwlWEhK/AgRwYDvO0vBgLxEKAS0k5vvdqepAKLsl9uY17IvR0ZFWNjx6
3nA0b1NQ0eFnskzBfT0vvohq/BaEhxy6Fu6VaMTw7CoF+Ucn2xLeceqa7qLoJZBi
s9rwsAWte2rw5rSWMAveQ+y0PcqTbt5wCgC9JgQkc3yEcuHc35e8f0kSjsd7+VTW
BFDhV0r2xatRa5cumsabBg5HUIZr3ffCy2dZOvqsSUTUHP7qGzHtZDUMzp3XDLKS
X7dnXK6TSHkmkYKPaL9icM9yKq2iVZYNPNpUno8AukLD5GGr5da3D4njaDlysOmS
WhJt5iMh+nUmnrMmJIrmpRU8jWuEAhlbfIsxJK4AcjjkNHVVQTD86KauzzbOjB3p
KiPUd7fUtUAY1IqCHXaVXKBNMa1q/zdW/XRPNaGUaOe8KrhEWCveu+3XqcE2OKWb
loiTzenPBW0Pbedwn8vPDK5ho+74n8j2HhngTZkaBBrkm/AZvauQoEv26FXiWx5X
fF1ZsDL1zkp6hMsHNOA2sEI6hYXO7NHpzaoT2tfXvn0K4ZMTMw71MxKxZBJ9HkVP
VVGqYU9zbV502vWmPv4vYkPwmP+6FVhM26RQ7fY6T8RcvIa4xB5IMexU2viiTKnK
xo3URBif1azjaCEqfr8nS93CO78OPznCzIjPhOC1nEvPI1j1fG1ex/fHT2aARcbW
SfsBvCgvlqSAXya06lt40Yyq+re4gTd/y6ZRKgWmygcgbOksZAKAmUX/AlN+Dr8y
PeOImgnba/hxSWFrqaGNn0plQ2blOCFlYc0u0PJSEtX8M7b9wYkhWcSsxz/y/W9G
iKoe+Hfu/sGX1B1cHPTdlLv7VQlHGFVEkr+/uNCUpEoQkdj7JLeP1ZFszeD/0+MS
yRTj+EcxifRJJbZTzINK4ICDmsPgtaRkNBK22ymzCxwOl1EDEfGaMc9ZhJhawxrP
kYR1rj4m7Y2AW6DnaTeGSKi1HTQQIlMCrH683K3AaH/O8Eotal2k/lNnRUl46F2h
ESmmnljZx8x9MFGiA2YISSpjiD6N/G/iw2jUfgIFWWWY+GbUmUOK5ROh/yz6+fJT
i96GbdR0H3ILBGVLJ9+mtorgqQ86MyxOsmg/wxcgiheqsQIFXBXBn2xaLXPMgXpu
pkC4Ht6aM/fhN8X4z6RqBH2vxVGhFjdxU8O6btHwkwsOHl1Is49tp4uzMDW+CHga
2EO9K+bPQhogDNVo7QNC+mTbZJgdCl+mSsQESSHoD1nMRyfuXixgzDn1c4W4Hz4e
vazEti6gyoClIjwtDy93PakZMQlop9pW+2aWfbZK5pj1CR+tAfvQhyiVHVGYqzg8
vzBpQkDtxuSBHaEDr5ItUyr+59Dw+WjL2ATsdy1uId3zKmauCnis5GV9bsCP7aBc
MrvAd25qIfDyb4NChZaw6PwbUgu3NUXnyjeVc1diuTXxVWj15HKCCxFcjhea3zG5
JFUFKqOj9xjf+W66W19q1JX+bRNDSqGABV/d/vsbE5G2JXOrzSrRxYgmE8PhglCL
/BU7n5D8iaRyV3gs4WstsVNwCcjRqHeetYewn6ilruQ4mE5sUbfCT7BXX+Es4XCv
HsGatM1qKPAHmgd6o65wxyhH65tXwjFAyi/F+LbFhfr2vl09lZc0LgDm4YsmbUkA
sscnNRvuQz8PQEMZxzdnh313uo4u6RnsOV3wQchBAdStK5GfpDXYmVAqds/MCcy9
jatkuu0krOR/DCwoK9FjPwv7ngPu1M4MZdV2tVEonYx3o9cwXF5+nZ9h1dVSRAvr
CgtOOEvhN8DdpAH4TsnMe+l/ay/B/DfRrCyJxqr/3Dh4l0Z7fU+IfaEwx0jzorDL
Xc9tA2sqwj8ltgRIToAoAnfVHsSu26J4uUYyjXozJsiOmGsO5NuhsQp85FIGkILY
zPEoaom1jH6zRHkkQW2GGvXlFXXFGh5MtromCmLAJF/0FrtaUt/4/pyykRjkr3I2
5q8c71qB/eK/LWlYK+r9QBo8aYbWtHqkQ8EE8S7g6nEf4uYxn883E7CZ61WlD0z7
zwx45cFR9folxLd2M8uWTDxu31GzOUd1uWAuQ7LzlB0oTw15pSKNH3Y7go8U3zsk
6mOBOQibj1g/GNV1pQOxqIC7kEEpp4loxXpLbQlRUi9JFFSstBd4jEFYPNJa+j2U
jTsDMXW+Je5F2hPaN+JU4Zk9Uf+92Od91QrJuyT49zZFEo1Pm/nE5+wtP5RjU5E6
jkTfF1BweS/53Mi5Ev1oqZ14MZfmzk3Y6HSLNshlNNc2dxgvBigxg49OU6FhubOo
KQk4E+U4bG9GlnNM4KzmkPStgVWfmJConiY25zaxeQfLoqCR1z0JVUI6YNceCLTd
xDi6/NlqkJLQF+9xxXVKCoK7thlr+am6eUAGEilKKukvSREnzWWXHw4mFKe1En9R
jHmJLpjbUhMvdj0YFHsm585XumccXJUf8ct0S+j7UvbyanDi1e+YrmRc0a/Uu3za
nKW52MpquPog51iGCweXjVxwcYsd6ZX5OfarRh98JkRcJOD/cML+aAIta8p9xmY/
3HiZ17EN5AOxWZwQQSlsKHBJOvU2ei5E+HHlMhxhhvcntptOr7Tp+Bf2PhmYEdtG
vLlaor/F+zPwHwrQ7wEMspRroh00w1WoAlUA3bX6kQEtRW61WVABnm7axMAR6Shi
CFCmPGMIUPsjf2Zz2JNeuFgYWlaBrEjblioYfeeg6guaE5x4ocvdwzaJZD2/E7J1
y/6wOJMNEziMwNmZSoS4Ds6MZpuFgb4wUV/Wahj/7oBkODWoEvqRAL8VExOEunCG
x/2OTxfySG2IweVGtF3rIBjItnWx30WEMgN+/TNb+xx7FO21YGz4bj73VDZRzqpN
YG7TBMxR4M4//HDew6hAtDSxsSvNrVX+9NT86XSyRxGl62iQEn40Dl2nfxWBLMGK
IPDHCLQ6znqqYpRkxLa/NpJocM9D9yTcNVPQQsFCQ2Z5PXDBaHl1whYNhQR0R/TJ
5dnG/1vNTCAigryVhVJkBcKtCq6B/yubDdNB3BssHI34BPnilwX2ew+1S1ofsRn4
S+lPj8IGFpC2F6kswoVcX9IL1acu2aJq5vdMuIwNcIuo8vJ8XCANTZYUizhJHfdB
WUa10K/4G4vLJbKHFWDK3jcteQcOLDYGj7nMI580LCVuNcFJbIXuOaEllDOL7avO
1JEyfyDh9HQIvShr4UU3CD3gX7hGzFLb83tF09M6/znwacjj29uGGBWLdxzoepWT
fwowMiFEmJE+erkZOpozq63RZQjmvmi/UE94RtTf4iipH3ZS1yqagADNBsa809EE
eOOzNnpHhWADipBqd5uUTnXfcibsdwMhufW/KQfzffPHR35z+b4fyY6lUkKrVD3j
cwu9I2GOeBfS+ZAhJJYw4EnNDmLzAHPyOl8xAoR83swN3kiV97G8jhIHECoA00yI
h1SsEswbObw1IWbj619JKB0K5cyCJT5+bt0q9IFd8Y6mHFsQtHaB15ivfUPNtEEO
cPGUaMaFUZ5noh51hKd3fvu5Ewa2oBzULGqxSyRCIrTu2MttwviOCK7vygxR6QkB
9CwHXH3vt0L/YJ4SXeIWbyzCDU+h/wOotqpC2gdl83P6S28rh0BzCq9f5gE6zcZN
mCtjwZKJdPchzsK7X+L6JIak7slH8HXdjhUUOfUpF+tjVDpJLEP7ybAsMLWnrVoc
4M4VJVbit55XfKGqn8dpRdfopbQKwcuco8dsx8DsVD+f7PaO6lwkJEMI2LT05oUf
ZZX5noUGe5267iyyH/CdRNNKOpwEqZGE0cvrWjGYK9xA60QaLkN3f2BJ2PGPJ0i+
msDcvElbL54IgtUUkAC8nmzViY1jsjrqRug2fPNd7jgNMgz60coTgTxL5QVtCLGL
mqimiXxSSfivq6666I/hnE76ciQ4mamT1c3abh7xNzNOj6z7UosLKDJOu+C7nQox
SNS6+ZHOKAwJJwTbzxIKUGdHVuiAQB8HB0G5K5QOK1jgPWnQ00pqMwA6PWOJC22d
tcL0CQtkByFvAhMNRhCyMGY8zX7Q7w2dtR+oNM70FpLwiLPsuP6qWJX00eKrV99M
RX/HJtbYSl1abRvsjJ+qjysMgrpftVU1TvAbfp57MIqawMzNPYj2b4bwpHat/Com
/JTJGZXxvwDLP8qTI2mXon6W4cY2FTLUny3vzVa+Y5KVk7NIjUqwogGXuTsto5bt
eHfBKtLGOv4JknTyWPJHJ/p1s+XBNoG8lZ2fvlLMY4gEsiW8HkyvTQbNZ8/fzIOC
QioeaYrMJK5YpXT02af1UF4nL3qMckU3+mFHvSLyC6msUA+fbqgrfWb+p25fmatY
ZRDS4hfwhkjVkK78XWoeRx+azgL6rUJihTaCvIULInUMcftRC24mU6K/JzMwUI4b
MvaCKywz0Wo4Cv1VsRJOXHnHU9qy0NB/o6rap2DEfp2dnc+wNXMCsh64ZFWrrs4t
Bp+iuJqkgpf9F3yvM/ySqXXO2XhmOM2av5wKDk0nhVx7nEtk1d0JCbjj0dn+1Vt3
SQ0MzJWybbkpkEHtLaTtljCF2d6czWIy4H9g8eWpcEHxHKfQWS4v1wqGovOtn5TO
gAmrYTjGMO9QKCEk8FQ/cuBA79Zg7tgGI+z98MS+Xe1SpP66uwsjCKwg4rRH5wlq
z84tXn3yXjGyeZmTMc93wpHzkIjfty8GKjgw/3iq7YkdXnBbsqo/Kq6RXl3/anjy
VuNS7DUWTNnTOKQ4PnqaBgksr2P6Ih1796QnkQSuX0/loNsLHXBN2ojDGOYHA8vP
Om5NpGcDEyChcOPvpoXuiHsuYlNdj7W5bSkgOVzFGedcdvjJ0CvmUVmAOQ7OwQF7
9h9d0YfdlXFs0UM1CJgZj5Q8g/FWzO/TALbed098qCeMQdKZWJEqp5LOEIa5o2w+
/RWx8SrQU2JMR+Z5N8QqG9hxxY/FTVUp5bHw+BHXOO6fp2hC+Giw2Mesizz873xY
v8YhL3Yk1+QFgwdodwWhLAA9LbWFsRkdVrTGMdBLi6kvImFwcrc+qtFtZgGk80fZ
2INkgR2cUUpdPxLBrskFJDHk6ZTRv8x4/EY/bJVxiPgmZ10clrI0fBw6SxcTfXoK
1eCWFmyUTvU3xzS7osysMyIMfloGzWdN4RtdFO5cwGiGbRsxqve3UY61kmHBvZbb
ecO8tGFdcv3M2SpmGT7iCMBVagT6AVG4AOg+gbNcH+LvQedn6LnfggEIOk5asgcZ
tyUMWTphl3XP3OTUPTlu73ehjKzRPnW6hi+wnCIEp/xOLt+bvWlK9UVjhdUFAdmB
YMQZwIxWvNBfTRvC4qWgs4RPNhhE5KJQLzkqj3SOmtddiXSfh2MwXVoPLjlcV8/R
zjL4GAc5jSNoVRRizcW1rhDS2APjTRoiTQ2ZJ9+13XfN5RNrhxSbj/EkLku22WhJ
OUqh61vZyIHmOKSRNjc/p3rJ4skMxn92vH3T1aON/D8JdUOQMIIEQweX3xZxIP0N
nFfw3XhZd3N0WwmdxvkS8uG9VJGhB5vAu3fmWIpKWSIoRhDbXsMBYINslfLBXCaW
FStmRloj7kuiozrbgpQ3S3pFempaOkZBBpgrTTjpPvPpQz2+nmgMAoC0PFTkQMPR
ik0Ia/luUt3V1D0mZJY4A1X6hPLVHfp4PC7XzA5To3PC+uSbN6tPmYbWNmuB4m46
QWtYWXWs95dvdncvyiMTV/nc3IKmuH6on2ZP5cmnFOifKys54y9EFuOnH5150AkF
bgwnTVMIyM73oTdyEgjfTI5JdhjTK1kJoDEWAqwkE0C4ETEwGRBnQ4cat3PRMWW2
a7MpODV5SFrIwDbb1I/miVDiTwXqwQZW8laphItfs2KtgDAz6voHLlVBdmAY/EDQ
cwge5JVVOjiBzGT4ijmbJjq4sjTsmrfrMJfL0Cu04D0uMajVy4pKdtcW17LAiTr/
BRVr1TpJndDlHrQDXusf24YQLx65SG0z88xbwym3lS8AcMJ8pp0Hefe969Eomgty
jZHs4hxyqtUZ/PkQ5js2vG55NEyTsW4DM+bGBYIm0e09azqjjrl+kPJAYagrXqbf
zrGHnJAuIM1n+9j8UmL4j0J31pEM54j2VC1qdbOgIomvd3wst/tJ7sZH/d3xxBvs
gjaox9MtpyuWVIoaJkxgYhjBaqZ0Yh4q1XquqcOAukiu1kmsd5ZQXJBKpZf9l6G5
HsMBQ0KryDq5Lt+eVMaqUSU3cbqNRczh8qe67tB3AeZ/fkzALfqWm5bJlzYDE+xW
Oo96PgOBND8h/ASmuo+tVGBvd0U+YV7Pca1lHbqXsA3ksnoAlGudGl7v+xKbO8VQ
RUzDQB2c6DaiynKy+YTGTmRjW2Ypk2VfiVq4IUwYSY4/71Vg72QljxqGdrUidffv
RMkfo0+UX+FTxlbRSN1wxEuJLOHk9Tu7Wmid62nCCnnJASCT7y4WeCswBvqlJjWU
oDDodAy2/1/Xr99vPMRO03P4N4k5oLAOSypE1Og0RSKBSTRxj66pCiO8wdmUrb5P
byJPNYuqs8rX82Y686QqPxqOWSHXGZBsJrAotxn/0S5De7UeRcNWvxZBVlkkywjj
LkUCAKGbmE1ZubU0gcBaJI3X8Pv6l0hP6xvO4v4vZKDOrpz6ZU/iwcXx1UYl9VLn
ZI//5b2sVDJ5/g6EYp7zAj/wXE192ErDUcOWfBfk5HkVUn42qdM4WzqCisYEfxx7
jU5CzawajEo6cFJkI4NDhwzwBdrfcylocwE8KT3tFfglkYMRntv5ZwsRo5F7PegK
uKo6dPLTepo64PaqLdwH+/MMp3JWeYTamw9JK8EPU3m6WHzCUKDqfF/zFC+ALX3g
sGe10fEd5Rg/DV6eDIqsEmnZKSIAWF7PjCczQ8F8MnLWDM7a8mbJ7rXPNLMQvLsF
TQ/bU8LNYN9fHlbFrPZO7zjc6Z4l2GE0t9ZiQorPBgVZp/3dQlD+X8WFlE3LScJF
hR0Yqt3ZYEnnDdac859dmyx/JEbMiHR72//ZMP1el/Nf68A13tF/TpneEpoC5OOP
MJ6VldLFi8jvfKRO7dQzdBwCXSUThoe3ORUHTEKcpD+zrLicx1F5ztqmqRvsQ4Xg
8eMubrIrRBWU1zqzxlLD5DOHhAwTE0kd60e08MNM3lwnJyI9gPHAj4eIiaMywQ4w
336W0VJnW7Tuvx01NBCIupOhOoXzXQzppXd4AcRCDJYK7QK2PI9Awnxo3kn2PYHB
Lp723hUejfajYMhtMiV6xPESYOTLjmjgl1zkZC17pqB2JvJJd/aiHCrtDPEeMl2J
lZNKJPRppkVLJFb9kt7ETYWPUGuaZROo+77N9lNjSed861ZhVjKkyuN9KquzimVO
sdxDOzc7MgKvX1TXxIouNrScvvpekD5kK/R7zEa3KmZNSTB0HVledAogdY+R9P5w
RD4tS8jVnLvlKF9qt8zJ8IN+QryvKalluhvWroySL1uN5xPEEBSLdDm79vTKNUjI
ExDew/dfj/luysXkzWlIrf1TCWgEhAWmQE9KGOZC2d3lw1kLdl56QLYXjyqDvn5l
Ny/mYwebOr/Al66vRdSz1ggmia9aUbsr8lDoJMgiMXAegv5ooe93Us3rInBlzyy8
dkR//sosnKy9TeLwbHYnQ67xZEcEsHooGYFe+e5Rld66Cz5bNEh6XL7f6Yx/CyMz
8hs8VNpeYmAagp0skcl54sNK144Yj3liSs3Wbmy6krVTd2TSnLgaIxwfUVtr9unO
OP2BPYrbO2G1VZLQ/y1vLaVkQaciQDWrlXkGtFn69imIg36BPyhSDaWgr6oyHUk0
If09KcXcfrudL2tj8aTZCjjookKfMjB8eX7sod/JxxETcqZqMtiL89Jzux1kich2
jUOoL4/ioYbBrZXIR71x8jPdnjgVpWGPKTd+lYwoZgg8eISO5CRfpHqt38IbsXB2
AFihZXZKMVOSf767XyiiECjEghsvFHma3zz0wuVCp3egHstQb7+BTBE7PH0dOPc5
n3bqHlXQiwXTbnqRfv6sbfYC5B83urbuWI3u4TZ9tXj0YVi2P5wmzH/8Qlp/WCGB
FFjy1n5TtmESVDmRJ2NkpbLYBaVXEm4BGY+MV4LJ4FoOaDUf3Cra7hID459FjIOA
uTO0hFIKgihNr0hWrdYCEmIXs3nX9bG+FmGN2aZeBxzYl1u+rtCrrFR4U17JgK7M
r2z4VD0mINe0nVxX7ptDc8m5QIIZAsVdJkzXqbsZL/SjWHXfkGw9v85CxGzxCGjj
+aPS3kQQlklf3R1zB9KXIGZ38hWPb0D5RcCS4REVjwIRpRtNfyuoznPTY6CSXpxG
yh+ILQBMH+9MqByQ6ScedpfP72YM0G6la1LIeyLS28+k88qjw2WyQn/rwIeLEIHo
34+1pP+9yl82SVjeRmeBdOHok4uKsWg1cOBIJx6glbB/3xRUV8BY4laMMlf4jHPP
UeAEgooPyJRVjHojfpN/WLacFArMqnq8zWIy7Zm+B/IrqfmbiTnlwixNwwPKabcd
lZ9wMvH5MHV8lQnaBreIntEQJjejM3HXFrsiClUP9KaQ4yt/anpnpU64LzLmoVQ4
sXt6psXnBB1xlEWORzcOaPYQ5dXTx+bL7PcqjSSgjFj5ko50gesZxhJ2tJN/yMT+
YlY7BNKGkT3T1RldoXtdxmnbRckWa/Ng73SDx5zg9ewBRLEaWbERfY6lOH2d4mDR
3Tkov/o0LZaA+TzyiLhFyhP8IZpv4lfjk6Ts32F04FRISBD/ICpDZifRTvOsvQAQ
EH5f7Wt4IpqMZy6760W3FMi158M12MuL25bQpAbeT5GXTRpdpdVbbm52+x8HxieY
eLYCQ47EQRDWOBnQJK9gooSRqXEYuQYoZAF8yvts/iHvIYsO3faOHgEQZbrs2zGk
VLEruM+OsbJDGBnd61GmoCRxS1Ml3dVeTTVXV9SwMU1hatmfFx8qDTO7l1G80x+p
0tEHHf/5tT+riNXembz/p6AJDdjNGvlzP9AMI9MaWhxGthOswHzL1YqTSo+R5RmY
HNDvDlsCnN6GyybASIHVdfssGBfAgpywlIcVFCzJ03HlcnQz6QzMRohz8xJIYj+g
Y+Df1UD7IQXR4lHwUMN1oqCkKuQ/d9hom4fC1Ko5GRolAMEKe88hgvSNpYQwKFMU
cA4TPnquKEPSyF8juT8Wh9mVc2reNNpwj6AS4zxpt13b8i9A8mMEyQPgmghpYXas
MFavrQutFFffbz2PFXy97Pd9ozwc4UTEXBUIAfxT6seYfUXTMUWvLT4Wv4A2fQxR
HD9PVGe5o2IIKcdunleICcfOdhcRU4Mi2zJF+f6LtTrOGVH8sKB7vLLb491evvDA
Kyo1HfnOF7/AzVDchR9Xqks9g3/HH+Q7dbZn/tjvRYvc8u2992/3NWRO8YfyWndk
r4wnQQC2SOdc6QHyGDxh6SP805py2E88y0tZMgd+tLSvJyRRVio65TfGtBqGF2Pl
9UVMWMlXabmar8DxldTsMaml9VfxTaH32VdLzC0MRc4X3jbj2d74C/q6Msbisqc7
gjS/T21/FHLyrlPAZBzmi/Mciby6DorkxnnXQn9kmHfIiQkRGtKUMK7s8H7l2RNN
zdBIUGUNiwqKH7i3pREbEJReJaVyCBuzfR7Zfx1qF6Vw4oG1wbdDNmegVH5t5cNm
sPY9NZ0CFEsDOnHYVGBBbvVeaTG4cR8ahoYZFQjWVU7V4LMXivkg3EHFiGXSRySt
wdLuXMvPsiDFUdJQIt5QmEqtlJB1eTF2RqSCwNYKb8Mu9wKfpjRXl9uIL3AOMDwW
FVUOYZbD7EToJbxWPUtl2TEEf1ZGZVXOyKWWO8wlK9B/YmPggJzNSYpPalfW4Vaf
5zxbqK/b7OISyJXBigI6W5beWGj0eUSuPF91DSirTZbqXEv/XiCCQvwTOSiFxSFh
d/bE4lKgEk+qjsy02zaO9231yPvyMpUgmMZbCym1vyHu4d1Px5oe64QxVZFeV0//
ulh5+ryEcpLZfMzSoJ0WyZjmNYpKGNCuRr8r1FpYkE8dXyGy3cR7cb0SNl+K4x2V
rXQXv1L4tlHiySFULj+ZgY8mVivT+Hfh1m3lk7qfFWzw4DufJc5MPyWZ9EW8GJXs
GLzXDJ2POWuFUg74Vxp4ykAEZSnxMnr1ZEIJMlbekmljTl/zsECi31QhZD1uF0vM
DVKR8+4mHvQAPPW8af4DmY/wkejy2wLtAqly/GDsx14En5GIScva+V7Hu4Hjb7oO
NwwZtDj9xBPuWfiyNF+X/7a4tAorAA5fhjc0gMAJgZtwXtE9ZYm/48/D3kSrtQWw
lga+Q41+oD2V8HH0CN0ElPZklUrZE7GkO0+d1dBs9NFyxl3MldS5iR92hrYptoQI
8cBwK8zaakdOtp+gUo1Sts4t300QY7a4LzEfgdtRSznbyod9Pzy6Jv7VAGRXHd5n
79asCzZJ2gMsJN6UFNNBWeVCFggjgYqi5CuVLg7CNdok8e8YpU/Y5RPwSotrokMT
Wzp8jXcllTejuLLFun39CPDrlX08zwqaNrDTcFN7yUVz7xV+gE/eDznpah/sUGv8
SAp1kEp7Wq6D8vtUStVJRPaVFjIuCSV5aulPgyg8qJ4YJHRtFiJVyXMRNO5PhDf5
V+go2q66TSSiEhDAela4FOLUkLV7tK9x64dywWUsSo/TtsojnVY9t6Jqh4A/t4ZN
mf2INnlUY3qwne3wFEOeP1DlUy2QBNTXWRqud3hfJoEI9ymO7rVqUvNj3HsnbHB1
IaJ355qTsYn1og67hMhngBoWBnZqDlnI4XenRr6MmqGhr5UBCfM0ezHYcgHu1L80
6/1hedZD5ESsESzFmCEcvcfxQNna+kYHr80k6Q+lUVZEVgt3hd69QA4TO/lPVNys
EdVoAHadfX1UcwMmcEraDIx0l+DR1HG6wa0CIMbnJ+ARfrDSHI7cXWw4YF6KHQgm
VD5zOqQzg89GGln2bH+dzcRnqE+DvPAQWO5YRYl50Y+TzlZsvyVQhNiLuyLos8Lm
b5fqZKddDOYEbfxUW+9AzC4SDAFnyzIoSxofmxe4vXgeq7JyP5IIFUzkKu9WXhEj
lr1ZX10vZsefX6TOhPtIUKAwp5vytHAWO7wqX2PA3/qoS2t4LEBnoZl7dvAdEtFC
xhIFkm2DzGojFAkIXk2oVdLXjfkAe02AV+pr5cpJ3yQGESBN5CtkFPdFY7p3LN3A
gX9SbtjJWMdaO4TfP3w+J0Vqh7gjpv0X4DNCtUVWR2VxHTFsrKGFnd8V3VQQm6EO
5A/+J4FatL77aWKU+ilBejuuHrqCnvS+sQEbDpz+jX+dnKnX2sUw2DiMM4Pqv1wx
NPyFUM457F+CwYXmHqPB8gqXY1pU5Lls0pW6KbI3/1NY5UYapi1407jhrCB7RtL8
L28QO8s1uDoOVJCH1qHXoJx1Dwh66vdyuPDogycg6Xrqn0W/iWJHfkm/o4cAytHv
5yv0mjaZ7X8VgmoUPtKfPgVkGzFEAkDlLk3wuXtjBQVKMbMn2CipqUQi+/SwGiUl
oWq66M0VLtTZoC1pjCUhI0xwZXCbq/sbItGA6i71Iw/RjTGt/M9ub1Gl4Kl87eiO
wyUAUVxpFwuuiH7z45XzUbE4iUB76Qz8EOAsoY0TeXKacw3pJ5SolnTaFv2xASys
OA9W4bW/7AjQKyOU9RW6KdgX86s6FydQApYrlnOrTB7BwCI8Ci65bL2BKLUnyNov
KSzZcqM2FM2bT+0i3RdNCfw6ubA6MoxU+qQJhyYno0luL4Dbc7rWE9SoC0YW6Pi3
ruvl8/b72jIjspmuQ3nlZV0LhmTHVvKeEfxqanqpt1riPSWgkcWskC0/BCC1oNkd
+NhcBd20iuYtwL/0srE218cBKpeQbyYPWnawg9iLil5RN5xSCJasxf07dAO9081m
uyVuzGQZ/q61N4XloOl3JAdlVzUSVs45lF/a6ugKzVKMCSDQhqw+j2Vo2T+gYoOK
xDcfnE4D1xZFl6Uuk763nN4bg30HLB3HiyZD1JOM9JxfVyBoj5RfH5iSUEmf/vmr
VsjEN/uCrc/8/R93xWW46vTgNOf9zajuDw1vXT2qMhDQ8sSBJloTz6QTfdmoWoVA
BOtEJj3vMUY/Hw7pmCGqv5r8Bju/+zqv+WQu9r4F7OyEfBZOeMfJAuOT7V6aFt9r
cQVnxjXzNaOII32kP+n0u0CLKXaNQQhIAGumKCE7jBX9yIXSPJNxHs3zFOTXs4pN
kBdE8p41ncIOE9g34nZdFvzY12PkLzSSkSlSs3x/26BORJl1EqY6M2kVHStK/t/s
PfbHDCACdyVjhl06ioliZBQ7g3ve2ChIAwpkwCIwf5uttjK94tXF/T2fSiG81A5n
0pYK13m4PyBoxuNTOXagdf8S/lbo4icH9jNipJuhSA+tMhh3AQGJrLp1raRDz/Fh
RWARLWX79Jq60rAssf2Ue0D0TbWmhzxLmkJWY+AokfWRLC1ZDNSU34AIBaW6lcMG
S0Io6Q9zWlYEd3BcMnBlice/aQ1cH1bX3D5P22UBOEdNQp+VhXA7QGjhDBLUhdey
NWEfqoMAEEl/SrQFopCN1N9AqEiaZaTSO3Yxtye1oBcWoZ/u2+TXemNrDPaCkBNN
e7KMMnB5gECFgwfDmOZ0VZJL3W0uPwLDrBF5qWTcz4baQ5x/QDk+NryOr0xfk47i
vxsCB0fcWyxl1aP1rQeALTSrhE/EGZtziNaaltQXNqGRYluAOWV+CR0ua7n/5LHO
owGgfvaQ7xlnol1YDBCHLgH69Md6NwD1XcqotAtjv9HelGyK9T8zvQPokHiqq32S
n5Ei26YlYHLNP+OOeu2Zck1zhqAw+2BD1GgE9jAtHTcuc1kfPqCXWc7CBQf00h5Z
l47DI2483y5Tm+aI+tJUjFTP5BMjsFL81H9Inxu5O+UdWkrb7hkoaACKMTaLFSjD
B/E6s3CqNEzx5cl4CrbCayJX0ePpanmcxHTNcNsaFYH5I0E944S2s0hZvcf2HOG7
bp6kCkRoVBK9dMUVWResOwV9ypOdC+MUCuHzRks843k0iXQ0bzEjdvO940dB4CUV
8g0FjwQIDgZoegDwJIt/gQiL5Fe96MIej7d4gGysHpeCY+IcMODNcDFYJAnLlwCm
ujSRGyccCHknFQ6q/izrRIkD7ooGTPKCNdcFSkiVXJW5RR/unxF8NzX8/H27uk0z
fkxdPmBVxaxacUF7RfEZ9HRVqehhQdARr7bORY+wytvID7uPVZjuxTjKCdC1MtXU
7UFmdUgqGvhHq6n8mRl995UvmS4IDlZ46otpLhYz9mZcgKY92EdMatubPqNxcI0H
ZLQPQ/D2RRk9tBpr27JAA++NPDvaTQALfSPXFVq8gbRAODVEhzSRask1oejxM7WV
vOQHL4u4tYFiWmYDmViu8rxLcfCVeXaPKNawVi4moWZ+3F22a5O9I7JhZiIfVk9n
IrxnkkMjnUKWQQEApQH4/M43qCYKbIEb/ZkXZd0cBSv4s17/srMKNeW1u85oE65P
tSSLo8k3ZS5RQ1L+Atvi7qHlaBjIVydic/uOrgl58MVng8LCUozMUicW6WhdIzri
yfmSthZHKBNdsd2CvDOfmb38an767lqWWE7ngD0WYsuXufZH2yj51lU3EwPTPVwb
RC6K5LzjOayinHEJ6h34n+mNC0Z50aaJN6jVUFAc2/OJHCdodCO7ZOF+8VdbqPZV
BEYtFB7WQTSpi3cGxqiTfh3cFfeE9190BOX0Lq3jmks9whOJW4Cdf9M6DKGYARYq
453sUhVzB2++xR5dk1W4pixKSG8/429x7FJgzTBbg92hlRKf3PxDHCixOYmxCPU9
SYv1LakR8+z5SSl9f2Qnj1R59TrqSZTobw5QbG6peoyPTVIvpHuCfnajrAT470NJ
umQURHTrDslzU+jUhi87oeq7GXcNBwB8iguEPEj7jZ/d8IEfdcg02Aar0TAVAb4c
j3wCKOkxW8EAB0x/yutzULBmbonrSId106J89wA44T7lJA+r4dfrTB3SwiGkXJ8x
7bNraDG8ex1k8DzgmSUWM2RSlKWf6D6KyPXQwj3R+uAcFsNnG3bWVXlsu+1lUoZr
b177hKfWJ+P7JcGIrM3QRGo0dbMzHuz9d71RYHRd0M2ifzVpu8YV4KYRP2OeNA+a
c7mbd8M5jssfTbbHHRX3E4ewQAsxEdzPjlDIw/IRWWnNZrewJNiEj7x+JPfLqYGg
p9b+tWGTkvgRCDi3D3OCcRSK7yrIRPwNIpSi0oKiBygmpNgR+V/PsAxwf8hB/F9V
BGPprAC3/M+knJGE66T7r49wFgYg2jq+Ezd4jAq5wnGJUOyCIXKnhPeRnmCVnVUN
ORASHB/SO7NZ9A29CxtJssX1/jlG/x4pUovpcpHECv9CSIzrPXl2KzuCWEyXD9Yj
p0UfZIlb9m3hQNQe8y0nHLHO3nNX+n81RSp4muEC8l+ClfR4mt1ECD+ItQps8znT
xNf/qxRllmqCSFzdVGbnE64byGHXBGZmHYnNn2DSf/FE8GgvyyBd9I/5PJKx0gnS
HU0rgwH5Up+muRQOg1dtKMT4ywwqKaaOUHfvuME9IA5ySieQDvxHhU3UQ5++Bxfm
VuqCSVUiApPpA4iqNkp1/RUScd/ZmTm1OmOIUWs6qshh4aMGEGdbNikELjvM01sP
wNZ2bwxhqOsETNORL8I59Zd1kpJpZ6RkoOheLvHVJLqlP+Te7rTZWEGW8r4RvNZ/
6L/M9jpRlRkjpIjzqX3mdzmNSWCD3oXP4+t46E16Jdf72cYuA2Z/ZEr22OtAZFuM
FCIf63qttcv7h9s6I/37M8BtjJ1f7vq9WhjI52IlyrHXOUH4lg9vSkTtxJmSjp+n
LayLV+IRSmZkKi+R/R4bBt3fhT8pylqdx49dx9fd425R43C5zEgAOhKwAE+zgc2v
xAtpssQp5lyPFq0YjjWcii+3HSaUpJySYOL+SjNjhc35T3YR8Ti18tLt/eqePrYo
C77BV2Anp464VouL1rS4JLbLGQ6euMdzPJWVlhbWSiE0udAiFOZhZZ3MjWRAodRq
Qx3LZoZZh38jyt6v9x8KHNziDpJJXPtAAQ2uqVRQTazoiVCdxiOYPiYWETELVqxM
F8XLW1qbHsGdNbssS8MbrLdU2E/Aq5lqAhmEDPSN8hoCdg8kVN+z2e2EeDuU2IMI
PZHsViqCPPHKaUtD6tnT/tF/I8UqxEfeAdiKlSoWBajVBloT9lCHHd56/VBqDRQH
F9rqASEad57G7HI5gl232VqPw+BiJf+FypNksvOeuJ9CW09baBHUJHENzmya++se
7+2wbIGdrEQ6JhMmjC+UZOW5xZImDqJJ4oSa9Y6X2GndZXTyZZzXbrosw4xIMEyZ
SPlexfkG1A1hvzNnu/3yrUgE5QeSrMWmmgH5ch+UKlZu2XaBdJYwp5nCY0ydWGDO
NkGC34oAHXeBT2CeOhPcyiJ83aQ6p0rW0I2yVWRoETbtt9pgR5qUJxZpjGIcnaAj
4Kldb34GCj7QCm7vPp+RB/i5zFv2hUTCzoDJhi++Ej4L8nA00vzK3rVjN9QoclBQ
U/nBXZaw+FJEbEspO4UQ2jf1flMtdRP7wj0WeySkP3mO/daytnPQ7G7lKwZPLRCm
nc0jg3i7fxe8zFeggEcMl9ZQ3XQdn7MD6DfGaJAfy2ovRw6D8dgtAGgBsv7LfoEy
qbhdCplw+z9moBkoJ/QoeVSLeWJ/0XrG3ZHKjj8+4hE6jYtaYhSP9/Zy45VOFzx3
q0ycRTauzuHu10tKy9kH9ZV4OYJoal1rTo2yWycnjxsc1mSq2ruHlie3FzYQq3/r
GA6SLFXgo6SZQnFgXn6mHy6g4/0U4SzhBP/A8OEkGhznUNGtP1hlf8yb0PIiPnQR
U7fHt6WKVELNfhqKvsPtBcvLxKcUBWglCSVZmWz81G2IOU2dkk6eeHQlk85emwfQ
08wslSOoKrZ36VAk6R5nPfHSPxFEwzUwDQ55dJm+N+XOP/b0dq30l9p+fCePbevw
dtMk+X+gZWitkQCor7BtFFJhmAn6o2pkca89TvK3cnaSnB6KSNqT9oKozFqV4CZ7
gGsUun5xZryJFRVm3xLNFZOPUhSqu/ANFobVCu+0pEh46bYmucHwceLk4v+mvs7c
HNTiGg9qIskMwbs/ZSjtACdMutak96H3pV9lqv+1dNMj7coKaCJyFy4iL6LFp3VY
eez/F3ySy0vQeo80Momd0BW6gMdZGeVLVVnm9/XifHvD/yDC0gZA+03KXU1adF3k
XhnNW+4MwmNDS8iZ1SkAAy8fFNc3uV/8sJpAkADNh5FrEfv0MSW+5AjokkuB083Y
fsPL2z4QyRmPNdnngTptZuNl8SFRuHR2oKMD+IkGNT7j4tAdD9Hf9EcMNNUg2CSC
F4kHqoR8aXp2VN2A4+1M23xXo6scMd7JnZ3wafaBc/FxsrfcectUcfd54MvAzKKk
L79DubY017sKGpUNLO+/1Hs4FK55CEOMSfTJ6WJjNldDTabaDf0KYmwjpBtbILro
6CBASkF/LZjHSYGfNjYR3j3fNrY5hb+RALBtFTVtbGm2pHxG3gcBYVEwoPfxrcII
RKAA762cfaH0f6pTCsKoJES8cDsf9/T+cdYqgLZhtXjKVZN0/Lk0NeN7pNWEUQ6t
+4uwnE34HTD5d8NCfLcxYx7OcaNnppDu9LYn+DRFd4K8fu7wvrgFMtWC83pdAmIY
YFq/danQRUKcfXO38Bk7Ro7BxDpo1XYcxQNNNIoTRgk6pVtuwSJB7vB6l61f//IO
HaSB5Ar8x4cuTGKMZARXbCBYCa6jFnBeikyxwd8mDdj9zwxm8wKB22Sz0h6PCM06
C+Olvz4dvCigcVyY5g3DGFnA6I2nUST+dFMBqAgEgPAkcavjbXF3RMqz/nGf0Cje
O2oOzIQoBBMtoYoxvc+l8RVr5Q/mF/271yo33qVHNCya6QCMIMQWjhi7xmnUG8PK
meVnc/cg4WB+9D/+s1+hBLeoLFw+5V8BD490lWEgQRIxg+FquYQPpht+8XLn8muU
PRPWUuImlgmlG1Z7c993UM5d2opRkSU88QbPZFZBI/RAJkiJNVMFbVZ0KK6W9QfZ
3x+3VuSph7Ezh6uvYBdc+3CAwRhWJAvbr+WsTO9G9YHSdWi9GgRSJ0qCvZNv+mLg
b4lUpcl/7t+nnfT2d8KQqFI+z7G6jJXrWR1l4oHnqOaOcPcMkEq1MDAO/N+Nz0+U
AN5LWe9ZmQ6XupfBR7NCL9S2l9I2ND4sGuquziOpmWOzEXq1q6K3XdkchmJy/kJi
a61hoRRWCwuT1cWaHY+IELQKV2qi9OMzTEy70/15MEshBP2Y8g7nfm5B5NCkwUUa
5mKh9eTIGTkf8Vfyq9iS7CrQXtrWt7gtKyXNLSy77YuX/NJgcRpbI9K7/2xvcP5h
7XGLEJgN/0hUwCdUvVGUHRaWQBlCEn9ctjVUnnfQSfqJRDaXalwAIB054j+vGZk5
/UsI6B1PvwZk2wheGAzAkD0GA6vDOM0PI1bbk64ZJ9tdHkqIZ0Be6YXhQ5iNrcuA
RP/fTwqyMXAxELlAGwmkk0ljPRggrA9ZXMIbw32Rs4eOJC5GnOYZ5pfacrvDhxX0
k64jS7lQLCAzk9sPSiv7hzNhUU6SSoOwYqM4/ZAajL9w5HXSBgSIVRtp8jukMo8z
GLCDTZsA55UNyNQi3NsSe4NfW2LjWEkUtEUCd2+46js0AodCM9BvyaR7vcCdC5cK
FD5PBs0WRZBxfCGi/D+wFFUS2+sMr49aUqCqAr+9ydBl4vtXZCBYwfxc9xlV0E6X
9oLg1jUM9zz9QecTRhTuBPvCt+nsEI2hz7CyO7gPPB1wcjTTxhk0gALk/BeTwZi2
fjf5+8mlkwX/dxT63JbTI5Sb9waNHvIyBQxpXDMxXxQzJVsWby2wFcsV/Em4RzL8
KaqZD4M3e1dkYapSGztcwULPOF/l2br93fBrUoZObPyz7HPtZy8cQ/iivtCU5MWV
HFaiiKKx6ka4HEsAURVP9qat+f+HPr6NTfTp4hzxiejRXPaGUEElfD6hzhkg1yeH
RF7vsbP71RYiYXyJ3GZ3SPn35LDKRjh9vn11ZRGL/30FZ50gP+wAR4q75I36tZQK
KGzbdXbKQweRq86Uv+H53A+2bLx9qEYr4nCWe2O523smJRtpkaC2+oQUGNEQK1db
D7PB3nEBd2MvO378ffULV6ZH5rlT5WJ2EuPNXjwm2+UPyiFZYKl5UqnE0+820oje
o1uGGe5DkJvIS4ykHBgMCXBtt2+WfVRpW9M4qTlJ3TX7pmEc+4GBGw4diwddWvgb
MQzlfHxxJczH8+oo/tlbL1EFRkoBlOP1gjgGLHb20BaU1ScsDXQsCryWoKg8VJAw
AmFlN54mnFUDPftLRdLcC/8X/2mHOdmFvKwsxWBfDtSJn4VLG6SkDpgTRheHVvYe
rQTN/gO8O2PEYaI2y3urRPOg2rTx7vjfc8xYI7U2aTTrZLJ+gbg3LWUOkhRw3l18
0ZXFi5wlewhhRDI+NdIxtt2K9j/cBAME+R4tjRqgVRDCAeLPtOcDHcq5pfH+oQZM
ku5kUmtqFPNawafnQ7+nuGztzFSIhjU0iCRNGXDZ1ATilXhgcQLtaSnk8tFsNIQx
IcCWloxVqrcVAMeaoKuSoilUeVAsVfkGgB3UgneC6tyHLLLqXM4ejlj3+5BH01NW
i8TttnqWGOkq5veqKQ+iaTjMAC7WBe5vIYGyZsQgiXfFtAwaro6aOsMkeDsB4Ekw
cceCWiBZhKHqMol8gbG3VGMgGgzbndOJEsRzZ1rTZBxQbut0aMvJWGUyYdameLPf
BKSHnumwd+xIQVsi3jUAeufCvLv/p6/uOENHXgCy18jP/Ot79o8PAchxXcq787By
7Q37/iImdmYJI/x6kOHPgbdDXzU5eJwcF5snQTimj+LrSNRnXpgVMzhNo5lReSWt
42Y8Ho7AtFj4BeCWSaZ1PpSeoTraxj7uUxCERaORPzkk/Ype61DEFr9J43Df/Eh8
MKZGXKcX8LzbUjPAWXuUBM2pdqyLto9nKjBA+f6qn6HJ2B15xIKy+Fur9mbirQ+N
tY8yCJTEE450PmeMSCjDNGKgrcekHLhKH661eQRWAYnRSpQz/vhgX/PU3F4OjLC1
PnJ5KWrVWCMu7KmlB51esBIPFfwk0yi123ydmDKbaLTuDhH6x314QZZKmbfpnwwV
A4jAd7THJVvdWH8wYQCAJ/+Gf6RAvd19Kvnjhk/u5l7bB33sG7DJ64/RzZG+OLy/
/7KEjdoK67Mk+D5sfB49pvm+m9/UJ7BuuEX+ufCYR4iUv6GYzh9lllUNCLqZQ+Tp
NL/sRYAS1UU8BUvMTocRWSEbKj9SwG4DwyAOdUKryG+6/r6ynvGJaGoCSTchdDEN
UmSM/w6NsCdi711iVerNspxycuec3gjaMmA2o25XOPizGoj54pAdd674aRYoxD1L
br1MyRV4Oo5T+KKZ5GrcC2H5XxFtwa0ZLmTgm/eYDYN3Ol4yTESecTP6AjQ5NMV/
VCer3ztQnl9wtRBDZF9yErJo8HXf3zvSKjjN7UZ+U8rpKC86B4y7/9PpOUVe8ha9
bMhuB7Fl5lCac/dI+z491vdoDkvS7rZ6H6ed7MfcOC9D8EN+bdGl/Kp5iCXC4RYJ
JhqnkjIVzoFDCtvjwh7R+uEbuvg8sxyDTw522HK9lkvJgUoMsAI6JEoTuLV2qCav
QfrLQYmzQN6uCkjulWyyHHYNdsjxJC3UPpjI/WWx+BguHOFMNX8mQFAmnhUtwCE4
rCR4HZNNvhd84CcWuaoTvOxAoZR3QxjznkQ6xdBd8K1/pu1VA1Z7h7YWQzoe8QdK
Qsoxd8YnYAdikict4MRywClZZwyXETm74iXNgRm2Bdm4bSHPGkfrEK5KYNSl9XDr
ldbynjCf5qJb2GV397qRiIOdIhIZbPhekRZb3+M5Hcjl4nMvKFCsCx2xbSsHQsn4
erUWJGcY43SE688bV3bxt4dLumyJw3uYsEg1pqOb7tz5sefJHfc54pfiu0/wtZLa
CTBrt1PVTX+hYkCAfpusr5cPNOtLW5ty8LsaML94wtR9RAgpxeI5dDTfQO4jVhqu
+lrNg87SShzxINW3Sq7GT+zEwUsvSTTMwrPISkGIVzf41N7Pc6xlz+vA4jcTep+b
HdPxTFcbdtz9UbzeSg4I1Sp/STIUEm2qhq2gV/GSyxuK9Lj4VDTa1bP3/ySx3IWp
OxHK3pdQHnLgYwu+wz31z6kwfjjt7nfkTbT+a+XcnVh+K+gOCdQoQKJk6OMHKPHt
qKhqUzSZ7UO/zcjmKvmk9+EPQvP6Vp0++I4C/by9J8NHXzhHlB6vMLDSImc/le63
bW/V04UDNI8PGpceZU6TG1/xdXp4xUk7OmR8ZV1P+Kfg/gvW53kXpLwbrV003v/Q
WeNjBVS+eE6Sae7SncY7hOwxOGeP+H1SN37hnU2RCGRQ4GxJv/VpiLJxwj3o/p2N
UU/eRn2Zt24cJcpmgokdrHLa5tev8kEoSE74eSwzlxlAx2BdK0e24zaG0ApqfaKB
+x02guSGjOZXkvAvuv43UiO7H0dY0xOl/scy52Eist3qLGV/LavnbPdMUH39Pd8R
qMLOXoOJk92QgxyYvmnjmc21yPrG8t51UkdAT01coK/f9+bDD1qdXsQWddvxCVzU
NjOBFCJhUaqhB6+W0ryKVaktjWdMb+1s8OUIdg+g2MGkhDdpKD5nFVWnBDJSJPrz
gon6mjDNZZXM/6IwM5YgDKMB2VfEgp8KPUx9d+PMlXUkjaWLzRx+Da7rmbJTuADJ
LwTdyDYdgRUwEVv0uBd3lJ3M2XDEMbn3DoXyaOm6v9oAZbaZIIBbISevV8+09a73
FUGxM/zvz0mpN0s3g/MZcBWRyTn0k06FMVJKJkBe+lrmIeTi9l7ww2O/VwaJ6ezN
h0C10Jv+rUGaFQA9S84WLF2aytXu+pxBDZueigKHaN3PlTk49eoU6XpKABOZ/SLZ
9aoNmOr8F3o4QuLzZSjhfCqwxFdVvmCtgrf0eYcwifuQFqoppTJ7vTq4OK5Uy1rh
ctiokYeJ7kD0ugtQ0XiKO+9e1DwQZvJ1UYtBlD+qc9i4+MOefm2tM4YIdK2llQoE
9m7lEU1paqHeTe4wi8qTsVKN4DVIg4fbvmpBrTaFFvig9aZHsfnSeLPFfPHWpC/q
Cu80Dte4+TU6ouO/9ECFdsbyN3tcc2jChbDTwg4XVuR8ljaqyOJ0W2qVQN6vdwRB
0eTaasBJDa7ynwf6M0ZjBNXQ92T7uSpLwHt3rAQrHsa7JKcxQiEKCE5SU5Oc13gz
PoRDyo7ZcllZvrXR1gHj5wOQ7Rc9X/bgSC2FoX2KA3iMRnGP+hKgZYpkG1GIww8z
y+7SDBnivpCzBhUDSTy5FWG6ljyALWMJ4OseIrYW/7YDjUMSGotuv3+H4M/adUVM
WkHuKrGAgggCpE/qczHvIhTViM1IDDeMXYpKbSsCsEO957WyCbYmyxX5u40s6Zsz
PycJrV+UKD7TsOQd8B5yq0u+NSI3uS1bPuiAJU8a39WQNtMkIAnf4U5k9e1xOlRr
9496590wNZsHs/Ty66nLJKsjZ6FdsqGNRpaIluCSwUE9NAXKGJXgIJ1K6y8a5KUt
nBnn8onHvd0kA+HvwDO8EXpMKet6a6WQRK7YiOCG5PcU9GdPYvtSN6T3nRdujyhZ
UfAxGMVb2r4gwyjmgmmuGFeSiWTpdhIgLPI9jBHLkT5XeplsbVQl5ijmQBvmB+sL
j9R7MQUT7+h7C77KWhvATrras5P8qy75ySRPtpKq+EXRyB6zqy3ssZ7lsRGKIE+T
hmdS5EYy7v/gk+CkYPNCwHiGdF+Tg/wjbrj8DA3zSYuCWHvWh1BveaMvt/A6AtKM
tjqKHfUiKpRBonOLhj+CXqe6y6uAsE0SlWp6+ttZcmCGHBX2NooSIns+V5rTNM33
PK5n0307b3/8cwF8ek3NLs4VWhBRveQMLZZTvNIKv035huPvwSckSHrLdZI65ORx
Alq8aOJXWDOt5SOZjltUr3ZMg5cEldSZaQPTzI6Eplr1KFlSfXy2TTQQqVhTpF9k
OJ315oyrfvX6olESM96/1Xw/hlBgN0igPWzyFrN0ergWHCouIAUpQpSTxjeED9oN
qgrn4WxoprfbPce2Nb77f7We6pC9ZX+ufeg0zr6S2b5WOq7ijWe/m2YFCxZvIdiW
VMA0xvDCmBSHC7ZqprVzt3YXoaoldjmoequkgIVAsf198xvgHd8VnQwk9RANNPfD
BRIX6ZIDJLStIQ2SOcts9giykj2Ls4CMPQQX97td6BuRVuEA6pjtNOkyKIvSxd7P
vc7Y+QgyMNP2n9wwKgXQhw3A2XHLU2luWSCoof3Qnu5vAI8yf8AQeFNPAWBsfpkv
aK3Kyr/g6lc+LLSlNoO1Pf0WVBAUmuVjqnoYrDq1Cw/22Q3mmBFHz5jXxENK9Zdh
B8fl27mBCM0KNIQRVqSNxU3B6b17fLk1ienCUaNIiZNHvJBpmi8PV/yb+uYO3S7B
m+tiiHiVOcQq+4zSgI/GkLVieDL0l1ighPcjJT2cb/VnmARKtgbQdGQuhlktVa+W
VmrxkftYojQx8RzzafO0So8XEXF8uWg3rbHbPTbOadfHUuf/YaF/6Mljtw7I3P0n
V3YAXS9oO2UTn1ChyrljkvbTaYCHczmUPdXr43oh0WOx+QnXDlfE5CdwPS7iML5R
MjpO8qIIrEW3yhAj5LuDbnu6sRf9k+qNg+g/cQFHqToFYkBZyXWY8Emwh2IxswIB
3vHlWbKhTEPq0slmZro14RgP3nYfcT3AJaYZ04eFhdj7XmFbnHibLCYb6pDdszPl
yG66FcC7Ur0PesCvjb83IgSWeC1DUz8ucGmPvDy9fgUljIz0IVsrW3cz8pVgpxnv
HcsWJ0c4bX1WaHYyaTLqqcc0Ek3jwmUjNKAmUwBwfPqb41ZWqjea2YogYLMpBJhZ
xCHyRXcy6ocDyskFBcqHHmHQw8GEgleV9OgAo3BBMtIz7KB9unYAC+r9NIphWnfJ
J8GBc6W/gngS5u3rT8IQaFK52D+zwW1iqxuCysJasDGRR8zDXq4GPIigyKSt8KsQ
EQvSr3fXhLZWYcDhqrVw+zkNSUyILPd034HSn52vs86kKxpPEjRMoR3avwrUtvwR
MoJ54V55OMj0RsUtsiNg+biytQ+if+IeYTSjBOtablkfxgciy/l1GJI+IosB30T9
y2N4WLsJ7KnZ31CxNYCgvrqof0EjAsKCA1QYjqbo+DJ0ruTGUq3QLFGTHhNpbp6H
CztYHhhhhk5+73tjbQsin6LH4iRVFf1vy9g8dwJgxXlRQzXOET3uyqgqItSwWqTL
F966kmnfa94PaOgfEGg74/R23KL90dUuR8T5A6x2U0gyzxmlbBAKCveVd0cl2ZQS
9Vzw1Wb/0v9l5tHvcYYH6T6Lrq8HlTAJhzXwPKZEOzWVXVbLtXH9ucSIjouoRygj
x4G1oqwUZgz0toiUYW3AabVaOMMeyH0UYCr70FMMCReGm4epwaj9Polv6yzb/T8L
4aaEkTbwbC0zcVGplZApOXeuMFl7A5GkItnXtVZzvvr514GpD/+02uRZn2XhPCIn
I6H984tr5sgcXafW4qBXA/RrhWhiia3B9tNizNAsBFggX2Dij5cuE6BNlshMpoo8
LgltvU0H9lyi2NJ6tm6NBGpd/GnC9nIin0x1s2aUo8HEHjAWfHrOz1uKEWyDfj02
i4OLXsAUtd+28HlBpxlxrWY+WnAt5ga0q4FJHvEoNVkszBDuy3+mZ0MAsuKDM8N5
M0feUfaEbfqN9CBRpGJRJXuPZYkmNhjrBkCgQKTiWu7/5P8Wo+u4YoDKen1XAUG9
JXlJY4XH22G+5CBGKEtt4pwfy6QHUg5VQ1z9rd/9ZbE0L3mW5dDebXz4qPXYt0rp
sgbcmpNsE8mGY7NBBqBXsatS3DKi1+qcXpA2lnS+9QesrYJuDexcXqSDS93Y9UvB
zEQD1znSj4OxS+kmXJAmRZgZ4SDKgvYAbzGH0m+lncLeYXhxSbLQHf3OJpvg+Yss
gSmarqDXxFuWG0Cb9utkGLNHWMJ6Pj9aAEGpR4PbATLcBNMhtNeDCJDUjeE3lcnM
LbYMFCt9L3ZSrJogfz6ZhMShBFjD8QpJ6bJHpRbPucqFgQJ4AwmsnOYee1ra39iE
WEj3TwDyOEqYThBy/6Z2j0D6bOsS5s7yEIn+VZMc/8Vzv8ll/cT/lKKjHXQCMwpG
iXWVCSjG2SSBvr2OVqZk5YbaMSFUcW/zEBvC3dSAQig71ujcCAeBq2YB4X/NBrPK
tsEGOM2ynIEwywehLz2KdzbeHjjU6cLCtku4gbd3Mf0IzeVvDx6rNdQOFxHe2fqM
TBoFnPRELmerLfDcKO4IBk5l/V55VbpJTVgvhfWRfyPj3xNzCIYpcB7djQ5E4t+r
QGKXLfSGtaW3o27XIXeQKmeycOu9FVKuHs6Fm4+S8DeTbsJDW1mbecN+5syKeKJn
UvDg+/2FL0yZKHxGg1uAjCbItkwM6xlezsJ8BLcKpvgjnQ5DuwDfV5UsTBPAP0SH
ph0gnWFw0XgY/n8I0jCjB0FkCaUnhyqO4mUmWNbtqsVZGtNlrhBqcxuUWJndeabR
ebG2i0vHcTkzsC/0bwX/prJFzc2HYaqNaAjHE8o8NOV7ipQdyfH9/QAKNqguVWWS
sdiM1V3vsWKzkIqaL116AKivbNmv0LsffAG8xEPsOBEAmANdinYdkGJEMyY9swCO
fZTSMNhDHTlcUA6g5ctKnEzWlR3pmT3LBDPnL0Ud0jiBzVABoKu5nUTXOzO9+rwu
qd0no1nToz56el3CE0MWJ9A995rOyjQac+A3eIKWyDy89+mB7idtrc+W7ti092jz
BgQ9oO7uNz9LhEzF7OX0voS2hZowa3zL2eWR9OL50YuoqlAYE8n1+1P5zDbAnBKo
NMHu9MmYDSxsuxGCwAMTKePYuXI/CmGTT0EMX9v8XdG7ljL+rq9ZuYWV+YW7+S2C
r3uG6u2SGa7YQzKthovSljP7zwOijCAqasr37UMZbwgy013lac/L6tBmSe35Rp1e
VMdfGyVL6vM+fQ5GgZ7ionS/GvdDdFQycZgaBr/pDihAXkRnewySrrARQtgl2rsW
GpRbMUAdEtxW2vF3mYTJgaJUhlP4YavEsp5P3MB2TpYyFBNF9/IXjpDuzEZDBYuh
Vi5jawZhBySKgS7PtZJpyFyXq+SrAJ8gv0BGm2BlHgNQGge1zp2QwFQwQKreuUrJ
He2CbdIqKEZJUiV69w4BtnRY4dIFvQ9Ahnma4Zv1bzAxLv4PY5mhUtURDg1MnPgK
R8nA412PiLr2dLrwMpz5hgqUG55HIdWOIqKQQXK15ceHJiMsLkwq/Jn1ccAYe0Z1
oYvUYIpsp6Y/OnKwZFOl5MSyZle1YOCElxaBJnFxSL10q4XDMh2irl/xg9c3H/N+
teTuiHpzvAt7TbdhDk06SssWcpuoNNBf7MyfOgpSNAZM0j9Mlxaj7pW7LNKLDQA2
eVjz+WzhuEsALJNDNVwwjdNuuwuUAAF2SYHItdHNUWu4SMphYRvbjFZIzWsbV/f5
5If7etfbHEwPprrvImLmN514ARjCLNtbSI8xRTt1Ft9qSnFSlQiDWJbGqNLqHnF7
wl7voGwJ8w0N+w/5Rf/TYRiPeuku9UtnUdrOSYHIsbqz8fmUMtjfM28M/IhvdJmS
IbLxheV4jq2cq2TihL0e37ciNmoChqXRpjFytfs9IoK9Js77/a5XyXKvWnZItEu6
nsrf0TLiRsyYVOO8PRVWHBlFYx3qH78fF9mDYlPewrXzty5bnf6R3EYQEkE+Bx4J
wgSWLf4sAMDU4+gu81PT9zNBrH/CJTQimsH+W0EjDlV4idsa72yCCq4+4Q7q3/EA
JgAIOVtsBuG21ZAzPJxgHXpVJ+tDshltWomOivnqrdVLwOmY1UhegRvSJoLVzVTn
CBGudZ4/YmfklxVZfMD2GSXrZkLTsolBSUiPV6T/1i+t+n7hhjYg03PXotwMyQl/
oeTWU4Du15oI0I0fKYXPxGd6YlLzaSihe4pt0lBJj8rKxV8bvVOsFhv28pB60EEb
mDAkLbuy3tl6hcHPvVw2IQ+IS8YYkCv+EoWgavKJ//pyXqyVNq982NqLOnn72dw7
zsZGSePbyZVOMK6k/Cky9ASvql/TCFDGpn9dWcc10qVB322haBdn1SOoRAolQwli
KDav6PTikYYtlJC27Wb9LNCnFaEhQeQ7MIn9gRZzfKmRIiD91B7zZvz/A+uYAIwQ
IUs9nz6XYXuVZ2aUJ6jrPYLy0DAl6hLO+KJrvjhzbeBKt6O2u4yl/xYiD7FTqa+q
PYZI7OzPmTUp3MKixUCOs6G/xCqzT2EPRKFHW6QO7o8NqiLFjbrIsYubif+nLhbm
ihzPgqsp+re55HH33kl+j8O354ZtzZky41tEz3VQjXt/Z/sA7qYYFBCuq2UrFhHF
5eBEWcTUolumFz1x9XLHqafPSeSI5CVTNoLWzdyDNMCkyH+o2y5h94laPfR0lhQ7
ozf53OGoKEEDGrD1crmUU/+tvbKnHq7oL6lJm+eoLir2f9axxMM3lF4SuknI6LVz
ja3L6YvevPEsBYeeOwmOq+XUaRN1r7aif0xFyUftIwBYtinYpViG9ARbBRpkp8De
HVGAcBI/CezS8yA2D04RRP//Tr71384v8jimXyTTEGnwiBQ8k1LFxUm7ugUE1kwv
PfmqlXDrRJQsQYm8RxLnuqkA3LxVI8waVuPyyx9gn1/2G5rI1KZc/BTs0pXG2BWw
SekRjVn7WovoQqpPLhvAek6OaIeYiYvJW+6k53SHzYmyfWrTZzIXtA/6s8eEOiBr
gQjmpfvb4mCEldZKo+HsHb4o2aBWdjvONpi67lsBGLZTrenN2tk2suymJbFEqtQS
R5ogQUtQquplNyXuTsG1G549AsLMYq6GRHB+8KMWVbpKRGLcwxXzoZJfxK34q3i8
zuDR2SeEQYbhbb0TSFLj6pE1rk5kJnAFXSMYd/1a+ZYj5gXs62ijz/+8mAo2gP+Y
xlrBKezGREAVQ/BIFR9QMxgER/B67DPhixJF0RCclQ2Ym8vCadQQJVQlPaY6OB15
RcjxFkZ1Nbq5DAeUvgPxYjqIeP1RI/oL88zwea+RSHgaOT2ba3zdIHilSzexQX69
SeXa62ZTDRdwcgWK3plLxXL62rS01wUniCesQquGsx3MGaEOWKE5dHz7sSkZQyIP
2c3j/7U15YiZL/gztLxsElP3wS9cCFVOtcuzmW4nbynt80tFG/9L8HLdE3iDPaFt
nk6RCZtZSH5NL6Y6YDHulgBUOYaEuVlBC65MHfWRp9V5POKBpZG7ISEaTKkYf7Mb
EkCZKJJW8KoaQTzTP6reiuGQi4MiUXVpE+wHAAIqhZrPZa0jlE/wFePqILsFToWG
jcyZ/xz8Zs4mTiejZIWUf2k9wr8voZPnd3dKsx5nhv3zU66rGXURsmgVks/ply1l
vmjAW4b3GTjgZ0/WdStfpSf567cjfL86C0n220kyWmcK/Cozi76l832GOsYssP/B
HXRNUxCezF5S8Nbwr3oeTJ+HVhqd5koQwEKtn4wo7e32hLMCTUXNCGkv5eHk86zp
n63NpJd48OJir5NIYbLwAmuiSKyKpwq/h/St2/MVHpcU7MFNeyrNETR+IPa1MrWs
vjDQIimyIyyYjlPUHmwVvu3SqJ2gPt5KWboLiaL5d0+dF6FHyjenNPbqm6TcOV/k
8p54/nSjONoHcjGxVinm7dQUyZ+Z2dDahL1gs/nP+o5rwYm28R9BcsI1aWjq0qK8
6j+5CFzv9mQkfXvbfu6zbkIZ7B9MqqD+8FRgSpOlLqVeSyFnWpCJkouAAkR8jPdL
sbzrXqcxsh/hUafiH4a2itpG7xPpFji/3BOFphB7PyXNiUvvs+UPvLjYWKdnbd9Z
qtT55NnTTy2H/7rUP0dNUBatesQ4L0BGofl6GTaRZu46L3th6CfMwHoeNLwVKml3
fHJL06d1F/fYf5b29BLfon7PQyCGAISy4ock9Znj7hn43X4ssl4uIZWEfSTWIVQ/
ZJmBKizPlblhllsnS4y0ia4S8uoj3gswIADOKNEmFrP6G3YJgTUmVnZVQNGRTRvs
G6RtahsSO4bneLpi9SnxihhBY+MDR7KsqAzG8X35wkPnapYWQympgfdAt2Gdb+gx
MMEs569YkSbDjNI3fSAHvfUg2HFiV3o0wmMdXEqQAqpKdoLYsOmBFe6tMjy3xs4H
2eH8AWNJTdu987bpO1yylA1Zle6KaULPfplW21T1L1qBfyNvU3+bXZBMU+BL0GuY
bK7gQ5ReRqRT0oa/x5hG5BoV+OektYQSscRzT2HIvIrHevPeBi1KzGUWQGQedDY4
ZU3wZhPX8czcJrWiHqB9IQmE/TTtZbKl5cxM6klgE9T7smloYZc6sGKniwYE+KaQ
IheKarClz0/ApsahugY4KW7s4gu22lKgngI3r5ExSV5xlLJPVapOOi68+fl9VT2H
d/zHXh9xJksXASWcDeq+WE3vab3vqxQJMqfTGSoIySaruzfeq8frjnpnLday1VbI
hMdm0eNJsWFFGvtq7FP09nWPrw9uts2lXCQPZh+PTEIXa9INNaDw1hFDreTy7J7v
OoYloZSIzeRElP55+C5gz+gSitERsdRLuQKMaNf1TP7mfqAvDzJf3XRyp/Pzp/xO
eMNJN1G1iM+XnNr3401qE5NB/p4PIqdV8WeLqVDMvjb/t87D4tCSm4goe6yHhrql
Xm8kF/WEuq6qivvCTPKyKe2O550Eoi36Phys9ttd5wpiUdQzPcIHP91mIhznyBET
7hUy5pG7U1nswxPFXJoGnxZ4JCiilNfNu64pPIhUJ8oJroyFAlornlT/9DT93k2o
UawSh8w+ejnvEAgcW7uLxQNsO5ZKrIytnWVoFZxMYpaegPkAtNqa3LyqYytdL8pq
65ZkRfEDTJqCmROHI2o7IOKIg56l3cq5BmkTo1ZSRe3S2kHUTYY+9btU+v46Qn9c
VxWiiOyaQhOvDENod/fAl0m1ou530GpMSO47Vlvuycawt1G1aZ2mAcuLmjsPedtb
kKOQDGCDGIrUxz3GIfLKFeq6j3574ZZCTC3AcpQfAtu8U/+vwnzy41bkxUoNAoem
uN8qznoSx+Bonza4dV2XAHjC5BDlhNRXftLzCs6m9qcfcuUCM577sGy1TJL9ku5M
ZtI2zIi4E+Tad4K0/Ub0Ew1iKsACPzEfAoZwaR2EOYRERLnRkQJDeguXEBcNtEeP
+WvUWTVYwaGrxGysaVZ4YJBVSs/vcjmKSeMbBkeNbfsPXQjdrSLut7QfunOalkIO
xKlmXRrWqWNwlQgTqqQQOX5uvTZsZ1aYEqt9cFAlSz+yrjP8sC9X1kvNso7BMdpx
5KXB6ln1nIkxkYN4XI5RjkFsCEF8Y4cLJzzThVcP2rB2ozqLn+bAbgDvxO0X8GnR
1BjjScKJZQSvukOD/7GywDK+ofk8GXj9cvaqQuZJIIZBPSkCI+AOHEgMQj7UURDA
V1oRHB4SSKou8/pxJrLV2tk/UTo7rPcChNYtS1ff7fZrqoQilBhSKj/PTXPyCnw4
qAZVOv/HqQd4d9JhctzRdUYo4ZekEDGIdfosXB/V/2gQC0CIjjJQlQ2PaBClmh5q
PxkCsigSadXhpWn0wNnT0v91Dzv5UMBBiojANvclR6alCXNaptKugET3AWWyBwMa
riy0dqkfs1LdU3s3940C/LNpQMBeU3QYpl/cIZw3skxqI0T+YJH/jm9+r1bG5gyB
WX53+oAn/uCLjFbuBfofowIkLfBxw5nS/rN1In8b7VLIW1Fp9LRCK8bfHWRIhjrD
f5HNYv/y9UjZ+USFO44fd/Wj+gYGpOq+ylWhbx2qHG/IRb7kVZoODfpnrrx7XTMJ
dJXrN9wb+wUJD70gizEQqdVe49wMb32mwfxi5l/qC6Fj4tYTNGk178YiJeN9RXcH
v7ZU+xfkd4CLc4Abfgt+qPsuw0GjiUbgTPiqUrCP3m/KxeEa5XRbN2PJy1JxKDpd
ihnXgRrGrDyTGMJMr7uiQiMhRYSLRZAj0oaTzqlag5NROI4z7nb4ziFyfspTNyMu
DEyzCp6zL6kh/Ut1BpIroFo8NvCLkQZN2BAQfXjjtoJ2BV5Gv3nUCZHZtWcRgqM/
b2Z/ts4QlsXUlmDicbmPK/+DJOOLkVWjYiTRGckpqEbj7F2IXJ9TQ0a90Ezg7BvP
WHAYYBIrX8eoY1FzFvwKRqE1duNtGkJ281lo8TJ/xtsA45xLFt9eAqxZ3jF/5WER
S2dnBAhcvHvGUzJp4VYmKzvNgMkC0kfDcGlwyqqrD2UQp9buPKbSwwMJd2tpeReU
KTHX6Csh+I3XxJatKLyQpObyE0rEbDI80GKI5m5bQAkdXlVUZgbD7QSCXIurZUqd
iv1BXnfcRyP8ptgsULJXOyGC0OJPvYO3rs8phQcQTCjRqzBJ7cN9Mtqf3t199yYH
tuzLjwHvFJfZLFtGqBQGOiPVXzDSnEhD45X1BPujkvicwFMjcMCzjpJvq0+5inqr
iQYgbJDFc117dIwUu8kY98IzNisrpgNuM6joYo/zEGOcqJvmvamjOnw5DlgTG26y
YeVpDPzbv5g3ejkgod0/M+cHjGABCzescmQqA1t09Y2DGz+j1pW5nN1tvokwpl0e
REqDB+MbTXhXFpo8CIe6xODqp9K//d16zLfLiuMiJ4Q07M4izbA5C11HQL8eDFt0
jnp3HkeOH9GK4sGJ4gfjaSgWr6YjuRBDnwhcgjZqJVInY5uibMymiEAp6BNGJ1AL
60hladYkinx8hgVcqz64PDdB9TTNiswRBhg9q8jXeCGsirgTFqwfRFglLR8k5eW2
VCSoagj9nd/wKuWpPK8sywaDH5RUumOQNzrGbtCZJFU7td5L/rB1k01glP3ag4cf
kmzAq+g3lKkgnYDNoPuyCV1T9fBBfjI9LSShFDyVY1dAE9qxduosw9WU6POJzqH/
kpjl7pty8CduUvi5gwIi+U+3qf0zNeZMUQ/T6oYnskbvXlISabf548kQhoCmYjIb
dqPeocH39aFL+vLobpc/wc/VTFoFrU0thE2RltycY/S8FbwOfec2C6u+oVIjNbW8
DmlCj5HjYN83zYel6bixegwoLhR4Vz4lq05emRUfu9Mj9rUzcZTvkxpBE8L8zBS1
L44DLZxIfQQ4yVonI60zxSZyuLzCprlbHFA5CJgzIUtexsB2ebnX0CCJgicnjI97
qFyJvpAqNagjMngVvHY/aZCP7xosm1P5GIzgqj/6rug6/VWMJQGiTjSLgZdY1Ixg
Zk8y6PySQX116q+gN+vO9yxaoCHpZ1IA8DZ93R4mpbqodCoUsyaf+ZeC4y3JX42T
GaZylcObcfxh6Sau67ofOeC4uw0PZEG+aNL0jHqn4u6WAcge9nFw9StPJoYFbALd
HUX1Q7KfLmr13UP8sz8ypaM+oNcT4pTL0Ebmm4Sl0u2Mt5IZNAU2mklEzqLKETp5
E1eSnn7MePcj2xQzpYkeZaZMszEJzS1dQpkvGP4yEhIgx2fXJW8EmEBJlQO17jSs
ZCsRBmh85GKHlSMXH3ixsgHP0UotjD1q7hXVwY95axv4alSjx8CndaEQOdYMToJT
bc45JIq9fVWlqjT+fL3olZiiNY3i8FVQKwnPkgDYiTE6WrQDW3wdFlQuo3AbrvMK
iR8cHDsKmOr0QKtpRY8QzCIeehTUc6f7CCgjlq6kpayounOVAD55wBIc5Pehwska
lEhYg+BX26V/S9FxO/HEHoUpWCBtr83ImfvyHQbnMkj20oQ4/rGkbFLKzrbPsMqI
Szs0WCN+H0I8/enOhlj7+p9vAkwwPV7L6syWZ154BOfPR6BcNElT6YLOigKYJDju
Byxzdy3WQguZpWoJmy76/1HpIynjBxMM6RffH19cETxiz+/JUisANnVvbmNdGu4o
SlDXgrSgdTvPdZccO/hLLeCTRw3r2MA+3u9uH5T8o3I8IOh3nV/hwd+2sQYOd9pa
RdmykwOsF+tx/VEryy/0ooyKnfYE94j0HKQzfy28dhAIa7DM+OVP99lpNdWs/84t
2zmbUbcLM3F1SIs79U/J728+IXBuB/yz3AK7YMimKOys+YwsTT23pikjSNVRm7ZW
pGaTyyfR7Wo9AZeOU8TRbloda9icnNJ5tGHa4yZGzXFjSujliYta56NjJulXEyUB
TKbv/NS0VNAvZwxFnhJw9RzekjwpVBOQbyDLrTwZARgBTBXIDFyRx6V4utbnPzYx
O5BZQWjSh3zFYIPYTDZRR1OKuP64t7+48c66SgDoDRna5/VXKWaXMUucsp3nq0u3
wnDsh9vprlPPTIuS/vt1+aC1aG2jH9FY9iwszQAPkhr034xMjUmGDxi4iTWygz1b
ZqtwoprS3ZmDVOWWkBQD+xlj1DpLOgrjPVVVLdluqxXI1SYh0DhsNyepdWofQyF0
tycVHIGPyyMC/EpqXIRC/8vSl2FoNdQjOhJCxiwSinU53SXTGCzHkfbgfAADT1rY
067i3PiYerjrFVDhV9Oy74cqfUG3/4GPnzfAHeUVjdqJFn7ubKuoLmqVDbxR1v9/
WtlZb2jwNnY3kM9tvN/H3FCaEs1C/+ZN685WjLmqJvqeD6gjfD1KLLfHXikSwbgS
zlQUwCiFWh9YiNUyadwqQe75zvETwnnwyaUJQ6FdgOakiLmm2SQmFr+DuBXd9w+s
IXLegJDI0sqcxzLMikT6JX8DmdCt7N1GxN2UnFiR0xiXSLDIz7ilARKM2PHc0eHy
AlgHSHl9Wu9j9tgqhJdw/dldedJsumma8yiwihaKl+XvXc8SBD1ei2qjJ5NMTzcn
DbjRdOxFuDLmD3SX1wM5kd76rN7FwCzMzxhrQqypI61Ga18ESFsOG0Kr+ghWraB7
fPXDj87DEHsnJoVVOBPo42K8/0ChtL96WVwe+52fRrFFp9trt1mIQ7er9JyZALS5
q3QJIie86/GyIp1e1FVnhL7jitiRDTQ0w1c9AL5zrRpWwLqoXa3zxefk+Jdy+Du0
+jLu/x1gUSclQ2Fsk5qDA7XKSlTllxF+N2t3zLotYc123aCPTgnRAr4nRjm28BeJ
P5+MyTSGe8SGmJBmybtDQfYCm5K3vNJE4QVmN9bWCflJu0UGEelMnnD496VAaFJK
JBFiyHdKVwx1sqgTcIjD8EcSbelDrhKGHvssihg+M5zrTyPY2fE51U5Hd8scTrlI
kojZrP+uXsO9w3R8pNjNzG2u4PYTSVfGEhV7WvoC5sz3LVGgJrw/niQQJzXgmTP4
Dr+2zwhjbGUQhnq2eLqIFhNEQtakniYewNOda4/7clNUI41tWYYw3jmm+wUk0ASg
4QMf3s4LU4xAsWoODwhYGQGYdPWmYIcRVhBWKCQz9lAgtjViqBKKZjyCw6zMJ4HC
jyTmF2QhQFKfWIP0VJej8uyfvUm38V5LDZGCHj6eELoce1SEQcO7izyTnEfPb5dq
n3V5XASliHsSAPN7gKd2gHA2/TP4I5eJfVcF3vBVvweIAjDL1lOdHr+JYjxEchLT
GdZa7/aCG2M456Xb7FlONGvZvjw6h1t4Rv9dwVrnolrPA6QtG11tdDgBNVaRIPLW
3Fm2pEoRUKKLUXvj68o783rToikPY3sIoqRxGSEyl+li6PFIc3QTQVy8M9d6AK2X
TNa7TW0/yCuBcV2f67GIAodTrdu2mtk2evN9cMcfQH3wTwZe29CDCk5H0BKPKNnn
ovDI9jCyXGdJo5Z6i7wweAv1Uy9tkJ0ZCfho8YBwCxq1ruf4hTkRI21b5u5fUBHT
Ilv/8fbUfyIQcjkCmb3hHUYEM1p/KGpaXT8am18mIpcHVQ1oQX4OaWiEgVG1s1IV
9SCla7ozbEBbKQ3ff+qKaUfT0Z5uhTY7CKFbm7XsPzirTUBbdAGan9Pgh0ZHaxXQ
3gT58FIlpFsJ3zi/xgAhtyrNvAb0ygIvdCceFKTCX7OqNzD/znwQfkSmZr/+P+rJ
6hlwrVtdxRWqwnf/RR1dxDLaBZCTcHCm6s9v2LHmxSsr8Zj4zR5AG3B8AEVDa4D+
+uZ1bAcnMHnQpBo5dNlLtEfbJIhsyAoLMWfRzbapvvK6Wu15ir4o3yzjLYSA5vCo
Z9p212WmuE9iG+0WRUUMwUUwmcBES3GWFCOp6arqhB1C3XZETWeOK1ULM7ZXdk15
rlOrNZns2BzDEWfKxUC7Oy8avVlTyhhIDJCJYcdREp0Zw/5j+fOSteKr8EEnJBnI
zU42fLwwdDSsGSZ+M5cSlX1iRSLZ8owoPMwphuJ7/XX3W2D3ZEYh96O6eob6DGhJ
9BmTbEfTDF/XUs0sRPywiy5tXoaz1UmTHLTdNUJsinTAupIdzPA41qVR1jCBEAZB
fAzvf3uZyJUEllfU7sY0F0jur49vrksfBa6QhUlIUJ5bC7ETRU1PdCgWBUKxTcAD
RkmRBkeo4WxCYINK0vHUOX7ZU77HioO2zHYhycgULPqxvxFnUTrfx8mPPXcOJ8UA
7Ne6BMILf6Nxaq/u2dMYgt9EJV6EDNzcWyu7DrJvcz5caJjJNIrH0imyC7Fzs6P5
/f6IcfgFYI5t4FAKPNmd//MohBQ7I1qtE7Z9y7BU3NyBSJURJVXm7UKYyxokqOWk
TMzDJJHjSCQZFSAeTdX1lzH5XzA1KTp7T0uW71qMgUwOl+zAM4O4+LlQ1k6aP9C4
KfZeks4oNp84o574r+iwhBSpruIK80XryvSssGKcZsY6UK5Q/4x43hqTL0+/dzzM
YxmwNYdOjyhcyqmuLspUWhq2U+iJS/y8IWqidOsPHngZu86IrxbymORxCmxLcX0H
GtJcUYI2ywASkV8CsmLM7PUk0siA4ZFXzVSDj0qpkrYiSHcdg6VEp8OJYHBz5Tzl
D4Fj4aRslQfwEfCqpcWuV/zoyNX3yQRHsyYsVskApVCz2tMbb46J53uis2odxrB/
Pm0vUQEyP3WcgQIy4ABsLLjnRbsARXYyvdHKfcqondY6ORPHnKxgHymVdoKHSqGR
HhxFYavvFI/BCTFU2+ydEC70o3qve5Wlxlb5QMZJrmspqqpvG0JWCc2goZHlGXCf
Avtx1as5CuxZxJ1/LkPvKzVClroEPnX8C+LpNHfGjfgqxJYrjI/lAR6m1AdFT5mw
/DWzKXvM1lDM56ahjnWR/jx23ugHfi0RvcM1dcCbyq+T4dZ6cIVhYcu0yYbquoJA
bBVcfEylV8k4vRAElqEd7ZlOm0ReK/Sh+rwUEFmpRUN/2JKgLkS4kwlGGRy2hmFE
tAFmB91y3DCozJVmzsEqYeu9lCxdIOkoGmqRohb3+RcSPTSm0Ira8C7zKrNWw9e1
gea3vNUMk3z661Ju1WNJ5o3IVlcrUxuFx57Yzf0tcCDtHINmwrGyio1kMgpt8QIG
KOpagqJhQ/gZ+0TaBUO72TofDkahFeRdhjsVbTGoG6NeMVfJqrjT0PFikTnNNc6R
5xxF9W3XEq30wYgJge8HuhZvN3Wr3HkST/bfLL/8vVBjujfHzB4VTYDjF/scfkfQ
RTRdbWSbq+AY1ygQAv0qxRgtmvpjZ7qQVfk0rS+X7G7iLvKjm5qdCniVHwLonlDg
HZNAy6qwxgVJUGCx0K/jrdWK8SLFnfRSufXsGqk7kkh5metqwCr/Jqx4FmmyD0da
6IbZMWcHGal9oK1sS0zh6kqQH48kw7S7kYto2g4rPgfsVK5m0ojokrdKcNo61Y7x
diaW0cWJAsHq6tQzvOZzPH+rxYqn5aXazTpv4fcaMhALVHBH10saupfCHKEUexsR
hEy16ujJ5xzXpjvxdTT90MwfPdR4bKvWTt4Qm9j8ayOOKAsn/2yN0/RROYi5pRPD
d6HuE+Oz8XNPFwZSNjLaF5fRTDO1iHz1wFFml8wKpJOBK6Kom+kWo2nieIUznH/V
9j8/v1utvdeAWUOunCTvt79kxZjWZoryKl7onhgF6EsKyelCTUCKBjdjZtqC7GJG
oGqNnDnn5kJ6Mgzvk9auhn5fHc4BJYlzkaRY2IxZcag/vZOCj2TvS60iuwmGWJaG
HEGZOBA1wjHTWBseMbqgJN6P67U/wMLMm6LHiTWH+71eJC3Sx90+O5NwpKlpk520
zTEXZ+6O6vzmqHG657U520pqqmKpdQvoWqcbjFL2cUyrdiNFBL8z0BEaIrbbM9xB
4+uFVU4VsxsrsnyQN5Zl3xn+YsRO0VtOPRSzJITftj/Hj2cndkTaULSjCLp4JVIm
wx5JN5ZquUmQRBHPJF6bVhactClbjgsJ/Qh2MwAKjHD05CSEi5fHYa0Q6Re3TCCA
ANP4AeSgxxxEVUJWQ8Ra0i8vhyo2mhts2y4qhEvPClNwUGzH0bBhzb7+5jJwwOC8
oU7VSMEk/pDJJlz8MPU3ruAYZsdgRUOdpGNQFA1a7ufwezHtmXW21re+gJKgWqqs
hT8CtFMn2ES89HbnQWe0e3KpwpHahD/VfFCrrH0keg/C4U2fK0uitbg0hBR6FtJ7
GE5nwIt+bo36KUu84ZjGr2L4jvVC3uWRINrncHk0fVhvNiYStYdGL9ALb59Q+31f
GrXolC+RPqn8orH+avbj3UJNieFJbjvZUKJNbQ6ZsEouow9Sh/KyUWEviqfHgvcb
O91FAGr2d4lXS60J+85LobQm59Z2jXNpai7oXN6Cw/Lk6ciNHwqELtHxE4Pq5A/N
01KhNbmfiERC6qsatBRsrlgjRu+gfewW/ErPtzSVPuHfFAF+K+F7suXdzvjElimz
0asX9Wvlh1HUCdsvra1vj4RO1CTLOrkmrg90w9UGFbC/ZKaMzyl4dOLghyIYNWed
fv3gVuw27cJfvXHPB8Mz5xGD1M+AWrJfSkLggSxarm4DfDhOlxVO9mU6B1VRTQTk
cBvanQ6lpWb70f9+gZU4yV5rEt8cUMcgM83aD24Api/1MtrUtZ8EdtWKraStzx3X
HpMgOpEujxuswl4aR4XIYgvHQlsD6el5Is4FnC+1cwSxjj3piiLrtMpyCTMHOxww
cBDgv+cncTtPwT+fu8dhGafpb1D8kHZ7v/z0O4mAUIhGyBEay2uSXQC/1NFtHFhh
fcjuKVqVQlUs5Vn8D747MhkpBNhVJN19+8VJdbLZm7DksTAMULE5dO0JoxCm0+M8
dQvLsw5AnKk5i8oK2QDO/XEPDyeQoEoVsGKznilBpYS+tgWPbrwK2YIxy7+0KjYE
ZM6Q7496Vf9Un2UsetxnZdIEgxGnbbdAVa5T1MQlXOrZlfOaDovxt6luhhLCrsIF
svwZdSXvY5gUyDnCT7QSvKGwOGmhqshmUD5igQnbj/Kra8TQWwqWZgFStWMIrJQI
ac5sqTtkj2Q/JJ2VhoJh4+LE7irAebwSosuN5uAC3yMISrurpiYAcjqfnaGZvfqp
RbVG2C8KXYgaZhl7YIH2CLcprlJ5yfr7agimieZw0jPw5wWfgy9IMOKBfiU0owgr
JBxAZvQB1G99lFVxVX/ZVBtSERM1fpH6Cg1PclGlgZ1GtllhuBbCIijVYXpgr7Mc
T5CSTZj8F+rfiYJekfdEHNXy8U++Iuv6eebjlef815VBE22sxxpqzV67H0p4OR96
JayV0GTazjGJoPYzRRt7omZ7UJ34qAyi5TwVXnjh+N4uTU67eyIzzGVXC0LM8iL2
lkVM/ievkGXnSBAMvCzhK3sGRvAi3M+XqH5v04B7BB7DpQzUgEJc/WFVmcI9bssN
Y+fjZ2MyAG/RwBHXtaIl/f6osROn2Mv9sQDjN6GJca9tq5R1IMV0St4/I7TSdm19
9zdDlnWE9Ak7tnpUk23SyFUY6k32rPlE49EiJCz1hMAFCNNVMO7Z6kk1Z+9MWZzh
39TqTK9BwohMPHPr+kdQd+p5/ViLFqJX9kMX1WoHc7h/RMphuydLZJ4mOxbvXeBe
AHCozPYf9kf9a8D6qFSgDwz3ryjByhpy4q/QWh+5pM36N9rL2ja4jIpw7EvslyCE
tfx6cYVizOwpgLrDuDGThmQAgO5x0E8zS001SosazXjNvl4dExK1Cq+dFEy2bp2x
zM5J6aTxa/+6WgnLFChNRJAZZ8EoDd45Tta38pd6Yph2qEzd9hpPLpP11N6nb9uN
QWRe32DOAW1Kvv5pKjYo0FTu4QqrEyYB1qiEVmb70chTmSoF27FRcGMCaJlsdh+V
ohYrQ5frCWfR/GHrh+S4Wcd62Li67i03GR9yg4hE9rZTZ4UctGBRAwxiIi3P1Fk0
EobrsKDKznbeppefjKvCbk0JJSJoHjQ+N94cMsTKSgi9UNIk64/vffeCCP+B+8PG
pK22PZ0eSkWOYZ+mQXhTlNSKamFRs3RAjIC3p6UpKXSctLN2P2WHxlTwYo3/sH0/
TUNTATRLB2VKCQcRA6h6T8BM5JMxZ6Ta5P9xcIqdL7PnoyYlO4yzfa00OSnpEunQ
NohuA96LGYApGlC3ffuxK/5d6hQ2a9QrXw/i1t2xB63ujnksWVuDK3NoErY31HxK
N0gvVK/t9SLSbtRJGrRf+QS4dTFuLeQ0HMATMVPNG9bacYqjjCBppDjyk67DLuS7
VmR0APpHWD2bhEEhnUXwTkbG0c8zs5Ns58iDNbfq9+5cH3kx7ia2yRw+8Y2KcdVh
jIr4PPsQew1EnDGdwGjB8nwaIUZ6y7WYQqJMq7gTgWjxhCYKa+GL7dZbeWPKnV8/
cScNVI74faUdk/504Th63X0tZN+In23f2TMPxzOPTqwm1czpdLECaE6h51YuB+5G
7lwgPQtsGgVt+O0/OVZmFcqgp8yhltHaT7C9cCNpDI7Yk9LodJEdp4Zs4LL3700O
HUUwEBvI4CLVcNPDkv12eeJfHYJlllKG5phR9qqnhwOl6b8kK4vMkYEaOBJU5hQ8
LbymuACPoqkW1xv9L903HMNfkTxLGZDnquIgAtCaay2xguPHNdWaXp+NwrZj3tWn
FI954IL8PM6ssQtRyNOVnJMy1iXKBUyv+pqw6qNzG/HQnixcJDJM4w1r2d/O+SjZ
ip/qvg8rwavcr8RLF02Oa/0MvBfO8n5TBk+jjW+9mFX1/QPwBHcdKprglH2BE0nZ
SsnzLWcBzxJSCeSwvxZTbHx9Brj2n1Ty278zvZIJAEhLFLGbDSAN7T9r8lq6gEZx
WgeArg2BNunWiaJXKz+EEzEoFyd+ORbC1TY1g4PbrojBCZM1jeoTrPnCcMYHiUXb
3UL5ESwiPl4Sc+cdarHMXH3MI6zJHOLTq/soEkJv6pG8vPozMW41rReHb4z67p0J
ZD7IN3aAoWPuBPD7ZsISwe81PWZu0TUoCTm4wxLI48kLkEF6V6F1o1SsMXtZz136
uBJDvxAh7ls8d1mMnbPiRypMY4G5u+WEi9O60eMiUU1JLOcPwYBsjpbqlYsORfB5
osJkgp+FxBr2XWnpfhXG2NAtq6ii3ag2Ipofueh6gMgrs4G+RPWkfmydhtQlwTUM
W5bDSZpDA+i5z7kIy/jXWzQCsEGnSfovPth1K4HiKkDi8Ukwe+Kw/23WAXh/FSW4
05g3GefTPPWw5AHdcx+WF3+jyYAqr2LBh7uImaXsv43FUYbcjwmlJkg3LMDItY7p
+Syfu2jiH6SgsCTdiNSe+SaEwMa1udfdTlxUDDhUiBdH+aftV9qEbAKowWcPBgXh
PR0B3qz114Pp/1k1y+uEvdvi8OvjRiW7v8fL71i99pAaxJ7jhprXr3yAiWsgetoT
qFpETDq0SAYypxCc5FJire6m8QDlXRVvfdxouM4VY8ZX3KkfjYbMQDcXKylJ1ceD
mIKlHRgJU/TdPF1dKHDCWOV8X7UQdnINuSGrxcurOBOt3Ifg3dpsq17UMFEm0zBF
9Btyb2qN0vKhmPn/UqcLbGR+fIhzYP14K+fjElw2jIjsVKW5MQqfTjQU36TcpEHA
s8zNwyAxPpGXlNEd7Lovc1VyawFBt4LIQCAsI3PvyfkQxv5dxmbU/2DcUyw2Oqed
ediIUH8gVFwfQmKnruZ5qEiw+xp5GMFtCJMO32qaFgjCooMgKizg3BfzKDSUnay1
MSPf/CfcFFRM6Nb38FHKP7KtFis5M8wN30IvX4en1FTxP1rw59xKdUDsVunVYpD8
wJNSGX/7w7ic3ITXr/LkTPOFo4rBKOEy+/VtL+qdovW18CCtGBYtE1JU8yZ2R1zI
3d+orPRp6y1VrDruT7zASaFeiSwf9akku64yVntOptF5rlN/9CIiL+ZPwOvDZCFp
OmhQvRhUBkDdH5qG4zsSfDOLYmlI2I+JisXR7y7Mgka4/CgjWt3FG/rvTJMQD4go
+cltUvIkCeNmSQriCMSM58YqnH0Rh82x6ezgMi8Xzv7uWdl1Vy2wO0BNVDI3LC3p
3AmqkzyN64gE45/rLgW9u1WiJP419sWjl5XAcfxHffJgyZgAquKRLSovzK3eH66e
KWcfLj6X9FB63e5E/02EE1XLLKkMEtE9BKZaM5UAxOYpFS72Ga9HfEadijS2AqzN
3a/dwwociPh+JAJrT1ZiTBAF36F+knr5F98yh9+lx7WW8WFVNNPmsbJfsar7hPuL
3TibJc9TArO5u1omcDOAK1nkz8W9pEeFkV/12wgE1rUfTbN54dDbMwceIXeEi7Yx
jpXdjkZUolHDTmPBi61h310+kJ9c+6TVOYlKyD1yGpPykRHfqpmHTUsK4ixkCOHl
vk39GVAlyJgu+d2ybsjGbWmISBp5NsfS+X+ASNc1N1xDtKQ7YBnp25TCFgrmWPA3
9rFGwIUMqvrw22PGs2maeUDNuv0qGZOBOX5naNAaMVPWxgCVUBuG0nLMlTHQTwZq
qwPbH7G+R20rmd8FECn3/r5KSGQpcYx8S4Ub6tW4fZg7ncqYuooTClUdbjQYfQP9
jAZfFARSBrlHAGZE7LqJMx7achFJK61jm4vYgg1MXRK6AFaWttUZJOid0rcvmoNc
Tsff6aEboIa/skL/Sg74WsKZZkvFPWuvBvdH3OgbfjLXcvTbXlkwO0owWioa5otf
kYNL30Kfx6kQoHGgMCDRExMHf5AX1Qp5HI9yhL7cPuoNxac/Q3EpahrAfhvymXHh
YmTDXI4gga1sGvwhzUX8tAbMWPrEYK4+VWWf+xTaPCKVfnXA2AnOGVxrDW6GGyXx
nTcCATYp0ki/BQL1VrMVX96GCOvW9+cyiaGWj7Nos0mkfOBKSF32UNujQDZFNCSy
Z7TT3VjLVpV9CkNA6A+05K9Q8hUVXxLnZE9GI2/3vY4vTI5RyUCBnrL3uHfGhqIq
TSmrtkrB6EznfdlPfNCpBwsWZFin/E7z6q+8DARILFIgQLc8yJpClCUC6aEMfWMM
Orts9JgYdKL6ibZc7ZBwlsFMgNJ4jP/XpMcvzTi7DVbIuUHy+4WIV75D892meOg/
2OBjxfeqPhPsrb3OQEPBwp98k5kHtUF56HWqvGEepNMqkdGh5iW/iG5Bh9SYpBxu
NYAzojqjuWD5QY6AqgO4hrrWzjRUeDyCcNvzNJ/0igwrquXbnWP4tgySeqYsCC73
qwJxjqFHy8sqJ/FY373v/vbqAAOBI+RTwUGM+U+68JSqzlj6QQzJjI7G/JCs30Ec
hkOeihStPnP+VAT6iZyqY7mclI19/z80rZbkcf7lWDaV3Sg6A2AqnagtbhZzw2k0
U0NPSOAssJk4RFta6WJUuGbqphWCPe2uMCVZp68nAsWyXcSHDGbDtYPJlbFsD017
57+YS8xp9FRWnTg2bmjKYKo7dsxmAnzbhzof09FTG/kLENAu4W9rXAzkHej8Zw/v
kW0OsszzU7y2zo/We7JlYf9OYAZlsnUfP92AFXa/HnPzmLEzDdqW4wjCKGLCr8DE
67Zg8vtm6ENy86pIjzwSPL8nj623KylFLYjFpBdmyQ66BsjXOXkxkGAZ3oG1L1QT
I1GO6JvBulpsabfm1Pi+YXPmTx+W2fo3DvCBnXjwL6cwUt0eY6EiD/Xbw80oHerv
5I/FYPh/LOeLgAhcSdAFetVeb270D6T/s2/L0CLrcCanGWowIp57RBzwsb2XFKVT
QIPXxyq+NUQdGaSEWsSL4OLuEquXqU0AoqbsrG/eavHKd8dHKgxKsXKUEx24xoFt
n7udgxbk+nHlshmAr9AlQHfVDGylKLtsc28RyaLLkDfZKW0FtgBpQbb18/3TPPj/
T84Ux0CLzHrwI0OXlkWvQSvB7Qy8VNj3vxYcTbCEiV0txfE2RS/lYyyXk3RorDXR
xohm0PpHkXZv/Li2THd7pk74eElbLiyJue4b1KOspfDmqWOm1ow7mY8Ah1+4xwI6
3d19zLwT+lC4Je57e/FtkrCP7hKgwIRX8fbpuBOoRSS0Osp1jqjlC9jREKPjAotx
rxmtUkMHt2fHyS6sZ4+8KdLcHr8oCTfdYnXdzPWJ/j/zyuZCE7v1lpXXx4dU0Kt2
y9FitPJi2VHMGvUM09PeKmf9jO+5AAhN7XYmS6Jw89v473TdYj0V6DxxahGzIUZt
LrOuwSNw24a++5k42xNcALYMcp8JDyDP2+M5qUZS/eZbWUDlzpFvRjk4P7Leltkc
IYGGRfwzPti++HYng8ojeqgmL+lp+TvcNGct9QhFpvD0DYXaS55511yoJZEgfzKJ
Jse8zY1JbOvBFVqCUAXT5u2PJUTA+O5CcU+tCEg13LPc1RjzanNe8Uv677MBP9zZ
wqGlLGySGkCNf6iNJlnmkWtIzudddWMfvqknjg6tPfmkHa7Usnvwqss5MtWxSWYF
zlxVvLN8cD/TlvBum517f6RLcg8OA1zhTjFd4CsGSSR6TnA/bpV9bX/ZUBvq8yDF
Z2XrWeJvpZnzl6KJtlQ46XCUilBvZdofltzjnVREdgVEj2zxbmXwwSFyPABJb19O
ngH9zCfLB5rkFQbe/C+fLxBb+asJZNCU0V25CEuXihxDl8lz+4XOgygGsAfG1/ua
z9NO4GJ1aWos7j9QOx3KRucCdeU2P/S5C5i2Cpr/dZ+7//Turyk8m57oVEsJ/YEB
smVkWoq/GPsqTn866mRHXROlBvTIk3eZXkusalc/GV/1RdFNoN3ABe+uU6Dyhrcy
mF8mympvy1s8PHohFYodaB0bc5bYwXWqY3kyx6bifkkb3HRYMY3KMW9oHr3ODOTr
/FDwgsnbVxkdcGOEGZAmPlONE/t6+YmJdnhNOZ1oGdYLFjoB3zxigH9htgj6AC8f
Xc4IqRbKCC8YlrLlcBmjWlhHn9C+ib0w3ncc/4uAY/p9U0ZOLZIapoQonA5pxzXm
qd2MxNRnzO6I/jTjDsUTRFrAsM/RY+TUSjJm8amrosirrJJ2Ix8qGx9hbV5eb52Y
ZSA0vcX8bC84p0BD9brsYnBI1sTs8sxf2dv7It+zEj59AdQBCxlUfX3RusPwqMjk
9l0G030BNblXD+8YzvulIsdIvpjLNaymj277y/RfIDNf03qpr9X0GzeleoxPZ9x4
2/pAFoB5Pvxlk5Yrl8p4T+8y12L9hHKQEIUO067dGqZxSm4/ZGsiRvzd+QZlalYT
TrXCH9iqJJXz6WDL0I3quitR1rTiqglbTZU/DfpzdCaHr8cJlZ9YK1bDMQ3bbIqN
GulkAsCNkHb8hgQpR1h+kbL8OnlRVfAJZiRiVexEtaxIhIqPqxXThH8/PN7WkxyT
CRL6A3lWWknlBNZdHlRW1Ho7cSNAHi3stcz02d8Y142VnrFjedD9E+wlTWTtgQ7+
lstytubeSiQCsDXHQsAgKlzMEMwCUtLrPc0SHiq8HryDATPapzwM4ahwZ1N2dJz3
qIagzzo0zfUAH1v0LimE3NX/tIl0s2SBF25KExTLoyRB1cjX/d+oCB+Hd98NBJTQ
zHv3mN2aEJIap4gJPa+YZ3P/FmLNK/5agjUfsg0x6Uo2sjHq9g2A4PGfPTy7mrpM
MDrwshqxBIoIzL31H75mcRhED5rtYKp3DYyNpMFMycs4nFmcbiBqLMeJiQKdWSBM
l8zyg8IwbPXtoA+noRSOP3c3b3WsLz1qdKJcdVKqsiRlwby98/MZvrosPqcrizOL
46gytWyTaF2f2m6kPo5ZOgukpoxMObED9Jm95k9fM9flnH638/4stnLfEke7Kd+H
k1tpKH9k2RVWJ+jm3eY6xgSfF+xEWdlV1NOjmQ9kVB/dvL2n7ptRMOW+B8rt7K/A
4lzAGg5cJCPEbtLtuJ6yrY8upXOzO1nXu1POzJfb/ItZZsVEg7Rfg5qvnA/gG+O2
Hce9jM/NA/8HRmWzZDkl4CwenAXbUQNd13xuS2i4f1Hc9V6ESWpOWapHZQ9EVdJY
+Qrx6z1bPvdcChFxr8QH2u825vh7MzAibGFLoS9pfQtsJ/dlfoxSmVeQICgVucas
3xNfD1ytfwD+kkR0wz+ay3a1GbjdIEYJrAhjZOfyv3IXPxkDvQXZmUjtmLthiHkp
WafMvyvR2oDHE2VoZmbXxswZi0WbcOUwnMgSL5VxO7kWcAbeiNESS1QvyFTUSq8V
2bXV+eLtajOxwbQ5ohWgv/ymyW7qv/rTWq7dD6Y9hF7vkvULMNDQVMGhC29rfebf
oqrCaAX0fCeIXE93bnuwxSKuv75gcXtWAFxWK0xM/kHywArJfeAFlDuOMKKHHSMP
rBiKA+S7A7sKn1Yr8hRjJZynIk/iVcfbGJtaj2xyw4oelKY7VxWjHyvcZfViULf2
/zXABuXqlDT4R0zqAgzoLnXQ4dS8mtQe0CPKPpqoTDRQOH+do2YdlkxYhVVyLZ+u
dHkWrdH+TPmF1iDCeUhKlUFwqdYhD4scBvNwyUsaIlxzKUVLYLPcvSC2H+SdU/3j
B/04FC8MBZsfHcuOQR9YEqEtzoHrW4zUNEwyP7Jejw+22qdXmQqaYqyPhEglPDbR
XJcXXurHRbAE6NSCNAU6yY36Ct2MySR4LUGJiJaefrvMHzhsi1JwvYc+0BmGecbp
LN8ftIKexqlYnw5qSm/PQgVhsE+yofmL8h7CsMg+WYTjuk2/LZBNKks2EMpIZ2VG
AXJRC37RRVJfjwBMsLKfsNZP7BIDAIP8II37lxddwEWl4W7bTbM+jO1mOQbDTDyQ
25l0MunxR1fq8AfxtSgghNlfc8gQsorMzA0hvZj80xONgPQ9tVCAmkh/ibcdqM0j
QW/Zf6BC+PJiOzJNjp0XoCOcbvMgq3LPtD8W90VQiDQnNaJTOri1uOqzNAfdmjUl
xqcMgxx2Ls3dDL7gM0k+xOUNQS+oXLCVQnHERDqzu03fb/QWRLXe/ByR972uAYvQ
7owF8poWY9hnt9ROw5xgofFr6EH3Pz2RSsAtnzG4K8PTAlNxGcQ+rWbmMiB/wxQb
jPZJruhZNbnnqX45/05FOaRr0F2KS9s6kxSzDXopKGOyPQ4YWOCBF70luKoVqkI2
a2VhgMsuzhY4/N4rOLGKK7s1ZvYCt06wy74M+e0/dj712+4q0PJrCqFd+nO6OcfQ
Ol8IntcuwZmFjsRuIAr96EDohfULBn1bpE7ZSgSWjRjvwxI4FB+Y2WEAh9VIMb3z
rjdqV9hZkisJepKiPvlJ9D2DltD0MaK+j4+hLwFDlE4HVL982ZmfreCfstHjRl8R
KMXstKYrLuW9KTHnfODivLj7KBW5K0JDS6bcvh3caUY1D2NMeUcembWkMjIJM4Kn
XUIpku0GtWtv+3twNI7jAp/K0V5NO7gcXjeIAYm9GIBuO5crffAoGt2VX1e79CJt
I9ymRi1mvKQV1xJRq2cYHg7c6gU+VxL3dKSdE5aGVzsAIt3npzKnIQDK5ZmWjnnz
B3XLPDA57h7FjGobIicEXzjQdmiTttdzqyB98IQFxil8yLHKqyEyd9uurzowZrvC
cyeUfRuwykWsGmsGwSWXIpnukQNOZ5FJQQZbQfelK3wTRvlt4qp2+C7PXqqYwD9K
ZwMRc1vSfTJBJkKv1Oes0ah4MV0L1M++/GYQj3zHGp/SJWUdwJNlH7alvu9W1BFT
8qEL7zIzde3KokzehKIj1WyulzwZ+c+G9DMPMZY+02BRTblKnnNW06kK3WRKiCM1
5vzN6GuwrJ7NmpInGaxx17FOYhDRF+u/5viQi7ShWcweRUyTYtROhDuC+uEkx02d
cmXjHQ+IDHf/rGKixvvRiFHFcexb5nsAy90GBpXPkoSvnzOQ4I8hbE0TPwYo2ot8
IlDevW24Gr9mQuZeA6s4hpnMw7uC/p4J7r21e13VhwpAfyr84e66BqiJl81BIz1H
6DmVOpxWPsXZRhuotaLLhQ8Vmi8E1VmmB+BQXLY6EtnkUrlMG9lIPFJagSAbAcZz
gWhhQP+si2l0FKmtBsoHrkOQl+YeG20rlc500jJ+qocLEpxovNc4IWiNcA/XEuux
5AnbnIiKU7HMLccS8ZoSyzEEWWW7GoipAqoYxAFxeUspvx9EFDard4rzNUSJKPMn
UJkIPr1h7/1Qk2QxKfYIPG7F+AELE517czDniWSBrjWe3Co2cLD/QOH+0DhoAdQG
M4m0C8PJiVGGzd7bCMmR4gTH5hQr6d5Jb7YSnu1EskpbtXXiCxpqEm3egm43kFDc
EbOaQqrn5oq5xGytGl2Ouz2Hvwk6O80kx1W38mhdt02PbZ52S8TjliTUM4bLYaVu
PuPQLm2T6rOCmjS+sIbyauSVW8fQI1s3VXSp4TECt0l2xrw1zrb8Z1Fiz/RxBx83
ILP5wAYmMGD2SpKHSMZQRvNcmxXmYq7qt7sMAuNh0Iow6Ic4kpQ01/v1hBm4k1Fp
5XgJOKgT4uWJPzSC1Hp8xoeg0onVEqAiuzZ+MRkjRH2Lqge++sC1k3dGOERZYbp+
zdpIUMFckPoxhqT+iEY0TXmET4lD2M7oAml+XGTdoh0RUQ4WSr8PLZE9nc7GHl8h
iZXh5np7SovggHwikx0b3pseqHXhgDp2yh4Bwg8ui/qyxmLPoRFiGTaHcCUl7SqC
cI7xFM7GK8xqTrddJvrQEQi3rSFMfu6b+8jwvdDpeIiKfrnTlKx0vuOB82sLYsvJ
Y+1fexo0nS++iLTKvDJCowHltBcJYu/rR8qzNfusOIuKY16vkVD0NAQwFXSnVxA/
F7mouCxhGLjBQbSbTTY42ZtQNlnb6WoeqzLOmD0t2S3Tu0cdBBNcs13hV/7ngamJ
cpFR46kUaVJEl0HsIbsJmiUcpKxrx0ZM3BnX6wtNeTcH5rijcjPTY1box5xW+qBr
qHz9/irVIlmtTqHMfxvDpMPJhMB2/VBUApgUHjKvqU2Mg9Gdbebl8VaPJV9PDQsl
ekplqcJmyreZeu8onHZzOU8fTACds29+tNcgtWmiH0nC+UVKsC5ZldCNTl3X53R7
oI4a5Tac50I01NNuiCJ+WeyUJ0avnLClig92K5DiIDHOB4C9LfHfgkKi18PveUH3
tkSyQHpoD64pGiFimduuMs4f6D93hBF4cdchIa2pJVBrNHuEVObGJV0e0Bn9RkGl
uKD1aUTR3Xuzfpg0b7tRPXOASJ+DLhkA8m5QZQuBFhV7l0gYJ1iJZkbGyEN7S2lk
0Cuvu1KES+2+wxRh3h+5N95Fem0ZpTeoduArS4h249NV/g2affd0YM/0Zwx1rwVT
+tOfQZV/62oishSR5QtjV7SAWqbRyYT+d8q79ztcmyiMKEq4h47FScEnLHSs8UQX
HLLw+udSjbyMDYYgjeP6i5/fRJ95kPpuJ767jAp9jK4pnGgMT7NSbj8K+F2jxTYa
6VnK9hVEVo4HTv2Dy3hWo46elfccRIg0OzNqbyh+MkR/OAhhiWPvRkIMQBPNQCj8
lqCKcdOQZlylpnMxnZ3SchWvIKOtCwHp9Z2LQ51hiR4/+h6V8Z6LpNTzkbtQOU34
s54HDZWgpATlvasmqy3ZBtJIvsnHPXGdIzUEnLynQaZO8cml5+i1NTDPfocxM9se
HTnzhP11sVj8hwJMKfIPp2epd5fphSKFg/XeAXiyIx6UhrZ+3lPgDTJhtvd5U9Ks
Rcz+y1yWjJDzzFATTVCMJMiGDlT1JdsjfVBzjPu5V9Qk/f75xjEZXyzTiuoSp9AF
l1IDAzFA+XxB0RpN2N/py7WgFFsZeY+A+CYXrFHoRF9DCZpjv7NCqyMXwVznmwVW
+vtEcHliIbbrC62BHDfcv7bEAN22Lyg67Pk3u4fmT6/csj5/nxK2UrWNpB1p5KfS
wYW/XnaOQNRulX/ZDkai0irh4Xzmq1ArECPVvNgo+wJXvOwMcTQ0Yw8knfa3YwoJ
+YBj/n1yXvXlQ2/pYnWaPZdWy5ul6vn3qpWQpY1U4HGiKBbhHJMN7PZ4HtK2qCRA
oMP9UQTRYdQxa9rqDoI70Y75SQ+zljyFe2mLRfz/WHQUjSJLnOHVP6l53yb7XGVW
M+Lfr+inP6KsK+I+IFCkClUf8uWPVD3yqZiCcR+XqS34bpQGrr8kuQriLrdvkavG
abIMq8rBDKXgAedqyCaZtThjy47IVLEewjAzxG6B2HfFUM81jL9NlCEgMSAL46ob
DLr7jB/vPXAbdCd5+BMxFRbMnK0VH1tGyIH6mvRqd1x9iHrBChHbup6WpNRX0Ilg
3QXY21PsA/hD66vL/SJP3LL+8+a/8PI0T+mQCUhojtJbqBBsY9e6YbKuWj4C4njH
S2PGzbaVUPgBwmKPSE0nOrqN+Fsru9+sst2+oLFGc00D67oYdoi+7TGmDVEKg9Cb
pg/BZGIPzW4EDL4nmtPp4hd1H/q5fCYH/kiwkO7lhX42qbNFN46/nFJta12AWGz4
X2RnH5Y5rvvGQvJsUBHJ1Y7cfNOzSpyvo3Tws+imPrgUpXT533pVoqrRzx5UMTTq
C5amIZ+Hh2SY+T7e7/nM5rFVpKPndR9f5B3wWy8NmYy+rGPIr8n6Q2K6M68tz55h
JSYw9YQBrdA5Zbcav9kUbxeNXnxg+rVkZVKPc4FVfAn16Mput6eJZUKF8lpC1qoa
9ucukQSuHW5qwxe2ccxSdaXoLCx28BFHFOg3cDOaYsKzU+zWsOGymrron30DBljT
leohdYcYtcS1KHEkad/FXk15ABdq454HjP4PuintlVaiBXQV13ICAUGvmocNFCzI
bhYqtapIennswCFsHCZDLEfpr2PLgrrlERVH2f9Rl6FP35oFPpYjv8SZG3kjjsF9
6UBnHJeLdhHLLv4KWaSWov3eCo2H7HWVtMlYebwfjvDrMP5cn83h7KCHc5DiBqxr
4/tNaqMZJShvdw6U90omjwffXdpB+9zKq+/XDK6FHvSXmitS4GuApRXKBpvgpLfP
bj8tO+E3h5MlO0mVyEPrnIR3HBZ8zRIbpUS6BJ9Zlm6hvzRHI0Ig8MYsY4ValcIC
2nNRfGN2u9iG15btYjlLaBcN3IYRg8fJhncMRMwAx19pi7j9ZnI4bu8T1NAJfTVi
6OZuDXHEz8UFqQctBJpc6Uj8uJMoogujsQOGYHbFNYO6U2R0E4ijR6JdSwSLLM9y
NzG6KQpIc+rPIjD03jMeLHKEIwOcEmgQlq1vpupLUsQQplT1tPlkQ1O55B1Zvp/R
jfn3l27FskVxUkws0CZ3OLlKvDiABlfkUY/zaAhBHJEbjm4CGVKe0chDxnc9elEM
yO+abm3QqnbzPUWvXVIDSok3Al5EEh4CvijKyxa4Vjp9jaN5Dp82ppKr7k9WLH/g
G48dLU+O7+KwJvcQ5GJt0LKv39aW51qsoYC0VTQNy3eK8hZag5LjVrnmnPpRDhfg
ujskkA/Ny8IFUS0wfeZcwQT3VyuLSPipa3myhOAApsG4YJYOA8jc0rorR/uV1i0R
rAA1eRmMeHYNFu7ZVjHrRirfTYur2PbKwIQZGF3F797iBOyH+nrHZxIrUAP3Imuq
oYFTNdiswKy2C63lMZdnPbCocfJL6j3FWcWbOrFdsIsdvikI8s0fZfEOU+9qbqag
vi9dg2ringBRcmCZrlBnMxJAO5vSJj303xTVActqEjK0GKzDAut8KL70V7cFueUw
QvUvYlcchzkCkg8ICXfuGQo94mnvLzBrf3Y2pr2SzulbC5CNKiKohxnDpylRUjCs
ZTMFgMx56AE7OJRemeh9nhBpftVbI60aXxzORtvvp5t256yFOnFBFdYLmrNIogJM
jaDWDxhFcz+G7Ubui1a6n63gRWDZqlx3xPvxLLsOmGRg4by/XJ7Z/oHoC7T2KuCS
rtIQNrluBPe0wdHGsE8lLVbihwhvFX+h2UamcRxAHY0cLQnm6f/a2JGOmuN5nd3P
ZwkdQfQPohDICRgq5qHoNKqr7TknnrYNNsXljaiP4I2NsRWH0/IkyPj5dq5BhxCZ
6WV8zP03UUv4iIHwMQRwX4SFjv0KOEiSatSZZjVTE5LY3ONMhwr649iVHrQZl2RP
FM0L7GhYWFz3FH5ICKeJBoOVJuGpFc4pXq6bXE96O9SUH+VyW0kAeHGTQGvTHH+x
IO2wmZGnG2YrcQ8vS4bH7V744zwLyJbbiSFBVpxi+f+hWvVA2V0UddBF9aGVTneq
0LCU5BfZscu+INqQlqYUlLMDqFJJFoaQjL6zIKU8bdXm9b4PUC2luZHBwAjkRRMO
POrBD/IRNfprE5QWPe0V1h5KrJGg5bkJgsFzeMxe68BvzUhbIOXRdIMlvy8ZFJx9
UG5RSNNtlzjwbceB7s8vvY2okKXsRbwEThQQCf7rrDZYfAgjRPm28Nn9UtXmoAlt
fk+36Y/xudc5lzULDvprSYoW6aquMvib3A+u4exmhHxcVqFwdzcu7TSJM5+EspjZ
4Jtqjo2GgUVqBXDY7YJdk9lgQ4BZ11DBsyktLyfoRmLbHA77fybk8oCn7inJGlU2
lQWEvLaL//OkofYnLkCDdHvz4j3iKGx0sangGCzRM+S/Fq225kRxoqyFQ24wNryQ
FYZ/GvAi2fQQVgu5MW5r615DJw1V7XfoY6OKJEkEuAwWJocrXGmiBVu5bahEHfF4
aZiuo5KPVP7XwMLpgceqwpQAIwi16UVMIswpsT8NZOOnpawoIAGv0cksPfYfpgl4
ugJ2yQ+MiDMvSNrtKx8bEL4cqK/4ZOPHWU2QlvfzEYU1xtQTVcikInlkIyIRRwqR
jUIdZk5/Jw2T8spF9KCGaHsSBrSsv5i+t0AxZqadag6I3BEYfGoU13zN7qGY4YjU
T3gMHcoCeMM1k1JSSwar/GL7mbGE2xm4clgzIDrpI20Wz4wdESCcr4HNuJJXXgV+
3Kd76tyHeaQQBzZASgRjY0eo6C/whbMqd9mVpzQ0Zmzsyhenw3DFprNaZVVo/6XL
7NyoyX093p0S+u89lepeo426hCBTMBIMIAxZXEP312PUjYOWYcrhUZL4V4bGyZuI
vJ5WzBZhpvm0VoK+OoyGLYGk+qaPQgLKVE1uUBIpUPfTkrxQIRjYwNn5mCr/8Ilb
74tKUIfbscnpSMlMCw8NTaKM8UBnetCTnZfg3CH0rv1L+PMafX7TIgMoZAR9Hf5R
6oYW5VxSkjWUPB9Ro00MMM23Qy9BDtnRKrrQ3VOQ0R/IQsqcZKw2wFp31fnSM1An
HM285gNh2icBL43uQGKiSFxFlC+Kpmjjf3eLBzziUQyfSmGn+Ysiby22mwFu9Ys/
20Go+zSW1NWfgQHumvtxNHL6zql57hBKu9oBc8oOIO1rKvmmeQFmYW+pyvPZ4hsC
DgKY4l/imAIKiUUptABbdqjbSXQb+6v5yPZy2jSfTxjTcmlHwVEx4b41Ro8R7MRb
dcQj0+L58ozGUSx17ZwHICnS3uvk5ntrnzxr35XIsyc2+hxC86XZ8QRs77+MK2iL
+cyx8nZIJMhYb+GvQ5UbRR/iuxNFKBkXvlk2aM1E6MxDrz0VTvfxHi8nPmDAtHPo
1Xl+r0cON9eDZ5sL7/4lQA8qzfPbE18IgChmmNeNOz7YNqRuN0wzpJsh8zPohWJ6
7rX5yPdMG6kfmuxVs63biekuw865XRDjkJu32yCU3QwsVVO3pbKNm2B/T5XOEClA
7aMC8898hrxoFT0aGBgzmj5WFb/U6AJ66058zw7vK+f6Fk4LdmCV4TaGcDaDVoRz
buLT/cdqYpDxhtg5aLI8mCqxO5PHLJBpO4gfqy6kZzNRKOqjGGm7uUoBP0L8Rh/h
ptXtyyw6KghfHaFwAH38hL+cqnXNK/ZGzGzRp5wH7HAYX1jfnMoy6DALyv6EkaDg
whDnqjpJtM5QOPw7qFuJADbVeRvjzj+KjdG+y2/xSLxVMOxHI8dDhj/LKpFWLuxC
DuEQkuNmF76UW39352j1mm43nWqvZ5nA3nsUu0eMFocb3BNcZrIvDHt2gyJY3etr
2HpiCRmEXlihITwYU0xVeNxhH+nJd91H2rp3YaWHrtpBsPC2D69a8XSpRYyx8LDk
thlV/BVP4+eXU1zgEPDmLdgx7MqMkGsCuGS8bn5WW/MVRPjNEv1GiGshQCl+I3Ht
nGf05Ci1jbrOeds6ZGU0TdHtpBq1rhEW2BP5bORZYP5V+wv/5nVfc8lob4+T7wnj
o5DJUW4/MO4tCyrCdYn9pXkXxDI0n703t+m00Ab9KaHcZa2KubWUMJuBMGso+Eq9
At/DPbmTPLv5nn7WCCLAPfJ/O1WrV4MC/7lIrg9e5e8k2sTJ5JOTRntwBEal7ta7
3NrzuvwCLZdXsZKrdf2lGNuxsIeKdPBrqLVa3/rlI5TMj57cNk1pUA6cQ7xOlJJw
egkc81LhWxYLVtPvfjiwAeu4owycZLes81aceI3srwIar5qkpRtYokoG8/PWcHph
7ol3Akl4vE5sxD4lhMIlOMrKlzp3KhhHuhOPPukD126v3tyx4oC4N8uuTqNeYLGn
JjxzS9QUkrsJk3Hrq+2rc6UFze0QuA1lR595gVNUCCn0YnbxlR/DdgzO9OibZryb
404DiMuCvb4Ma63kY4WDA72mEcBreF+SgzEH1fEDsQiS3LYS2UezZ1n+sdR9vsWV
p1g4JBBCR5iDpT8+FvdaCaPhjC+QAjhPebUhjRh/RNvspHpCL43U3TGRBtmCRsP3
Cr6hY1432qD3Z+SDfatsWCrlmk9A7w4fLDM3XepNcAmxuAmi5qXK3E9rvLneD9+W
ikQC/wuBet3jVjnD2eBRZXJpeQucspA4y68wmOS86BUK2Qcjp094P+wQVn60ARaf
QpBGHzX/Sb5fzrm/ccF2R/DPGr6a9MBH9iR58cqUXKWcGoE2+ATUQ0+U5OEFvF60
1ri6klO5eaCkYpBynih8LO4GPxUi1qf3g7B+9MYuzhVsxDj7r6zYmc1CDHg7Bsog
t0DL8LLqh5mItV4ro0zQ3XuptHyhplA4wZC+NF9hdePcpinY/n53V3C3njOmi0Uq
Ed65HsVvq3BGP1ucvM3YOrSObqWd8fajF5Lrh+Bk5vAAkJRMUN0Lo+Y47aL6xaDm
jaGH2cAW195Ri05Il5DxnCHflfRG0D79CgB5QfCiYIreFyeRxSpY7AOvN1/2zXdb
XPgHVZMID4N+rd+lRF/N6QZLbf6J426451bE2jlEn16GE04Nn3mnXv+clx1Zk5Z3
1whMT8eGUZYjjxzG0zFi/pba07sIEmdH+Oz9ky/V0h3Z3angvBhaHlM3fL3CkrD6
VoPiOn7JxHV0AWnBLyWmgSlLA+9st6U8sCRWsJb25Tv7BabIImmHNmEUdD2UWibc
ybL3ylSXyOdQM6e2NtSGpXRG3WGJYPUY8tbRuv+TT/K1Sa9bXRoM2u/mxPnBST7r
X6p15Dg6v878silbzGnlYn5lltMk4mRk7Jc9I4zkCsttBm4L/R3sJmNgXIBo8rKg
iMK2zFd2dycwO68BMjxSaSrJuoE7M8mjnL1ZmcHg7Jipwdfy4SXS+4/vXQxY9Sbj
Hljs4FEDJtv+NEEiLDpFHB9Kj91cdAZZn+mn5WAW4XLNvvVmI2ZvWDdWA+D7H8QF
KgaOvVhrjWebD2Rp+JBLXszmE98hHysow2NHxpB7IEFdz151j9tmptC3D0xV7/Wt
KbjYLaLAIY971mQ3J+nM8ROqD9Qic5d9pD35Z7gDtYjcGtu3E/IyCivb1MvBkR1g
ZytHpjdINpCLkQo0HrsG9nb/PZQ5wk+Q/8VmHCAE4hpZtgPL/YoHhXoqqX6MmVjn
kZFvioybb+h6/RvgAn4SrrHBkciVHMDBon3BBsnNvUfV3JNy7hMsmvhGYnzO9cGN
3JHcDV4xjmj3Y7MFlscrhDnhedPWyW28xZFRPhID8i6enNaDvTq48BFRoi9vJ8uF
jPNy/JZzLYOpqNYr/OktVFtE/PqBR48jW7UBVeu9FL7lA2BiDNqcYqZ8fqs6oxYm
5A2yP2Tx/8W5a7LDWYD/tgmdd3Hz9oO1sNJiSebThGBrCSH0E1FzriNW3T9Khywq
U9SlHqtMFTGVx95lY7458kVd0mG//JLNSgZ9rVJTe9OAjmArMk7uD63euygyJ3yY
f+MMqi+SMxGq+Ey8r7202iZSTRdjU/Y9Myioe18Eq/48ZQZA6XqnWqd18nSRXdEj
r6zO0F4Z57TwY4GsvhzdjdqCNpOKcBiKz2dkRg2SrMVo8WcHLCd9OO2UuI7qahfP
6FGCfSyh2dlBZNxpe0/LAmwwGditwdFM4lkVZtOyVcHdLutm7emICbgqpbSbpod4
D4nbWvZZIOaa9zpIM6Ceo/dsvr9/GbzOuxQOk/4S/sEEVDdnFuo8hzaKbR2RMKNw
AWY+turNNwGWMVl2XngGxhnhj76OB0NJ44edYL7yE0ilT19bUpASXZcPSYzHvU+R
5qklRXtmd4F3rVg/h7kg29EyfIHO9UIkpkAFIH/r3W+47cfhwl0AjKHrUagWegnn
BA2PbDVwgvZl6+4f/OAJrlucwHr9KRUvQX9h/+hXIU3kfxhJzU+rN5HcO+qQz4g+
9uPcwUJbcARE98IsidYdo3iXAhgav65UWX3Zmnl+L+bEF/Gcy+xvI5hGhK+eYc8h
jAZTYAEz2/gAfX3LtfyoRzlhome93hId1IyG0ZWoF21/h1/dMOFZVA/U3r+E3i9i
a5zjblPU6wwv4X9Rnj71QfqZSVP6xLb9l+JyRpZat9P4tAeR1hZCVhTN+dRcpTze
LzCicyHJZwTSQ9R8qr5W7gbLYOXxj2iZNWAsO6WFxwU6kcgdo/H9V9t++6bQrNFI
D+80IiBOdFJv+4ZWxZd3GyOPO8ocFbVoMMgxfp5DI0/GESrjmYNnq6UsNys/omtB
f4jT6yu7/lRXZWUUt4dDRCJzDNTnr6R2GkNTCaVHffG2pnxjrzt2CVurI5+31M+M
gcPm9PTa/6jyxkwhvp2/ZTxQxu8nWjL2/jFDUWe1dgn4BPO+YZsJu/tRf2mChSOZ
Rq/G0/5PSjg4ULPVIg5F34x4kdVjnBAIvD2yaiEL3VRJ4rRz6gkIZbD30v1azqsg
3Zd0cVarjPPxD/9XCwzs4/yyA3mr5eQeh26vlpXj8NgquWwrreNDcn/V551s7CeM
k2fAZLLv0dnoID425V4NiTaYNAua66NCiIapmJnArqsw/S6s1B2Kht+B+WIFxKt4
8y058HjuEFaLOJRn5mekSCHWKN821enTrqHng+hh9PnWMlCYoA7ify1p4l7O/U6p
L6/KszvmvEjZ6bwEeclC6NpjBz7VRz/9OpQxOHPD58zZKShCdToZ3vQlJuaJoMMl
4oUZSK3FFUCPFnm69ZDn/+a7ChU7/BqoNpcV+d3+xWS2R6N5MDf4YaZ+bZ5OeHR3
78XXg0yAD9xQBMBwy2rPRkd4yrrImVRrP1Y3lU3ltziWwQfaRVWOkZMyd7itcCAP
H1KdHP6sjIGdNqfX3SouqGjjsnNQj9YgmoNEXfoHlpg87RrtAPLBmvTqSb6iaieU
Uudo7S0bCDRScXAK86Ql/k3Wfn0BJgZn5rbWD7QW3opVPy5DY0Yxx3opQ1Xbqp67
bxjNlgpej6Hu9ADJB4ihhFaKJd/JH4y758Z0VLJ4bk3q/uUYX5/kaHvxFqDGl7gg
l6b4Cz8KHMx+AqLGRVc3BXK9WC3rlzoYNAXIXbrGYefv97Qs0dgoVSfkULCmf0+k
T1UQVrAY70+ADpdG1v/1SFe2ymtjQMamqi2oYmoiT2YA64y4yAK/DAcVrPIIXONy
Jm9kFqVrJT6NLuhDYyA0cpV/yZoH7x1EI6Bdqrcd3wqNLozSiYeuyh3BnKBshShR
AIE+osIzw/fPa6W+ki2lecea6dxB7O6zu4lkovWxVTRc7fNHBuPlmTyYbBXwLMFP
xPHMzRsi8IJK3yk2le2mcWU/JFTkZNN6a8WsD5Et3+nwsaNsoggI79ZbooOIRLyd
JUcLzBO9iH7fAyR/PSLDCU7IBAb3ONY97MR0F7p36zgTRXwm8wYK6RSV+cu+6fkX
darmn0tNKuoMCh60Kh0tY2B0dxzr/rc6y8A0OFVL7wbCcdY79KXJ93xXifPJmTTQ
hq1zSy551wJyfyXNIWRyn6ZqUuabrnGuK6zHpDQBzbalQQ7qUcSOhdhO/c1NhCl3
jd5niXmXCuI9nipSy+HU9gPft9Rq7kIUZwoUGyGik3Vv42d2nF94b9RD4v9zK3kE
XQSz0q3hRNT47o1sKZkztgD5mJHJIAwajvZVgSg7sxUIrpUfRHgXjmuqza3wHlk9
sk8+Y7hL7v7g07nrPmoYqLqrQ1dhFf4DbTRdfs//q7grOBAbnvWYylqNOehi03uN
4qAKrafBlMAt1c1rv24j76p5lD/SkMV50LUnX27R6UToEbXY2MKxy+s2fZhFPfsz
enqlPaLY6RKiMM1DDyK6L6e2xjTLPvoIfgqCQwgFJPHOQMxfjQmvgTgs7qfRXvta
nX2BDflzaOk/cHMAd4ONvqeRQo6GOIzKWbpZnEYW9LJGmm8rV7X0qAchwMXlatdY
LpHbYhB7dWZjHqineUSUBcLDmgzDsa101Wz7xpAI54he+lrXJCYSshIf+gIETpT0
YZKA0PyBMcSbIu7f/V+cH7qZWuyzVCySMK3EdxP7TGQyK1wkXJ6XKepTGWa4v9c4
MZDgmSYHuAlN3wApp2EvfPtC8aqnVa0cIUuMKFnO6Vo2LLSRuXL9u51f17jN9klj
J2Yu/GFINjBo/QYJUKJz3CqFiKWLyjmvaOLOlzSx73tf1r0Y1u1EoSypIZH584XC
vVI8OjZBcfWLDcTa2RJtvyu2SUhOnq46uu5xdGy04rxkL7foH/1fA1BwFnuSnM9b
peUdr8o++Sjapbu6+yGt/AR++cfN0zCNQGlcLxWadmLNEbUqh3O8DcAtEIPhgrHG
gldz2cxujIy6NWM7lHUFGcWK7/ZEyetN3o1CxAINQvoM+Ez/sb+fU9mSSliF7UJp
MaZMIpkj1h9hp/ZPkPHOWNNM3sl3FyrDsRYcKSUIoFuLRaN2v9igP8UavLtSG90a
vYHUS8AdEJfrqYHjJ/upD4OqJBelmqeL+zvJCSSHzjx535suY7KTUce1X7p0vn4k
Ap0y74Nlh6HnslV0/HmUd15Ccx9/lZRdPQgH9EMLKavuyKbExk0Amc/w2ZfLpCQQ
coQGl8JY3mK3YIY2/ckl5MkDhblfdzzJ+L4akF4q97ypvhmvSBSQ5l8yk2EJiVT1
1x4NhDRBuj6oLl5MHzlJmWYHf4JCs9Mfdj3nJH3bvvjXEt2zr2byjoqe0+AB+IPI
1gBKBkM5gvSzPVcrUGEer6UaqJ999IYM4H/+5SSjEpdZHUhgW1M0jat7XEtyW/tv
FqSfZvyd8ek7Ogg1ANj0iv9+gGgQxKeV8qusfKgqGoky0V1TAoqCaqJGK17jpNy3
XYMWLnRR/cpu9wd7iiePcsxS2+TJbEoVCxyb04GGkzEIXxhxGGZDb2yiOQMSI9YX
rp8b70Lyy+X3o0rsUd+i0B6ObkGy/or31ONqSVswjV6fMd2+V1ymFZRzQjFyll2l
BZ+yYwvQVeHTRxhzWYtZouxpPs1YMiwnxSeY3o6iLp08UN9m6iMtUgLXWE6UXF8Z
UY4rZ+KMSoidzKjQI8g4OC9RhXjmFs26RNjTUEHZzbhjUBCCUhOe3+owlI3KAj5v
oXDuL+b2yzlrk8ayG7o7RJkZ9bjEeo2bn+wuMQfeR/g5aayRaHUUX69si+zzNxKi
f7aCBmqeYDgxygb4t1CASQMSBvpalbT0ZrgP4AKnhbcEEOtPS47lb+dW9KlJnGkL
BuW+nFUNQvBy2N3wFrQ+aWMlmzbLrJ2zh3phx/zMRnxQ+o/86+rE+PqZeuIaR9HO
XzX8m7ubSpnAhsRfKqEeCZJtN5mWKXo63S8yLLVL298CrwlQtgZqlE5u7oAc15Qb
1xURUawUxfrQ6GiGbqkVVP8RYVgTpejnZ/cqMeVTb9mDuTAzD0bNRztij9PLY4Xk
SJzh1PrIveYPFdLXyIn9T8kvvDZrrBZWhVP7WTc/prpUB9A4JahMmfohTLBSVah0
FBUcxNhIhvabQtrcQD/cOz271pmEGDaGsKUf+74ILdTX/+hu7HaC+UUfDjznNdDg
k4+xgpZj/CxzMqRuX3xL4gsY/Aod9e7x3DkR/NCnKQISNl59+dL8oZa5KjdaZ2qi
KKOF1E78XtAi/cnrozERc55J+N4UE6hztapjxqY0Cxgr4Jb5NQDxKfMwbRinwTmH
KAI1wbr6OpOzX9yJG1W7+9iefnaErAjDlJG35MCao8GnMK1gpXi14Bba/+XZT462
ZZX6TRR1UFmX18CRRsCT7WJsilOi/EGiWOq0+Zmr3Bk82Qleoku39AHa4IzYbESR
6GBMTX3FfM0piY07O71hGwvFgavy0HvfP2zWNGohKFNz7hdjYxDuS2ICgbTH9HkV
1RecQxyMVHdNMsmqKi9hwIATGPt6EevyQQ0i8xTxcTpna+E5rHsvBdon4c/H8aKx
rW6GLjCTWJCJy+gupoCJUOhJOyQ8spInb0h8hvuBjJ9y2qycg/bgtTWo25v14knm
FvtCGTfOsL/A5Plg/ChArehtEAGES6qYyem737w2DBXKJV8s2fxmMhw2AAwcu/kQ
g0hcs+0HCSVo5VeHtiPE0415bwbkKRn8e21DdpYux9zszarxwzu6zCFo2LxiHQko
FGdl+4Fhyn+lTGxeI6FtTbSAc2VkufoAHoreyRSd2c2Y1RPA4+eW9Ts7L417rQb2
WpN+b0k2nefCf9+OUReyoASw9LGm9e7/0/r1q8KZksnfb4YDz0Oi+doDnymY7QCT
FgB7tAHlrjrV6y4fyh1iPkgZOG7LsZDLSAyJj7+JukINMlUd1Lvb/lfjbpkO/YVY
z0fhrGNduKvJVdbDtP9lRpk9ofyaM9zC9dTUrsaemRj7RWMItuhiYuEjU2X63mDZ
Nw0sSvX3Y2mYT1A2hl99XOC7gFOiZC7lBBcXN7neB7fjAywDVQfdRXGHKrNxW9l7
1pazp/k2Go40SfCsKfJwjEAJ8Dx8bqYBJo7VAgdBGazQvZ1MpVCN3gsbwOR1X2Js
qt02TM1nZruVSpAhMhon+ZITO63MHdUw1ORqxzFqbX6cCavSraG0TeUvcBAcsO53
oWezokNV44/qHC73nh51SdelXPz0zooPBSBkQ4JznPyJarp63Cuxipe5LASFq9AS
2LlpL9eQeiQLOyxOeVW2aJM+03aQ4lRBmYqDVUc2ijhanlFYrSkUQ9xH7/0JBLfl
n/ZLeXTxSHOXriW3TH/j20JaImEW5asNEj6Vt16HmUjuCk/OIh2Z8ocp411BJVkl
89lAF/d+6R+l3IDpZR2iYHMX1M9abrJ0O5gsCuXr/F9rX9w8sB2zXOZss/oTjtYD
esDySj4jVI5w3q/WZpuwe9o4/BCopHEH+9wsEEecpVeANA9Mn23ReAu5IqkYXQRq
NuvtH9RTbClcpzEMJPcEwn77Bvm0wB73Ov0Sb1OluOUiR2Jd0yKqVDO7TanR4E2i
+w1LgMTYLS72k6gbQQmZsRYJLtdLz4jVxSZ8zbg2IjwWH/4w3YPTOBlovzuUVPOw
Yuj1M53R4XbUIw163pT4EIU0m22e1OlYKcz5CIFFTer4QNx+GhGLgw9TiHFIcW+b
g+z4i1zr1rtP81q2fohQ38HamUu3zwggQDF00VwdlDp7PGXl9T2cpE7trCsT5yY2
lu5B+laxRqt0K2UCaGJqasam0ZT99cDBAYkC3vvC/MFd00GzehePtmpzg4cf+25k
X/V/yl66BfFTKwl2pJHrGJaYKyKa1h5VN8NdPvq7cVu0maHamkLUdh/bkAGPSpcT
0QmusgG3iB03ruEIThCHDFhErmXbV9xbTe0JyPe8e02TXnW2uCm+d611gH2t+rs0
0xErbRwBz1FfA4pWzru7GcfAX+vjXJKlVDJYpdbXRwZES3EjUoJjsGnq5zYMupM7
Qe69OzStS7eEEYbAE5td7AFdjmSF4e/+EuFrrLrdDL2GegCZdxcMNwYlMp+5MuOp
cM28BItJMIfYE2sCYeIiUHdecPhDe2gGfqcELVM4rMfS8fFUYlJybAHEty3VbQKO
3PICA5Kkhh8JYh7f82XuEb10g45cNUu0KVMTjGoolDCxt34gWZmN2rCH/0tfAktj
XQOzw4Biv9S28gDh4roHlC9G0XwegvHj6VkrcTWFonGNpL7/atPk9Zefv4Wd9p4r
tbp9kD2cbvQi0PdEreBW+Rk02Yxx7m+UBq/ujHG4qIqMyKpv0OfbxinwCMbpvEbA
P3FEbIgAisiuVoPqT+n18uzE8qwedCml7njqtnsNFoMkC1G39ENoXBeTWCt9+BvN
Tnbp6w1eRlF1cwGcmnZDghr+Osmm8OcgF0OIaJRdVORG+eJhhKXqDNcQ39dniK2j
zDPEg0G2hPf3KG2hPP60oB+JPsCDc88QOOGctngtM4eV2ZoXo7qq9rQcl1YRfzTE
PcFnA3rsX0gb6aW7lQx/onQ34a9IB9e1wwfGfWAL/IsDJl9jUQx9LbZKM7l3A4Gs
/6uHEpbsgF4TASygF6JcEK1KBxwwf3iqg9Z21zrHtaBQv+FIJWI7XIS0mvnVHEzm
HISeC/slT8UiKqYMhZNjz1wN5LU86nYexnmdzR7yD31FtEP1pt1CBezAFChFyVdz
Vpqze5FJkGqYBU3F/h0fnnC9SiS/Pb1wQR8xoD2Pkqml85cbQ9oyPxFaAPHrR9vF
QMKF4p/EStjyYy2Xm51s/mIktZBInHhAk9ai7XfKdwk4TePH44uiUrKEesJW/iKB
S6+Eixt1xvmJGfHeFzZF0dbTzswznRAc1IYITzXZQKHeRg5rH7OyavgcNdC4arwJ
QNh/xbTLdn54ZvOBU8CegErYwpjui8i0PUws2mKhWld8gM9qYI49cw8iIPjcK0Zt
uHh0hLEbi10zbG+sFlaaZhZpGj4WtK4CM1Twz5yRa6wY/yLRo7VCR4Xj3dytPdHJ
V5gSAJ7zAr34pNy//xr9jYnfEBEFuSWv2zshC21sEx0eNEKzRB47HOufVDD2+B+L
AmRFD45XaBokMoVApNYkU8xBP5CruYQgsyN790ik8MEOcO20PYWcffgYaTMgnOj6
PwGyq8ByVdABMzCFIOVApwsuguEOPtZ8/cBWTg1fTpTqa+p3VmpzUId0ovSs5GOt
VfoiuiXub33hvrL2mecuMvj8y8fa1RQfogfLyo7rDL8AbAwUyktvFsIHqDooQcGp
opzEckin1/xHKqbsGRBk+3fP2iK5aaiHHpbdXNuoOr5sU+xWCccZMPzKFomGUSGK
GHPZq+dx8UJNEnnjXFsFF7AbOvVevmc2ayF87+rD4UXwLU7JlRi6juoDkojNp68e
wp0Pm+m2vA1WAHnQfZmZLlc06m3v+oAxHAv9Fv8X5yVgV6VH0pjnGjH0DDQaByYm
8atdnq8+im3zY98Jf38khXRx2SOJUMWHBdQL0R2Kf5DR24KlSowxewQLk6o7LdGF
wKkFR84fAQpYVLNNRaVjQFstOty6jEYDXfzNB9x/LuOenKWOuolVwyMRXcEXQVN0
jQqg/jZKHlOO+eyxxVqtIxDDD3aDonmFG1aDIp455G3BLDA9r25KF1/ZnzZboOLR
VL7e/uDIUD1RBzPav7YtmpQ/ucUc1mz66wXlvFM0isaHvVUzIq8t2kUlmr216ceG
p+tXdROfSTDV5eL0IKG1Mb8z8qNh7s27nS4P7GMhRjGHJ6EJFxivhKab+fQooMlJ
iS4GwYc70zgim+RS7QldwXLY3LiwBZ9v3Ax+J+s2TZtt+zpDQgpBrOSmEV+L9V8w
RM91TABkouV/ZphhGmxT5NsX+vQtBdRqmCEH3NJZpxgBUVewV4XFQHUNn8ul9Yiq
LyFPV51qzJx6TLR55OHIYOvGKJzzLFLV/2OC6AfBD7NaB8jKqFScr/y/UQ4avJd9
FRYTC7tXJsagur+fXQleykaiv9UIN/QPGbt4AHj5+ot8YtRPp3BosVITAN+xzxt7
DgrNDi+zBX7MK2//M0NXFsTvfC4v3PK3ep7Iy6B/eY1y7XEeOL1TzN83MNxCt/XB
RLchC+G6bBPLRvAh/32OuXz9Kkq1gbi9NttC2l1PpJJHDRiff8skFvGrOAC2ubFa
cOJ0V7QzRQlUl5IE/xW2WJxOvS/jV6l/+g1m3q0vcnCEm7FFOU46buxdRHGZfyjy
w4T8MojvZfRulWUqMi3789wTBtuhydTf0kmf4aZGw3ROv3NaTyZVYy/DG76IOoJq
Cjt7dcYuezujw8m1fHjsJYk0HPoy2R1S7eyCuzy2Zu86oKkRlVfx8NZO3FuKSTLW
N9/2w/yK7x4lR8aHNwb3E0s6w5/D61FJTz/Qoq/K5NvNLhekePKo0iHDOGoMGyla
oSbReqJJteHIHlSKTkN0YNWn4rztecQpQQ3wMr2/vh3vmzmqnFPggNKOZV1IlEJu
EThbeyAv+SUHpDgleDCxA4j0iUrz9eNGb034Y24EELp8OZF1lQN0l/Jjg0Zfm2DR
iUUppdOMOnrZLJzmX54n77NpA+dnjPlVJCiAu2jws6HRQc/PwvbFl+3D0F5qxamW
abrAw4dT2TrQZq4/yTGf4MPrPtyt+AQapGrKzPoCi6RWeptd7huGqa8aLTedvZU6
Ppt1DIFLp7h7OeChDy1aV0DZIpWXHAnlbwxxGl9Td2hhzi2RXpw1j33fc7cQD7NU
XMqUOZ/vrCwRF4SpuDoZfHPFS0eTgT6kEGCNK4kELZTYc3BTQxrxVadVuzJGrA2I
AYn15l1/SvPwUuVtJ67yJdRdoDMXVJ5XA+Y4s8qUls2e6AIFvrDxppUn4IGQtm60
wwGkAYhg6xcuHPXbE6wtCqlj4g9yflv2V4NMGn/sgR2vcDYHWHQ+mxDvFlwVFkpC
Yn+WQxagVnis/sMtfGXBG6hWE+TpgLsq6oFFJbRlar+CFF45m3PvLO0U7b3V4zEE
gd7E1obULLXEYp3D1MyxMdL0hjEJuE0JKKSNxY+zqiNWi3zIpTOsl4SL2XIksx/C
oY2UaONo/m33HglCjm7OrLkJHjt5vXkx109pACxO0cpv1PwIKRuHY2iSSvU7PtLJ
0RqqWoCCDRi3Hvgh/NEq3+4Q+6uoyO9xhqKjI8gGJD3b5JAFnp7XUl6CQjWar2X9
M/WU3kZuO+5hOByNIm7kHYZUU3PpuOY0YtDUcLfGagFdYgUoGa0h1Pw7kyZo+ylu
0r1rKDpiD3PvEXssCvIEPnpjzL56y70/COlSrB2whj1+SACcrJr+u3Zr9tCAU1Ms
t3qme59vLlZ4eOhw+9NTVuzffrd4cbcaJX0KHp6RvwybzBwESh95Gq3i6qZAkdEc
xm7EO5TT7MEtKfG13QKOIWfRgXaYBcBd2kwUZ534UlHCGf9ra+FB/erd54nyBmXm
JFBM/rWOsRpnLQscKOnhMigQq0iUF7Ch4/qoQWwOZ5o1Dcs8xXuu8glUYXTbJbcX
PLydzmWyGxVXCys2ITfX/ahIu6hXe3AKbklNHmiMOLDNAH0bNWcL61BJmtvu83le
5MMf1FjjBWY9sUUrLMM7vOBUWUwj6h04G5ghvA+B1zhy4pjiQnpnK/jzPGpWQSEc
MV13zPX8BZC8kW6fKzbjUapMS1nLpoSpcvSMOgj20GDO5WzG9hSc/6VHvhmr7Tgz
K2l23YHmSllYXGQfPkECibLbHN06gRRxxZqp8GqPBJQjHxoukyj60fkJos2u0RaK
Hlcf+XSetJKU1IkXUX0iP5nQr4d3M6DecBNQ1XD6ROi9WRFUXwwUJomB1JEaZ0ai
B8S9+o8fAPlqHcrJOoSISjKYMtW5fMcTwnsNMGHlI6YnW1SNlWKSNRHJdbZD2HvQ
MiPx+7RAAA3C17hGx1tbkPvEWXlMYc36Bmlajl3HTbQzYJcfUNJc4HgeATNI9yzU
fP8TKYzT/4WbySxtFSM5IVdfOfRAN+KncKBHNVm3CixJEntHO3eg8Y62gBLspjUQ
B3azBnDkyLoNyRTrdEE9yp+tHrAwZIL5BigZFl1o/Bnr7uQHiFz9K9l0BFdsJYaY
i6PS4Pn4EALl7xm1JfI36miu4Lt2R9vsWrLCGBxur/jWrisYw0PCyJcrpYwYPuJn
UhREItMgUk2W0eXsx4p2tcSgM7rmI6eH88ObGb08P5da9Ug7shNSMVZ1uUPwY5pw
yO/4tTpB8fHkZZsQu6yk3fWxg4aNq4Mt2e3r30kkVCKH760QgYIZRBgKdCzC5QQS
KidG92jfgHOmgWZ+kF3UrjE4JSJ3BC53HpFN/BWrFAwAnRbMoi2hLmwjRUWaRKmq
gnR3LFlwiIdXH5CeXWrKP6wqw/cmY5+7Qk9S8IIp+JXyKOaV0eTo9PRtFuKBWDuA
l+4dfKjQcNNcZfsh+CIZbcEF0N+hakmeHQqtfhurGQNaeko/FIXmaTVtBZthWcmE
L9pZ9V38QKm8kYaviKK84tZRRfDA2ODSmIcU+mqrZ/4ZiyRTleDzNDTB+qum0Abl
4VPaJQpBN2AAtvTH998XJ9MHQqBZPEsaN4WUYifioQnIrgJZAikQFhoRv8O5Zlat
P1qf2LElHm8vEQH3wox9PwETMi2aHrAB0sKTjY0/3ItHAm6F9ArT4nRMer+OYIrr
zapLpEk/JVMIO9WEuvUAiqbeqDsjlWMF1Ame7W2gllZ4ldJVnVhGlOnitm+Uj34+
iegGazoBAUPsPG/pLFO5bhepkOr286Jf44ljRfnE5r35L9E/OAgT0gpKwDA0oj0m
7ejSj20Zl7dG28uCm30VGXqiTyvop9LB8veaIak3DSvgD61mpeEvrwHJ91PoE5I8
cRKJLJYJ3KipBX3g4CBerW/zJX1Oi5nbED0UwYrYYv7/WEJgash/tpHFsaso3e1j
M+xq+p+QT5nI6Tv3jTMjEzM+hJfNsvgAT4/Gk/WjDIcijfJgieDnxCMT+jWa2iks
aeijRzUGwI0kNUjOH0H2kC4qVMnTxKuK/5SQ31ikr6qvSGKxP0NKoLf4A7vB3942
iuD+YCBa4hL112467u5hriNUzFiFjIFFTSWJCnsNrlYwcTEUItWOUah/9KsNTVt5
kgre9YMOZYzIlikaI/j+gBowBngpCb2bXEGYw5vhv4XOecwUXEgjyzSzQBM6gY4W
XlzMaN3pksDNbAUxT3dXzcP+cQkOdH0zytVjTYr/WWTQTKdpvlSjsDFLmq92j466
fhS0c62O0i0LQE7G1FmgXMi93vYTyUagMtZd8PGOIDwJgOpQBkhQhmDA8rSzibB7
/NxkwpblcWZe8T1+QVWTObmEUTnMdhOlVG3z5moE5An0mSnYJp0r1J29cglyOPhR
KTD/MjcjmW/yh2iVWofrPrhrYdiNhFoWhp2nPByrJZS+GPbUf7N/TKutsSmY/GiE
p3DOodTUHNp2SoZMJjOhJxy44pm5XBXq295AhqiugxfeSjqsIbQFvJxYQ3nq5XgK
kejPT0YiddBG2uXo4D3LNeOGnd8BnICuOTny+hSRan1hcG7Prl6O9k3zWWYrlUnI
Q79AK0L1MhsTUfzuIyrSwVBYES9R5RPql7TqlpyKF77mNsXZPMKpGDTiKB6ka3GK
m8wSMMpp6Q7D2wYKljgWRdYhJHQTeAVGv4I0g8SyLs7jjvVhHs6+B2Z1FIq1+C/B
3VPSJE0Pbo+R3LRhopZwJJezLY+6kxK1q/osC4Uibhg/XR7oARzRBJgW2eQmp4tv
ypwOPs/gM2JzOoGh6Qc62jnFHayJsmEYAzdY/vA7v55ct845KrV+tvITB6VJRKbF
t1J7Qvkld66ipMizWd6fr475S/9pNqEeTJG4KLRPrAl1LmOySScrq/rEt335dCdA
uyj/Slg+KBqAPtG78vRwdCedWb2MH7QNjZiiA50vEY4uxEy/X3jKktG0TFHh+s+t
4OF720+/M5VvLSVU+inXEoZU0WX61/qdb9S+sWUQdG0KWUqMPzz6Crb8UVVbKonH
rMQIggtDpwhCYNDSwfyozvTIwwSIL21uSzwboYGdJ+ElgjFXYJpt8Em5ayNJzapf
Yi4MLGeftOWQPsM+lVTxiXsb5vhNn+Qluma6gCejSUWlTQ+FK45K0xoX8SSWazXT
9xLdVO9tXvFiLDUHUC7XP19awHv4zb9Ej0RjbxCo4XRserNm/s84/7RweUOPq4aS
sxNzQNiCh5wbQWA046Difq5ZBfDGLlSDRu2mib7kBtNbBML2/mJvCeDKVN6rLKuA
MIaYotU0d5jJUBwGTFUlgx5X5/AQj9WV1+9DuX1uN5HyLTW94UXwVBk5cp2STDoc
UOlvV8GX+41hVt8YCD0LsgLu+ac+EQMAS10qfi0024RyOU7Z8wka2Rf1NHjupiZT
ZSseiC9845us9KiDDNgneIDQHx68tTQm4Dp+Cf7eBn76Yw1PlWrB9926DenNc8qP
Ez7UYb2HuCLpl0UFesdIMuqpgx+3KJeWe3UOTNX6FOZa0xkIOJKtEaX0Wiz1UjX9
pauufKqNSIimWZHwwn6hm5bNPPlSyQVdCFEhN+xijhkrtdg2+SytwKA8nYf6PwdS
9JUpXqEHBPY6hMxXVBxVUD5Qb+GzQWWISCVivSuORNBS1l1R/t7C9DZvxpy9Jmbj
zClIHKCkFANv6Yp9T/oJzmtmbyLojoA3s1mxVR9Z+UBVM565hxCbE0jn+uJAwv7d
pM9+s418Z8NbFSDU0sYGEeta7RIQGjTel7SUeqb1/NwrCt5Oocfi3VXb8ONaZCOn
UI1PIhI6fl6UfNQ7uni6cApyHpvlYJdfbd1FuPfdoPATZLuibxtx19+2nd2//Lcn
tQXkByhse0SRRA6CX6sCamgJDoXXroFWCEgvON0frHlv2Uw6iPDI0rkkGNqDciDH
+8Yz80vWSQ5kbrxKU/JDzftiA9JIG2Llt0t6eRKkuvS2iQY0Cxc5Q2Aa4X5QFpqK
m8mPr8A0+kreOLhXdqVc/R3ThIGOzpe+jIe/AmYY8QB2uTKC4CTO53T23k063w6c
d18IeYVPoJQPzk2uFRhYbbFTGmTlrtmauq5sjU/NWOrQugckQoT8qM6MWnYK/9oF
heQUvLOHc7bbP3T8P6Wor5Wt2/+lWhYMZcz9BDZXMYj2UpC0k6HKQ+GJeWd6IVeI
SuxofrrWZPdhNXPUeu/MFxc0DD22AiNrh0hg/MbawN4fT4siU68JnwEMcbJyst9j
PR0bMDC9TiyIM2UoBz/M91EUbUNEaCX0l154z0hSgdSfLNqdoz9xC9Bof3EW/ICb
sb40xO621WiQBTyv4enkJnMclCbh3RUdssn1A9eNAlPaynNturou88WKhKxUH+Jd
fBfdLGisQ3DGY+hSw8vCOvq6l9bOya6zf7QKyZCb3gGdvKyAkujyL7G+oIQqZKH+
sb/BDne4D/dmH1rHiUiKOOkgN6h4f57ENgSWCcqtypOHHefmZ/xqQRHFI5nSEZIf
6kWZRo5jc1Uaedf/EwRVDrO4XsIRVpgLklepAth7U7KkY6TkLFQJiomikDmqKy90
uYDI2LeJTzrwjxc0meHHHn2K8f/YcM0tV7D/U+YYSXI/G/SK3GEqed4jVGLJIjqr
ekfOtx2tsZZYoXm/PMO/7uesCDDTbjvC6MmROWb9O1sCJtwCE9g+DNMZwu2nbOkZ
++u9L0s3FvcJG0RjPjJtDbHshwygbcFDr4XowfyjXIDcgZkmiOaqXWh4cuKwwPic
BcEcyx4TQqHT2LO7S+07GAza8iXUUkIpUjpOM7UqesxRjUbtKF4En/jheu8s8NYz
S/myXLlSR3Yorrcyo3/KebUrNZvupVo6bkk3DdJFq2pFHvLtO8jRO+lqXySVFknc
8JZS1Nl3hh7Uw2gsYVwPVdjHsCx0EsSfUxKWe4QanB9SbSP0/GO3cP5liqyhGSQt
G+qIXf8vn9tw1Ayzk2xYy5iSkXSIpK4FPbwUU6neS9bXK2mRPmOpzhyUVD4ttvC5
QcWXJLUCtydCQ95+A7cNcq+wFqCe+ACzsCYSbMwE3bx8Sav5dfLTWsPMJpOXkh8W
IrfZYAlV29jRIIxxs0+yFSahSbCRMR5Klz2SamB2jib8L5eU8ij0BQbeeKRf9S9M
ipu+I3Se636L9bZZzYR28BIDQUMLeOjkJScWd8JO+h4eA9YuiQzIiVmZ+G2IDH2y
E66rvXPew1yplmgEKwJPIchi/hGr5my6wo4RtWl0oiZYxhp9NE3djx3P0EWsKTGI
K/w03jqI6KzfZK5xMSa0ERkIk07ZkStviyt6VtRfTw2l/E4GWeYuieISznLOgfwR
y1+LJ3sbZnYuWIbBofK2BpQgcRGCHbaovEMx4HIdsr6iz5aL4ItRr0g+6YxWLVBw
dYiHHHdEp83Oz0axhGZPT/bHreSrXBfLS/FlnHUmX+kr3CSqKncprKzllQ0fJJMt
IXQLKtcfPYi8j0cZmuE7qQ5Sl9dZH0s0JiCnjT/O9l3DJ1X8dWb8FQ3OKGZNtbCl
bpJtm2nIemJrNHE1cQP9If/l1Sv/3PjwVmJgXu6autirWuxkDWbEzSBObauWHBmm
fH1BKIGkv+FMR54OhuVqk0O3aQBktrz6Kg58oZ1CB0eekEaYHPJw0mt0T/mLu4Wq
JvtWTtz0+pfjfpPXCUmTV/QIgHE0Gki820Gvmxi0IRNlA9DEUAG/1j83o+WRzfoR
TyAPN2WqJG26NbsdPj0raGx5rhfEEg+i8ajzn7MsZAo+ALupCUi6jsSZ+QdZxVrL
K2KwTr5UNmgX8T2mNBYszPhMAd1Cq2uonn6tOYpQNgIt8uxZBuZUHyPCw0215/vP
xbHcD70KxTL9zSZwLrOXJ2nbWZCP2/rBCGnn0UJF0MifkvHiRV3gY9H4RzGSX2c5
vpEmKMf0LRU+cZPx+iPRd8vMbNkHEWP8VG7p5YURxKyQwMnf9PM1Dt0W1wFaD9x2
yvmh3Mj68yXJ7Z5vUmfyBX5gGBAuB3IY9hP1UyIiPOsQfcKQqU1izLOv1BNKS+fa
LIJ0tP/RCdCuUU6pRv3KUcFvO7IcjXtuQq0NJe/9hnml27LTvyt6YRwKFM2W2rmh
WV2E4q0RxwGOek5ZJV6FU6mguCNA6d7vzX1pE++Tpdy/jNa1bSu527FufpeNpFSA
Bf4Gup4COMwZZlxvwjTZeY14NJ7MeiYxwBOU3dbG8mOsC98fMHJQSvIP1mxQN9b6
0cY7HO8/wiuTgxKBpSR2vUscDraaiDNjJvFEETeAo1LFcPxZ7nK9yQCbtapQkvwb
JZ4gIOSlhDeWmomZ5NI+/llhGEEF2isjnhWSZn13cnuCJU/THKjR4/E9rIWY+D3w
Hy/qRKbmaK8vhNcKKTZin6rUrT0iIW8yTpAsvyOINQ1CFrgSaEfSYl6UOjPksU0T
nOsFKk4Aqp7TGeNEUVD/g/32a5kGP42xvmD+iPNyn7RCFdoA7KAkzPfnsgEjrShV
0tE4gt9wPLCDfKBywiq1zR+tJzS9veIPyxDbubKBND0pPfo52Z7Io/sA9C2krXQp
FWocfM7sKYza9xeygLsjjnxU9IluYuegSe08suDYv0BzdATj7/kFj2NBfkBxAIlM
w2i5PC6DUL7FEnBNiQ58KO/3ZT39loIZoMvko2f4XuVucQvJtEqj+7+FJ81ViyoM
3glNhD2dwQp0lBrPo/3bHh5sFNDJACDwYu1Dt3w9yoNv9ZzJpW9xafwleOJNmsNb
YnG9KPZM5CpehAnS21pft3VdrHBQrCdNfMcPBsF6rlSKpdnH2teMVYRK8UXGCLey
TFNXKG+Rpu4tfhjt6T9FLURXjuCNDT+uxLJDEchRBnhektO+2VVGQ+YdV4S34Os4
YIr7rs1+8IKh4UeJ16KF4+dvZxgxdjdWFdRzqfAOI1aA75k095tbfkbQyvcaLUhc
W+p8KVnt79ehquhHK3VROq3GweLiDaHSE697EPygB8gCaKSa1AOzkzSCDp0KNRfI
GEk5Okaw1UdmEJpkWln6NSyQJHgBpvUTt7VgDGcjlY84E3QFJ5aQNssm3jBNWKyP
sp457yGv+6mURcig5VCV7EZvI3ZXG09YwUa4DODv1V2u2HxLDE6XCnpIhNXqzSgO
zQDDDzVukgdt15/2NfQpxjwnYGWgTGqckZ0N0OkM+CgO1D9yNzH7j6LXZFLUgfIG
kkbYQuJ5mF49T2KN18Y7+IZSuJlqlVBPFkUaj4puMG4CQZaYc/cJoCx3x28bqXEv
HKBaZoPOzsUcvrmgKVFT3QZzvy3FVjjKV7FDDLT4U9CAQoMINV+ZwUL0WsvzU9Mb
FpC/ohRxRW9c1IDhXkUc5UWsVI1NoK2PRZdrqNnb7Q7aLwPzNQ8v4fIaX7aiYOvN
0tpTWCMSTpXABilcijtnNe9awqVbx1LXmb6jPx9dGdO0YqRmfTydMwmcWGZAlnoq
A1kxyv4ZctM2wn+WtY2H5vET5BB8890SvEzD8t9qrZa5s7gwwd1dZhrJgeiOIwqQ
SgMHef7ElRhIuZqLxl0Z4OlAUViEcRbHOopRB0AI+OEHd5LavlbszqdDfNlgYkwb
HOAs2Yd2JrfmAagCRsmRXl2HrirvnqZtoVFQ/vh6JsSbhSAGnHdO+htmdGJAJAsv
wQ1ko4HiPZIGYLTokrQVA7zY8aWwZ4tCflh0EroT0olmYON9srKulhqEa8Lr2jSl
sWsoyZxNeYK5fx8Qdf9uDaMHkQ1qXdLPDmXUOrncpG7LJADRh5FWUnP/ADPXEmoK
ldJKKIByEtggTLJViwTZRxKkWEgvWOI3A1ruEKr8G0V9XxnMA7D/oQq3DVnZH/Or
ezu9iq6/lzbKtXBq4+wQ0bSRge3idR6A8f7hcfjKg6o/0ZqBclVRhH00yG30qvK4
AlBDixXm8w8JYBhfQVxDp5dmgtcHHZIpwrZLUb9hkQPjrOwq5nEb9g1ARxz2hyTP
hbe+SlBhQ+EkzcOid30cocLIGkYleWsRAq6k/dktPfJIs1s4Fb0/zC8Wgoh0sPm4
b40LnP5G8GNXMyiuh/CO1eL0y9b8d0yVkvWLm9BrPzTg4hp4Z1wmcJN4fvv+xxTG
Nb7V3clyQTYGDZTagISqVbY2InGmSLH9hctqXvRJRao2UQtqn+fnQU0V5qbH10Bp
SltiOl67+Ig9pKRm/Rw2sWi8CoSpxezghwGM85g9QN89gKnDPn0PBmYujqTRDg0A
CENcyP7Isc6P9xqKQVC9fktTMrMBrHF1XyDSymvFc8lybyBcUGGRcZdYSgFJkYGP
pEhT28eIujijy7TohWxiDC5XW816Rty1VDaKW5wnlFVH7iXsktfiJ+Yq+3Pze/GV
L1LTL7q/Rc+Bwdo/7YjftrP0ZFeqshrGBWnvwLMRGQmN5VlSFo/dzxek4JKKgNnB
QCy2UKZYDpnZppvoSDOur80KKFQRSHl9O5yvSxqZSn6EiaERkSWG/eI69tbhKY4I
lQx4hmYL6qAXi2dWTeunB4AqokF6U7ZPxFbWDC0uIplLKa1Hh/l6vPmAEtEOnlRt
oTJn1Y1Kf4DcPZttGLzTCEaHZ2bpQ/E8XU7ka9JmBfLOH+fhHtE1Sm+DhzgCAr/D
ZDceDBrxXsGu7ZPVxWq26kcSrEv1/TQnBHVrc4LXIKisdV4O/BDa4PsNohOeLNnY
nnyALXY8Igx3D3rS6R4b7ig/UgUCVx6uhNTdzfnxxgTxG9dcFJZarnSdbAUGVLbc
F6ErsAwD5mtSR5qGPT5+RQ5dLuXxHj1vJuqLvEH1CBgD/lSZ+Br50slUFpNseB9o
6kemVfVkQ5eD1nostT6kPNq7bRFkB6aC9344VWQZ8rog7YIZy4Mo3B3rGCBbWJa5
ANFCZkYPi90sZrWan+kFmCk0YWNX9N2iaBo56FOOxxcuLVvoat/gDzaGqnAcIbF5
NxPpf7guVJwq9z41s9/mh/lq9bs05tuQgUaAdnvE2rwfPNpHjVAQ9p/ITOJJvG3N
koBWJ5APwLIwtljd+uPr8GzP/FJblxqzZhqvo3mtwUf5ReWxK/rKTR3ZFSRXI9zk
5GZv8HTsGls16gFhPUo0zeYfmiNAk9VeX9jiazqjAELi6pL/3jGZuEi0nQvn+paq
fUtTf1jgMxM8RHmT1VdFMSzAV8HDqxlI7oyqLaZELeGFiamZJLg9p7Yp+n/2wpqt
K/xkpSQ6hdtClzdnlMbEGealrS7ruafmPkKGXguWnTSdm64JYoDKjMxfU9Kyo6+r
kGytsVbduVKLO1ogQBYVm9jxvbAvuA+Ic8WN85k21RfZZqX8fmM1L3NXr6IiBUBA
HZlkVQimKSR62B1kbXORN0ByQ3iNq3GhsBMUHGuPnHMAnvj6t7hl2KSEjbQzR7Hq
1+8ECqScG9RtpCgCsocxLk9y/naZCvt3uqoqr4WnzMGFCG4LEdSWxq+SkeNzLRnw
a7NhCDGqx8H8i3GCVvOTbfJPXBHCbhywIygb1s3kkuxlsstWaVHYY8FUslcJJO67
0GUyOKtZEwjjzqzhxrEL+A3hMfp8rl8/LW0bzbfmQr52xxysmCpQbD3tZsr2cqv3
1Si2SZKbYo7YL8/Y/r2S3I5iTkzWoWC1NyFPJ4J3Rxv42bqsrJt4sGYQdqTdCEM/
r1iHR4+/qxm2mQkL/bw1y6b8hb/wRXzFLGbMlxEWtEfJMgMPzt8/zH6NnRDi1rmr
P/WNtjc++xQBlDusEUZw6upuWz+yg59k/AhezvfjtWskKnfGOpBCsr2faZGqCzcs
GpSv+eU9q9Bps0AKJK46/e/yJwsG1CRrVjSjoRr2JE/cHwIGotvPRHgqstRc7KCk
BaqDNDq73wbXpN5dRIN/Ak7zq1/j/El3/d4lsKOk8fW65BKoWmOSk+de44GCx66r
jLfJYkQidVKAwB89KseV0APEryPo+vqYpd4vcQ9iJ1nyJniLd/O6zohk4jI3Ksbh
xnwU4eyXQiALqB3ST81sBguQB1ek6HlUg99xgGId35w3KRcXWRIPcaOULwOeao29
2v871C+T1Qf8yczmQh3s9FGmvwQr7kWkJhcksl2mtLxAy0WdvS6h2SApEY/B3MM+
GeTPP1MSFqxJf4aa4f+Xurg4cyHcmgV19W7BC8M2tDC7aopIAiFdjbxxxZ7Ai1/D
MMgGdqZQQbCbbeAr9Ej/iEXzSitXtZtdSTHRAGINzkVKBfEP4nCvEV+NgTCv7VnG
Srz973vliYHY5H1Hjp2C+ybSQDdyZJL1tsluyk0KJPDT35EktduZIr56GXAEwa4l
uU0gphyoWgVCWQe59+yh8VO9+4aiQ+MZH53BoPtX+DXaAsg/aIS1Nd7hK96n7S0Q
A7oE8uzt6PN5+DMoMMI5B/W/PajGundD8TZtxcv+YykE7GvgzJkW8ZX8ojVsCj9j
1k22ft/fuLFub+zQ7izo8hubeuIp/Q+HgcmuRuqraY9oWdL6XX4OkPgF5lHbFbyZ
vbCdTO3qxTrY/q7LF+LORJF0SreP2D6DYgULltJicwgzNVFoWoZ1dsWxrvrOATvS
IhiASLjFJS/pVkr8tyUqxf3cM5NsJuuO1HN7GIWPKch355MeelzUONxjfqIF4OU1
ONHRpAD32GEM77wb3CtXYLv06UNTegj6BbVdovTa89xeUsjsP9lOHAoBzFNC2xkK
VBpivnvABzKoLrQvf08Vn1nk9Wek9aup25powRb9u56EAUoq4Aj30+RMTxljSs6E
rXMyhDfj1xAweP4GegaxSn1H27V+MNyqxzkiZuxq10h57WhYqvcJHV59NtISnuO/
vl4dvcBuwgBlX5AIzpaC3+uP61Kt5/RaJrpUmVN9No8Vz+mp1pHbj/Yj1beY6XMs
ulgVOt/CkdFM5Naaxt3vOb7e3B780D36vMgTvKDLAvaxpNNQPuUWnmpITHcq1/la
QnMMriDDYDqsVkPsZfOX7guTcW+8u6kryY2hrzHlJR3u31NSu5yL6mXW6Xq+tCK3
Z0X9Mkj2Y1lpU4LymWiStWHLJdN8tz034p8y3jy/u8q/ypYST6Tg7f55E8oqOdkJ
v4uqf0SBcNcZ7GEVSplZvIMK98Ho2cKEcY+C9xJMa3G6Ltl3sln1RnE7buJfGS6t
fXtveiAiPf8eMxlQ45Mm0GHhDNY1ZJpqCfMI5JJupthnuM/7P/U2kaYLc6r9+eRR
55WXpa8YOJJO16xqzLDwcXMPEH3xHFZFmN06Ui8CSDHL5CHebqDuCUhYN9f2FiUT
9pqsi4eY7ykC0sgeON8Jso4AdYm14zeIDMKaKDxY2+boEa1XZdZ0lAiF49QuKpOY
mz1HKRY01uIc+C5p8jOA/8XOdNSq98Y5UOd8xj8eVjSOLtwVzMjbe9CslUHsPqE6
PSQijm8/bSMuWqCH+OJTKVcMaS392hZcLw/XvVSUIjlb3QRpXW1ovV8ufrNgrUZs
GTyJCKGrpBsFm1ZGj4h3Tk1c63ls2cLk3Y4BWSjW7E/OSuI79rH9i0eme/pZdYl7
nVWrr9hrw1RiasKfxVURoxRFrAtQheeUbXEae99sDDZGs0mvQc9pwUmIezmDeGnZ
wGFBnsQmhM15uSlMxVO7flZK4lv+ytXr7nz78/9wbM8AKG/8md4Jh9yterPG7CzR
YcR4W0zxcYT6/nIjF0ocZa8L2wegA6myr83dxbldocXzm7vn3Rry/D4VRyzK67sx
bKdUZ/cIhj55v5CQzbWLqH8uUZpy16iUah5DnC3LEy8wEHkj5VT8F0iQT9BSRrCu
TzWG9YYb9koL803yyGagozZ/WqFgF8i9rgwzvxs5sysPnv1k9BireH3d2QwgAcRn
FSaNyQjTZEt1Q3YYw8m/et2WWyXU9yeCx5hwJis/G9Iw7SmV9Ir9Jyg7tZpTVTfa
Kv+4tH9t2Xmx+F3PD5d7AfjUyR+rVn4YGXS0conf98FS6zIUTD+h0qt3D+c+vEqz
6C0AqW7mN1V9UJoDKTjXcbYQHMtIm2WtZ5h3EUV320libyhwjBRYdGN5C/EBBe0n
gVceb1gAQu4QkgN772g8iXQaf7dXjUfLpcE3UtHVXd/XZS6tbcQd62FpqLqxR56j
W5ZhmX66Bpajv1O3Ax3R+pIy1lEStArVSxMXnmGZyv652g7l8w2ShuVplnFW+/rZ
IFK8M4VanWnMEpd2hYzVKA54ZHme+nQUVmn0BLc5K47KnFz1zMQgdFAKCBWnOKp1
r+xNwKsaHYKzjVuaekxbpUIQ2/Wb+9/Z64lyUXYsrNqkkOStjvg9rX/JJwpJelO3
4QM6HPUO9NL+QW3psp4vIoSh2zHLz+9aF3gz35kfDxKoLulGO4uc6T6nu5WuAMfK
t6N0jKJdtx3w0+z6n3zwdNElSCmGAaOJL1gi60mTwtIFobC7z3h9uv0aWiuryiL3
Lul4EtGxIKklDNkUeN8n40csfOTbmFKZH8acilLvMyrRS+kmfg3wF4dBX0z3CAwp
WqUv81EdtIJsAHu6WVegazkv4NjRO3cIJzPgV/raTPitd+AV3sMUQOkMnLdsjq3Z
e0zOeLvRdY4aQjddVeRzlTdYPniwgx9uyOr64eFDLkEsgZNC7W8gBEZQBvzMaYmm
8N5ej9prI4iOHQ8sUzFKlGKVWWE0mexsLR16X/UaN+Y5HWqu1CKeCD9ryArUDnyE
+ahuW3TT1dFjuy4t3JrThLuI8189a7UoDEWKakMDpNGae8+wARI3aXjk5G1GHLTC
T42rdmoUkoFd2EIk+84ZsrGLuQg7d0V76oJ7ZFgFw5s1W2NDXXEUYU6Xl75R92hu
TFdjBk6WFwOWt3yG77Mh3MFvRMWmZ0OUNfl1y04hpyoW+WHmISL/WIc7jetx+A5e
QVGhYl0EPelJQe0UE9Ou7Fw7THmmQ4tNEgyE3PsPWzyVUbG/qYk29JU/VjIgiF1+
nO88zoQm1sEnWgTMydp989HHtGGcMKsf+hjSCUWt+0B2/gjSbjuQpqN9wlupuJTZ
wx8DRwgeTlhheNZyqKUClH2Nw2DTHWWT2TpOuq5d4oAlvGMpjIvZICwB1iHox/Uj
4tfOI6w1H9rYF9barIDVdKNxW4ZfN09v/S6pZGSY9gHXOWIb6xeDaCF6tC4HW1sK
nGOpbz0I/iW63jpKEB1v+avRcuwJFr8iwfu27KMlZkM5G1bfS749ze/uQyXi/SNl
epUz8HNxPLl0hgxPc5/p/1TdzgPF8V/hDqz+Xaj3v85gZWecmqYQ6ONZgHq7X13Q
9pXjBlYKvPGDA/DSiJubxrC+yXd+wFeCGClUSmmbfSk1biTz9+Q+8ZSLdeUXFmEZ
f43PuKlZDx/MfAUkb53FSaQA37x1zEE8kqVdZW1uKZBeX+gyclzhioBROcaRGj68
QcbQ9oQHCMP+uRB1QP+7bTJHvFpDowzwjzVEjC6g8exm8dayq8j2U/hF3udwalry
jpwLhxiW/cIfGOhjNu/TeBvFxmR0G+/w1DGjyPn0iPWLKEOYdDkJAmxV7HqldEVq
XY4gzs/K0yMBOgxOksJBf+rGIFwhU5pTEXLwSrmKip+TKWytHtZRsQXzChmyt3Gr
8rjVPQEirMouL8JGw+unOak58lXTvfbHkE4LNPuPZenK5OpqZkSsg8DtDqncFNfK
+gcjdNpXpb5ndsjeLisKcU30d1MlryJmur4rqf/M2sVYIC98g2zbSxOxFagLTbZL
7w6FOsaoWzjh1lZjTWR6AA8TFr4OUYi5s1XuK0Om9Fg8+0OlExWM3SzZvyvGPGEQ
ApZndztR78HXjOoPNJ0TsxUbqTYLzGAme5DpYscPr5esDsF7E77D9+UIivbAgl+i
rHLRLPV2f7aJ2qC5J3bNzJQ/7MqUwIWyZ+pgpJI+JgucwkQIdAxr4VtduX4Mpr7n
8ba3969iMe9KYFXmAZvRYkr5ifKE412C79pzBWPFg5bsg/ODoGYRU8kvDR02IuZw
bjWNvC7Hle+L8GlfVOE8ePMDyiKQpVgsEkzadazRgbJ4rgGBXRatcX//BxLAjk5C
VjP2wLqQlhYlemSb6z2EWmzIHQfmrTk2AoJ9HZlEVgxzpupxveXY6niw5v1Bp1wc
8m/oOEeBzvrZtvPX0Tc9pEwUCgmCdJfjPHyotR8KO7/b7wmQpCOQev33UKfHibYg
6tqMsqmm7YEHuR1Vx8ZqBlr3yKB5mDznBdwiP5pmLEMgQQfVPDvR1RYvXWAg3gmN
LMDli8LBUAdp7zzz3+OTnH1VHjfKxl673HeC0nsYTJpjgCrmF5w0fNvTOfEQGV6M
zl97U2Z4hmXtN44mH1OI+5lPvk2hjSjRISJSCL8XHcKw3hiNKcI9EyExM2SuOlWT
WcgqYkYlVAbvcR4nGKxYXiQ7c/XPVe31YnPrWepa3UIb/skjwAPeceyH5mFKWrvQ
B3+Efyya92pfSk/3d6TpCSzJSeg9s4L8H2GkgGKjVjvOHUfplajVyUSk5YMzgvCs
LmaplXdGoa9R683kj36E0mB8tLIl6+l+7bJA7l3yeruM6eipauK/iXvhqzGp1hdq
o5MBz/zkLP+5K32dyfJoLV8lfGrqfFvv8LwQ7nCJwO9QGmaf1aWiqc6sx97r6hAF
kFCSdQ5wHYHImAdSmYEJlgNZjPkv1QjbK+gSOru5KAOfw2r3PitMVuzpHS9/ZctE
HQhinCAKnebT67mfhTflDF6oPOzV/HdXGTNK95gQD0M8FwIDDDcV/PavLPCrfJPb
DVV2O2bAVOVaaW3OCOCIolELJosEqJ5A3EYUSxENepZgrh2JbLXDm/FLKdVz45q1
rW2S7EpvR5vN4YndfSUScwicfppn4o2i9fv1O77srw6+gwFZNgo1EoZw97P5JKX1
9hx3mC7Bz0orv/5kL5HYOIg2TUU2epKXq/wNwEtaud2K3agBB3JI8ltccT/y/11O
Bqipiu86B0c2W1tLR8T+KCTX/s9TWG6Lv7U/1/obrL4JKGwHxe/+ghlSSci1LpFr
U/WTJSBo1UjR6EK3HKLXwjMmp4BSaycB4IrCL/i+zzkImtuEDQxndE5bJ1Xp6U6n
7R2wgzdrXKLFspfSI+NQIDIB3nCjIOP2thcWehr4wMUrNFWYJK/qfMBpJ+IbvLHS
aa+p+2txu7I4C9el8iTdORLl8bytppfqXQlHxPhAyrnt+Qa7EMVZEmRktnfiMmDB
qzqb7A6Sd3O03iJswXRfdoAKo1e+mHvWQbOaR8YtnaHxWYs5DhJuBP96O3v8TCQ3
TpQeLC5YeumfkneWilYToj8D41Qr8fLNEHQ34Da5jjIHBpVr2XkZUavZOyKhy8kT
Xhnur4nScHPdS53mUfq8texegelxogm2++tENRJ/NXg3r8R24FLNhM8vU0tJE9f6
Zl0Lzyl4b27ozu52JUgz6d7CyYSyMDz6EtIGE9VyXkhU32nIT6PRwkwp3FzLymjj
y7pHpuuFviqEWpe1yrY2W5kEPfCWiLrrBZT94fQEwNRi7PWVOfciU7R0w117imvg
o7B9O0i/KejsGvJgNMdyA8hYVKd7Ky+kZbX5zWfM5H+YnHI/LaLtmkhgE5gvEvoU
KCfzRRJ1BQwxN9nqzyzazVZ6z8jgcBdlpbt+ZCjMSwCo+S2ngTa2AMIdZ+RfWFTY
Ffekfn1NT4IjdJYFSwsyo/taUq7z1exTN0rj1efa2MZG7sYlGeBO3h6E2C9H68hm
VODgCuPNgbwVx6qUpIgN1yJReHFHmtdLEIF2I25F2LHIXHW2Jjp30aOduJSNRquL
UerPyVeNVoaCjWeNHZB73QpQr7C3S1eLhCCGe0f53uLr+wFaXhtP2n/oTRNqHD0o
+BhNj1EmQnD0Z0UaRLeVM8sxB2v/OpTBy6x24YOctACTDb08k4ZydWuamb1QnXA8
i3rMyesB/n0GqSQ3dytleCVwOOqoAlPfR6zh/0ITzZaooUBafQnJmktp5TLkzkg7
vrVu8FwFS1mhHPmDsXvPIL+WbWbHVis4pj88tVpJzj0o55rIHerPY0qrgXItlzV7
EfL7lSbiSkNS/ePyHksJ2tVHR7ugYsB66K92YY6JghjrzTGSYngy8GteJT60/xlw
Mj3iAe5I6GNEjoA99Qtoj33V8jAI3qXm+NuUTi3cDucDBdSbZGoFaL7yq0MWmCnT
llL7DMh8zKJntLPxm8kHspeuF8sHFBqbtfTmPCNqhd5U3UCtbIQ0B1V7IZLEUUoz
GWkrPwbQEXGpP9zVNEXgqxUlDqekNDDU1zX7IaejsnM2fodonRSCdr8Oq1AO3zXN
T2JE8p8jZ+75Bhs0m4xjryM6K1lhYgQRADD7ZymoRFrUsfoluWhdTWyVGiru1KlI
E/Z4a2CEhAbn2e+0fRlqDR3ZWTSJHHx4pSYZyxZoCVBJcTv2+spUPssD3uXLQGbj
E54QMrX/iewIVHg03IBh9dwEbEATCfY31OGgY26fYthcx8mq9MvqFhyYFQO5G7c0
2Quckyqt2AyLK3HAnqsLMvXyhyolTFd5xYkYU3ZoHryV3GjiVRdrTI6SrV9enqPG
kj89H3sxHzLWhWO5kh9Sz09nHS/XrVj6S0ptayQ0TsTiQ1ZV7yArlhAHwFIA5TBW
iayYXFpQgY7AdBTUZkVNXAzjwjUEN54DPyUYXjNJLJajSlejWrs0IDCaJ66/iB68
FJlqNj0/Gb32jhwRRlq2XmVASBN0h5Uwx5pd0/TuunrtQ0CpdWvZRM+22lyCJ5YZ
S3tqLaQpylSCI08hN+Rjmbr/UF5SVU1N3PSACtOEBkg7cyXc8tqmrBAnwop5XPVH
Ioo+4go/gyewZe1znsfJdJqpEzowHpp5KJpiRGv/JmjDw4hL1QRMJyDEXoS2W2tC
N6U4pvXQHDNDkbIrKoCQ9nt6cGd0aI2UJhFJ6PEtjLM195ZnpdxEBPC/SUrHBS2x
tUNArTfjQSwZNKxYBsohOUkkZaaZbezak5EWqcrXC8cbDul8S+qT6YNfuJW0Vzvq
BBaqLiS4EAtzQwV0x4YuXVCo/MYrb6rZZS6rFqHi9inK5YKonQy/evkwADKnQFqW
aJurIgcu+hPjObW5rBo/28NqV1YOYvz4S1OwGDByN9UA9auND0ZuwqjSTaT3Rzaq
NNg8ALpUTxWa4cuUCuw+IbCLInY4pxcWri3Jb4LkWL/smlnuluiw0NNfvMh3rArN
kiERuHJpRiypgntZ/VJY1tUBEdaiuVQxcllfj7gY6mBamfkhiDH5y+mJkByLJxA4
E7yEsELXJrcuYn+5Up0JzmJAW7mYZsCgC2HFd15cKoq3gOL28UgrS3mtH1RsVdP4
JZG0nZoxc4i01Y2gXzg7M3fZgxW5gyfeXc8jnSx9oCK5U1BEijAZy3uXz/NFi/GF
1YXyinqoRSsqeTx2lkUSyAbnsWJyQh8yUL1RALDzXhYlJ3LlcWBRPkEL9/49OEaA
VJT3TxvpnfST37Pllz9nlN1EdkdEksqsksnSEJ2g9g1rjaZdykFOTYX9STHiMCpX
vEn8+3KNfo4oIR4IBVq10BAJsVQfvR4TSPA2KhFX46hgtMQANR/dgfYARN/QO4gN
e5J72602cOdr3jjm2B2e8zLWObsWglcGeY0P5npbXMDGsdObVdBo196we8LKrjYy
xQYKZaEmrWj17MtW8azDRXWOWRH79OrKfcN77l/NwSGod8Jh0ygjldPuzxzmISwa
XhWuSynF4Vp2Jf5+PBE1ziiUGU5ECyMYq9iKNMbNt4rsDXHWXWGkln4NCS/tChRa
2ABd7SVvp6N62XpUWxZc0ihA7oi1cCM07DXnvyYDrrk6115m9sBH5hcB1LwJuTiM
BEf6qZozSylLK3eH/sDstc2kRXwCIs51uD/XzzHQVUwcFDMXXlMchyYc1H122yWR
MAj6Pw8VobylPb/0dFJtFRpsruDY2BadP16bhBt/wxpNIEoms2WT0uGbvWyUocKG
HfB9w5r6qAIfkhe4yfIhMKxbr1Qt9Td9jAPwVSB0KZdvupqJo8T/yo3xfxz01ahM
Zq+Qe58n0QBN62ojlJAxfQWwdqD+1Yphbcb9nj30wdHn1y6hwyF5fMpQsao5J2zp
qoNt3EHXmbIPYFA3TgMhOfYE4A16UInmgCTJHB35T2kVcPOC3LMr1iYJsqKqK/6v
K35oYO7HuGYCqVfk/msR444nBSZ8uoMg5AHc0tvapxyWjyUfZeYEDeopnL+E/T24
Cl3roHRvZshnpHULbj5HitY6o/9Ys6r2TGLh5KvB+vFH69o2lR5B+CTI1XgWZLuv
xSlIGxSPIsv8WEVMsgVVqf57XD7SA0mxmEUKBwujxP1XYYBGm0mOWNF1KfCRtb9V
ujQayTtKstXP9R8QLmyZTq13OneSSyyXHc4OiLtoH3XgCDy6PDL6gUr9G0SCKWtK
hKS+cmNxN7vlfCfwE0j1OFgnmpQ6xgzaIFRNxaUYT2CRoO0OfiR4U5lVAAvB51ii
ldwDTFKpa15oaTmeq80PKZeMyqgn03pU88GGrZPgq7J1j4otqCry50uYHHElZbKE
V/tmIt5opIUSNGA6jjKCnxzdu6NhmxJvZGiGYK+/WvrmI8fWKWkqZ3okz8PpkpMC
9az4Pd0cAogQfZgFMbw6UC2UmxrHu7yhBpUuJhFRY6XGbBrEjh2A/e+6WWQOFEJY
1SAx3eVMpYDXu6L2BohkU132UfUFvG5+Isx6jyca5tZT3Yxjb8Ax93hJ+UW0A99I
edOazBuQpowrCs4tLeRcKWxYyBeDVnKTnkVr54wqo63GqRJh4XFEBvXpfjXrgPGb
Cr+vcx7vRYhtHZgFW2TfLp6l7BT7TWpWYR2KgfLn2SkjNrB9DHjUmM5XzO5D6i1H
sz30EtXGR5a1cbm1nmoWKs50OW83L+LsVbVUY77ZsXWbSHoix+xxinvzuZcJzfki
s5FPiuYgkNV1hKGQL2CU1qQgrBnYNmZWphbh8nepMiPn6WADK3V/eLsvhP8h4GKZ
EzOS7cRVDEc+uFU7/55VJ3O6Z2eGTj1aGzJ+wBgu0YwGtXsAcf+MX/Lc+LFVEBNT
CirqQFUh/NNBaCUruQcZE4XqluqWGl/Ptkt/8GIHcrWWXdBZ7eT38/hKjXmTCfWy
XXGq1E9Z/CD3fSHFZcLsDj4FIkJlwiglhE3+HyyA+Qwa33YsbgW9NUfcE87IuS+3
BkOeFW1WvqKiNEKYkWnfw5N4jJJHdm/3qN/4N+rnfHXT8pgh75iRLUDYh9LX5ZE+
Vwa71K5jRO5q9EGLHZvMhKvOSscmpnd+cOn/1fUuRJ35edtSgoweNTlYQLA4p7+J
wqe8lWrA5aMS1IIyD7pMxkNRs5cBN0X1F+Ym+hlqRUyepudTEoYaHOuME46zfMqx
8Gr3ArC8INSEbA84TwyP/B18xOX8u3CqYTUc2QVUEszACoxigPzX1rk//ZZtqoHP
hZiEqDD3X+fZvgKXiFYz1XMMRbXnljf6TU+hSrl9tD7T8hezRBa/kKpJ9YW7obFs
1ljYailIvGb+6lGTgVOf0nmHDR/tS40w4UzA40U99lG+04kZIBfzRpehRGgWOr+1
R1t8ixik0m+LLWsX9yf8bTU56dcR9Qo1QwkTYGyKLVUHDgdVxdVqko1vV2Ks4xKU
xG0BFSGLhoCXdqw0hL/KIQqyY60aTBjLw3aI7q20PU9kkTKNk0sF7OMwCi/Np+pG
7F8JYfrpicKhEx9ULRXzuTl3X2+st6+nr/SWW95vHYR3R3oGWS7WsZ5f0cCnkdME
iyiKNM8sC6iCm6/2vGAWRjrly2cpcnycDAM2Sp2nEbBe29w5pg0ZUxwAnLUaFbzT
Zk+SA3a9eN0gQgecX2lesG1AiJ8tzHTNedNusiCm2JXuuB0WQYGYaZBP7xFi7Csd
ujoGBpdA9Od9wcjgxOnYxSHIGpCFxRWkGPbScjesOa7kJ5OseUkqCqekhwxBv8Bs
pxEB/CnlOeHzbtFZDZLfCCbA5A1EENCbPoVwJFAJCH54rOfgbdWB0M/kUgRL9IXP
89rEl6zUcZAfCLNjcjJ+an9Tw1+Qn+6Yy1hfDYRYmm+HPk/kqhr7zWMbREIT9ZyB
/veBIVpnuQUKY69AoEwzdiDPG6R2tchT5+Ty8QDvDCho+GQOiBa7NZaV7yUdBvpm
px/eyJil/+XGlepIIJ94SOtYonf3S1B157kaFDJSumsP14YvWcE8OGBiRC7VxAKL
F8bUnvIOZngx/q/XvXAki8TsQrjCHu6Qjf3zB9lJzPkK5EopwDApaOdIGuYEsUHy
CEYZybC1TvbuAEMibbV5C0GocNjm8ALlX+XDezHejxBLFVVLJD/Nu4blJzlCsEE+
cTKcqLGNeh/xCCoU4teY8ifMaZPjwtNrlKRLQVEGqhPOPAYTMkKNE/8oxw0smflR
Jwmjq8yvFaRAsajZbOOa70UkotMfGp4eKn9Kueuey6VVU350utmZYIPruv5JijvP
hcYxQ5Kd1taLf5v76Mq7tpRUyVriNTw9HCcwm0NikITu1Ho69tQ18RP/XuvyGLvM
9xQCGeUkYL7r8Pkrjlz1vl/EiDBGZwyulZcRwhoZCn8z4gg6oc7Tc+9qcUmcPerE
NL1JDtMT7b8X3a+fwnrrGLoBRQrSIyKlvowjgWEqEFby430tu5ZkP8dZY3PaBRTF
kkY4pMT5v5cPvmoxsRjOzCid/Mnhlhw4gJqI9vD99N/D70828TREIy1N46mOQSqI
77MdWAWJE1M4ff+Wwpj38zl+ZmPk2NVa9S0aDKEnRB/fPxPIs/oH4mRGLZnkdUoe
3EhvXX1w92/sw9+5lgVHa9hA3pRRP4ZruhMy+/ck9xQlm/5Yyjs0BaCY5qpYD0qX
n/m+Q6MQtOb2dnkXcfzXqTmMuygvvj/IChaxa4sqmp9BYJ7jo0IiFWTqCQQJrZMe
2D73bdKK6lsHS+UP+kzxuYMU7zxopEs7/lOMWYlfaRM8SVwllDTUjZuSV452ljyD
O/MVEFNyMD9zxAEpAaAQHfM6yO3uKRVluvbTiWfIffiUOgeypuQ9rNmo0na6Fl1+
eWrt+BkPyUDSVcsfW3XCNIsOtuoqMLdpoJhuODrKwA6EYfcupZNyRsBZjaVNeLiw
O1qlUv5j5f5n+b5zVE9uAjrAgKh050ZHUBXR17CGHWwJaYDyXebD6beA37HHlKZn
m/kRhSNAQ7FGAEizDGb4FnyBZFm/q070ZEti19f2zfEFAAqEelL2m5Qnt3v5PATC
OBKUSJDa1chQgOLBz0xPiBt9gmM/yb4sQxaeyrTPxDJKiuB+B/722hj+p4buvB2o
Q0h3a38pG2KBhGxiXTRQ/VTJZ2XQWJF/z8U3J0AtIrrS68dFXdlBpUDZf+r4NV9d
XJWbgmFE1zMrpyDbuH7N89KDc4R95AlU0FIAqBrbcV63E2ai936Zj+ScaCLb1uEn
GE3mbx4DIomCetXP8ImNQ5YCdc+ZuPISIG7B7HviqPGc5UuzbRqaP+HE2zJTXDmp
3cx/eaugqNAab+xMGBohFzNlcswlS8ZAaWEiq8QWwnHKObsTOeijYPLW4W1CTkMZ
VVnNFq/YGJbmGQxQjJokh5izAYKm3UHGT52GBk3Roup+cQ3e/GS76+l4rB9i2L/3
0qcwk6iO0WCGDNJgQqjcbF8HAIg7KXy8VuOAMvssp6hk8psYQ+iBk6I9kNoUxRSG
wulG93AhVrwDOq5YO3cr2pirsfRY4LGc6tM+tcP3rAIhv44MedNsd88AA2lZAr/8
RhparEgZUQdzjqMOGhImJ/2uyzmgXqEg+VVDqhrEkKGPRUlBoKj10JeKI8B3XWVb
yiqHwiM8MM0TwWNnCUy1CfFrgJJkG1TLTUetxBT/To03Z1SDKKB6TK9n+BqA9pbJ
UgWlqqxKvFhy0/IUfqy54Rz42CFckg9mXNstEEBouukoIVGD+sidRHY6qRVY4pt0
k2qA1U/sAiGGUxvvUO9xn5OaB7rONSnRyD3dF2gHu4f7vOwxJLydeAJL6iFjrtge
XDs7hxUvanOAOl2XeGBs9w3fCzfl2sB/uiYK9v2zG2hb/37/58UEQjjI88XLcAuw
FyKefMiR47DlzzAO0StTnKyG3cb68MHawy9b3f0RSmj3PH/FQW0WsUYsETicBsm3
KXGmhZV40PIfIGWkRiEckcNlDcnkevP4TEKcuGc/5fbonxWxBJka27kdYc3z9LeI
8AK7M9CFiWowxbh0sYlnEK7/+HHgF/6NL092v7vpV6CrBw/goykKj/zHxmKcHNlW
4N6FgLn9BQoj7wbHBsx+kO0RzHO/PMPb3RqydKyyQB5I32P9ZaQXYLUAsDU61ibS
OfCEpnZsElmEwuBk76TLHtmqmDIKGlKPzHefjNOXjzUapd23nKdLnMO5Yu6Nnxpj
dgqE/sdDw5bdGspnEMJJxr9TJIXnfrwEm9j+D66plXnB2zMsSwH/AmUUpNgd3CRR
3rBYbRPERg7HqGazueDRLQn1CX5tQBG64Dr6Ix0yNDPkjkunSbhmrIfnki35DMP6
S1mWROwVOBWuUetMMpLQoKs1PfA7eUGQ5Huzp+XyVoUVkUO5vymc3s3JGVlKLxBx
jU4ZHeOjHOBLQfovm02NrIHK8oGMJYxq8e0l/PXmVaUgX7dIb3Bb2SspqgLYtTS2
Ou49OkGWTT+KvXJEkkEYNNNYnpabR7FofK/eRH9Yeo7YBn1CcueDFPGe1/vqAM+3
qozjKuN9jLMp3oKp1/dGFCggkmofp3ZKBozrG9yers2HfEuSAyxspxSyL8sMIlb+
zytZC+7AqK5yIV8WNEu+q57W7VoOMof3IfYIdDnAGOmzoLl3imTq159mHpzwk98j
SQ540z/oLeCfVOOkJoR8MNu70YGUCKcpUaKorQv9zu3RozFImB09LARNas9jHry2
WmC8LmBPdP/qliohYHrKMg2p5Zxa2lLr38GOc8tSxQMbaY91ygihh9wbA9yUhy22
2O5h3J/pQSjmEgk6MVm3i1nSOR6KygoyQR9WMqnLVcT0/7CNSIDvxU4MurH8m/Cx
HTbylz3fTLt5bh9Ye85fh+CUvvgBxi45S8VqoXSUCMpFWjNSATC/64cyQBJ8oZMF
aopM+o5RINr22/a0Ots8HYLn88yqzcIIO2j2LARcgF1bCFCGkzV2yh7JSKbqKbXN
FZizXP9OE5fXFJuBqp8yjY4c4q1a533rW/Wi/KsuPIERZphyn6PoqBO5FJug8H1/
8kZC2YB1nrzEWfn8LX0ZumPTYfQUNECk1e1GG4TwJ4WlGw0ZM2mUWsVirfhQS1ax
/Ny98R7lcOQ5N5p7rtHlYwMR2SPN54Ekyek8/LiPjRd+OkT/vytK/7dl3bcU9JDh
U5YfaeZSl00VSDrU+AQVHCrFQ8NEVhoazbRJ7I7j5QGj2VbhRQl2Xe75BF8yD929
xogO5865PjyFKdM5vyFBv2i7YhlMRBpNkRNOni4YeLsszxdMtkELWs5t0dqt7axZ
WUFpxmLbWnzgZ56w4bgceqRda6aGkqxc54dpWXe+W+0ggs7PBknc84ixFIKC+n/5
8FKtK7uJheB0oO0qEYhZqVTUOcgdPlsQBl+RFEv/dv7JLvHMVr7ZSa3M9oCN7rrK
cWJjj2t8b4Hdr1VF0Y/LXinCkqIDbiReBhAOgB/HfCQbskBI4XfpR6yMyDk6ml9g
NB13/28p3QNdrX023H4kjttl7nv7bNV3IBgQT0qiwJi4FtWcoQi3wQ3dKtti5nzl
dV4yvo8R94hljk+XmsCWl7npidVz+Mel9/ub5MjKb9vbKJSqz1b290e6NhJeLacC
g2Cmw20tZ8HAA8zs3Umivn260gFQ03/tjB+Poi0BfhV55Z8LExrRFf/9mioXjx14
Jcl5raV5ayKcijhtiAKlXqx8FSNL3wiyhpihc1VIYjutP6YBNObgvUfvu41aNURM
c1j6jrUbknd175hW5TWhhACUkf64KRbSiezDMw8J6RTzH69BEC1HTffFKMC1UY72
dgdcQkMzEkEwaV2QYqGBEBhFJZBd2LLKN+Q7xpaBmFvCJdutXlOFZL8NM/OYIeZh
wkKA2Dg7thqw67O1TiZ1oYaILlf9ZSM4IVWNTDqQHLBzbNFlTmPJQE7Luyn+X3m7
UdEoMPNkpWyNIqXy0KIUpr+U3hMjaKbVQIVNvpkBHjinWCVL7wrZ2bnKqhhEFrZ/
O2JzO7Xl1skut/VT50PktPUgaefSiuomnl2tqcOoGxUd9lwNSzwfwiyslalvXSgA
0onRJooia6rvBPNAbykYzy2LWnys2nGB976axomNeqxkNKTxm7ZGA2UKIysHjwLV
VutwqLnbVdHEr9w+x4KXDeq9yDRaNAale7IvhuahXv23vexq3FSGLtH9tMTDPmzf
01EGv68h6BnZQWKwrHRS4w9YyKQLhHQ9rqC9wVZSkhFoOUjJAlgyITLBBY5qWTX+
BldnyhhcJ+tjBGKUpjsm10sqfNnNOGZ0DU2heaDXbvgRMmdNKAnu4VkWBg03839O
MpUvmtF4cowEaauraBcaXuM/t8O2a8ZxbYTKTm8hO2Pii/hMA7jz0DQASx/8sjsI
PG+3j6ShC2yb8rVagD9JW277Gap1QJYOKyV8xitNVMvQcNX7ueQTVqOpcU639kU5
gH1jS27khW7jGPV/6uDN8Ejtuh13TTxkYHP2MfJgIt5idEpghnZqm9iBMv+nLSao
CWBK8Sxqbv0mGejXS3h/GU2rNRFvebjIi9hTaEUxgr/0tpLn3QAGxvdoU+PO1+jc
5S6yQ+P7qcLcg8+iMBzxEsVBaxfYRkH20WsvAd6vzzunWyd4KGOhl175BaEiJaEQ
bP+lfYShAWZcECoXTr5NP2oZIQhC7B97ZqP3N0AywmW5KxoQNh4WuPKftFTtu3at
YBBbU0mqWCjkvQJd5sqNFIeD5AOvclVbq/HbaG9tBM6ONj2XA2beoU0RF2OLhTKO
sgWHKaBTVh8jiAl/ojmi6szaMMYSw3lnaTP8MqdGBwAOOAiZYZnBkckdXLzGzmAi
WGLjj1BbmrpR6Wv9bO+g7kISrdxJ/1gMIB+Vyp1emcIQwk5cvamOtNUi04dVjfUe
eYEY86OEaz1CSGMnaISHah/6kgFOyuS2tUHllHfH88asAD8spDtkAX0zkuF2BWp9
jFlyYL1MgY6+hP7H6UnFiG7/at8G1pYOoYAeRWyw9QJcMx2pXVON4iQP3fwDahGS
rSEk55cfHnLnu7RoS0hNS0uSyfQSA2mSaH/JNCM6GZIHyBNo8+/rAdArSVyLveVf
0IJHMI3sp5rjmrJ7foSCeEJp7JdwxlnTMBCW7E4DKogqpPoqkfx/NVhjRkDzZ87u
d9POkpeXw5vyONncWgeZi6NhXeew6uqPrwLtdg8AJ/IBGq5eO8iE3fT9SvUBsoLR
BmtI9TkJBg3IZ9PlC4YXgku+AJZeEPHIWjiproziwsrKoBTfHSYfr0vACRRPl2Wt
NZuY75q2hFLeEAg4qL15hmLk9eoLwJyoTn5DgV/Rg1D1g9JE4JxcLxR//CyG5rJf
y0kJh7NeMZCQ0D6YIOKOuY+oOP6/cic4TK0mk/aSWyM7jqcHzXqB6ipedTvUZcjM
FSWB8fthImI8EWXkmsHQLdTCIrZFHuxBhSpWwthxGWjRMnXuTvTEm/ZPUAP4q0f9
GtOeobkD1Sj9ugo/2loqfjVEF/WL6m9YAOwzii5Vp3qU/r4QWbDF3M64SHCfzeCt
qa8fkjU9/g2zp/A4QwhyfZcc8+hE/bSKNiSu9j27X9e1t7rTkizVXCBaMWh4jnqm
EXu6es71ouzXaBsSzYPC46KgJG68IGTTFlWOiHTnZ0xEZoVOQMoEASS0mOxMXiQs
O576/G8S/iak9UlDAYRR95vwyZ31J4lpyd20croQ0qeT5eQX9g8oeFQGieYbHW9D
5vYiH3mjrLk5j3R70xYBWr8zmfDIKq40bbTfBvHPLOSoJ4fc/GRgYMv3nQ0jqgHQ
47zXC257WiPzMKCTF6sp1j6hkcaKtVjsXx2z/njEx5ukdMdN/3fr3kdioFcAp3GI
eZQf+VnsLv0iAGzKMimTyzq+X3lUlqU/oFY3EgFjrp5i1tKXIRJBXMS0kU3Hg8iY
VEKGcoezF+KuHZWbYfHUSH7xsTtD+gDqxvGrXUlimyJp9zcPHLJnQhpbGa30imP3
JolvoWPxyCgtTl9vXkSPhPkOFX9mHJ5J8Hu2k4YLN6b9XD3EWy673vOGt8pgSS4v
RnQJTg7Y42VawjWKSlaD07SjxFE77HxM0amE5tMICqze0tT+4ZOlyGudvPq/wm0k
S62RpxEFkW5srpE7vjsgI8DrRUcObqaQibzo7Ja1sGZey6wU5Ypo+DCUpry2hd9C
ZNdbaKzPl7XQ3A87duE+I8E0Nm6uoQ3YErZ/GKjRfhJR6CAivwBInnE0O0sGOoNB
gp32Kf83QrJ1jTzjWWnKWYLY3AMo3ZLWhk0z7zm5GMxvpenkU521rBMfhB8GLiBg
ExXQm3Cwwm4UhNtrOQN/J6mAXeBN1h2BlTlCsUevdfHaSKW2BSjq7O2kpk3gYNdK
7egPd+GeWenpahQB5mcNb7nDDyXvenxEraJ1U1HTl0YlwguLeobUKdnOz19Q6Xiv
DMh420tOeWNx/Uy1fgdPSFu4/R7mN91JnVvN5q62hZEWViKjsBy+L046kuKhYLqE
V5c4EDmkA+VQ9HpKMpTKb9vE6LEd78lGLLusZ7zTS/IBui2LQTSPiHSgAlxC3KiT
6g75SWMt25NCCk8VUPBjvnukx4C3gcCU/Rh2UYhxgB/Fl8Ew5P+VdHz5CsCTHQhR
sCchL2tPX2EVBLJATKSokFbZ6uhRi3D653prgK8LJaCGaLCzzhHxTvmuItK947vK
exyD8a3igBvY6J2+SWJ2yxMQDi202emzb/aHfOF4mNHp+k8UVkMRpNuv46ZWcsJY
QdNCAUbwtd2R8fr0qGiZzjyD+v3Bkbq9GYMwxMFs3dO1GBmgNlFAFV2WHgR5wx+4
38LosY8iZ24A0HIi+KCXEUAkdE1ZjoXOckkt3Z13zrq07ny0y0GvyLioI3GxUoSI
PgfXClqKudNv4apoeCe9RN2F0pgxNrddP/21AtHj1kJONlwVa1AL0QFI1WWvfTcm
mIj7TfnEdccepblcqmfhKucrSAuncNHwEzCDKjQievFpLP4ZVC2Om/XOTH0Jvl32
QFpQe4mpSJS1FIZmKari4J5PlBHgL4qdFypdxu7AUNCbEtCchQsyMxtSaZ8B7dHc
9nqU+NrFWUnLJovEOMHoZR7aj8FEb61ynrBB3Z7nABmKKFNR8V5XrLRt6Vg3eJmb
DzHKFLxb4dvQfoHDa1vnxiA3KVkIObAMHaU5uEvVPEAmu5mNoih6OHkE6rEAQrVu
egpzDpIdIClo//48zrlD4w1FdahGuVxWHiYVuhDLbvL591t2ANWd+4XL09UTvlTD
ihHzNBiC8RrQMRW8J1flXq7oxfhicAmpUijJEHd1Y4KIOLGxgfcCKgcYn0q6bwaT
FdIfOn52b9JRSJN3SG2Nwyy0c1NJbTw9gvqctGitImCkVW6gnS+vApYtDgwZOW0t
0k+w/sU9hUrJ+j0/Gq/sCwmDkMBrMnWVgQbCmveMixr6ApIN/M0tr8ZmSnlSqVRX
PUkInsumiL0IvCAjlJv1IJWOO4IFuqE38Yc2YKYZWcA45cRdEYGO3rvuhWJZO+lY
PPwdPejA8Jr/sL1mTEqBBxMyINk/Su+jN770UEv67vRwopbKhy6GC4/c0ob4jDIm
uAthOj6gn6UuSAuCVv8O3NzSTC9to/GmteyRSE9nnTvNC2vPMs7KT3laVySIL7wj
iTGdpr6C4ltRG59UtDE54p68wKEtdik+/2plQpO0QZFl4pJwBXlsYswT/hac4WxM
DDAtdZC21TiZUCXnOYM3NWS5VMzBMZRWrG77cCo1Q7TAEKy6yTlDpcTeHhMPkQ53
QU/rmFW95D+3gE5HGLCfyYY4i786Glmt/G5WVvTKQGO/CyEIn/32o6L26QSq5CYJ
wFIseEk++wgxaL+pUhymEL7Sqej6d54dKo5mil01ScAVy0StmzPiYKl5+jPZoR87
DRBXF5Db7ncEWVmzIIXVC6EWOz0zcYYGD4HotCAXhRH4YkvusKDKlBTeK1vzySIC
pyFqcC0BNBKL/Uy49ZTS7dHBFYWXx8q3ZOWHuhjpYTr9DvIY8HN4Ua0URzVTUwYM
45+2ZMQHhHD1UBby3QI5vSh1BhRgDKAWUCmxEAopn8FGMr+BhTmXc1PxgLI34Evo
J/2EpbmyvoflxrURFFqoGHZ0GhTNtHcUQ52fZMYLOFb6YJEYN7n1NM3IRxuZP1Jb
dk6PspcnEOVT/lUSd3IhpFGtMZqjAH7VAR61oH0R7kgRe80/nADbIjW6ZVvAalNl
mKWcToNX8W2snDcPy7thgiU6yItsVDYV7S6rFcdhDr8eEmuknoq3A8wsh4KkUEId
rONybewmiojqhWrLVpM05Dr3e+VbKZU/RV15mV1eQhRRE8JnOZuoBj8C7lJUYAQY
F7JhErXIrCABAHXYYDxWzrfeownTHB3O+nqQsGOXPWBSDzOy77P+mM341+0WUmFV
zVAB3ur8O7Y84BWix0U+xS7BQX7m4Yu/BUJY/14uQwmiAIKBwdoAEaVBCYT8GyWL
ZY4RkkaDExG+sePQFXfyYP5fvl998LMBX3s3HRw0Th1TFBb9qvvvQtrrU8zKCfIg
vd2dMstbqc6Xpm3tVw+kvJ+/I1IrIUxPIbRpS+HMXnmNJx5PbPrG7Mw0kHAyf3Kj
BO9QWnnufD6A5wbk6jS4bmtK/EDev4VLn6LLXxELoJOyUHVFoqYJDjGhcZtSy8Ii
FUoluRTyZAp54BTT1Mu4Er2QK427EZDj0odS8JViz+9FEascqjiAyJEwI6/+tFsr
mFuOdhCv7WNZ7aW4dhlyLX2oVs2rSxQULuML/p5Fq7qcAViVE2C11i+2zYaIU4qA
j+XM8wmW/Y/uJiiDo7G+Qv+jBTUNIsXEHrgcz97Nm6cxO1lG1tbVWAEXBRNn3s6m
dh9JNk+zB32pjsSWwn3QqBRdCU/EsK2JZCOEdcFTRzNgz6msquyELBISkTP4Jq0v
DER1iCVp3pqb0N2yOZx0JxnUBoUWLGQdJi8yNu9GlNcw71ZUDGkQvDV00MFEDoy5
yYRxGdgyC1eJlHWMPZXOMbIKvqOfNn/N0fEgZqO7XjHH0R830QfXJU9mP535meKy
3c+WJd2edx4UvQ4WaenwrQdcGA1jmYd7q0kexfX6oJS3bGGAYd0hfsHHSXlsZInC
092ek+NWGpBu41rl8lLF5Vq+XlTAc2XekfbpDlwQWX02h31NLkdGZiark72JcAW5
zYBA/byj9+VFmyKG8xgZ6awUlJ7q4XaZrzIfbCxgX4fE87A7vtDH/sJVVcgRvbAo
Aj8TMkSElY1eMxG7GL+lwfooXVRVyMCSPzETVl1/TEuSnPyXohakucQGRJHZyqUp
jKGDGAAKygJzTtJlTt8idy9SEfOpkHoy0HLqqH2iBfl7mBQydYsZtZvisPaTROBo
UqEstYkCTBzPsQ33H31gAaz8N2gkdFDSYcyUTLwAL50ib8mqGLZjjthJ0s98VvbV
fA6vUYhJhCjqs53qbcQQ3/SSm4Jg2Vhu5/L8aapBCpXJVXbHWFsfsTPu+XqeSs4m
2f5dWLIXTZJRhN956g7TBKhdm2wTmijGZwDviQMPuuP3kbiB6PkQomYNewPM6hJm
Tdy2mrYV6q9gONM2kGDocuCG+KQo2A+Yp/hIRvHGtHB77tpW8bMaqHrYwTPRWOwD
605yckmlRQXJc7DbJ7mb2Hb7sx5HPj+SiWrykI3cZjEUEcwcm2kUJBmNvIY6pdW6
f68dEWt+WXRWtIO4A9dp+YHwtD4Ocb7FdSRQNYgrFqQWe9zZRwGkubth5FR7vL86
i8RCDjLLtxBYPTcNeX8Y/UlgKN+SYa7niFdMjISru3no56nWODZbWet3S2rbeUHn
sbAZzLTu3El46WbwSAU4sba7rY0s4XjrLMNe76xa1eutbBf8QIzkCYVSIwSM0SWa
dUar5KCWgqnI2W8/rc29O0qh9yX2gOkMnpRzcBbVNs36g6XkGbIkBVaerSx4UCJc
7o5KXJN1YP9My1qJxuBB1jqfX0rEvuPHpqB65qCfAW9SCHgRWmSynC7RxF9HsTjN
uPaPY9QqczHS1JomW2WSq+JAeIcr0etmUjV+tMpvK09x4YIxnmLnx66FRkKsklsu
mj1OvyqdQnXm6vwgOGlH2y2hEpK1S0rjI1GboTRdnxMRAZAvyzTbTByacdJVzPX7
2enwWdI618R2c+5yN3IrS6WcmCpqhOHFgvPTmlwVQY3Gl1QOmZmUrYQ+NkNvOI3s
g0H0jxhudLEXkX/rfIjTtk55skS7dvyNUY6zwP4NfLJ3HYygle8MlJ+2rnxD+Se9
eXRQ7hOE+zshNza29JO0IEYBaKFQqqgGaYNl1qv4SjjFFBKTxvzjs5lReLynpT3q
nY0I3G5AARB9mu1QrDypBLe9rzSdVZWKrhJGyg41SDqgbDDmAbyusaXE80opC9py
Yf8LpNMotjMt6DLGWkh3hL9LbrAIQGqx4gLDtth+jQS6s3jdM2uaYoVtz2+gF2lS
675nCmWN79s51x0IfkMeSdVlDLOf5uBKEnQLwxDTs8f1dPitvErnmjzEuCmLLlya
h+Nx4J4F+hXxEnQzaT+HJ8uYxv0MRMdeY9qn7SogMJiXYSjGdIg0bbRboaYFSU0m
G8GLYSq/R9O0SmaiWb5sghB3d2nfWbKWa6AyDeyrv/JJY3buEdO2FWCLjA/CmY2w
x8FVKV81ucQ2Uk0iyhtNuRSybcUTdKvt3Efkkzmyp+R0iRUaqZUwdvYIqSWscDqc
qp/bejpr8nykAQD5zSiBZ0RapSa5+RGAZDIibx6nLCt5zpCYBjzR/ploJVgrf98a
3S3sZ93B3gldiZJbqUdMTCvtTArVgEo2azppxauhpQrI2zH/p3mrr/RqiKCWZGqI
oo8eH5ygHQKy4pvDjJjPwBWpKKpwljMKcxxGJ879PKrMja7Eg0YD0ljDEOQ7FgTk
LLi0cLQ6kCHgRSP3MNIaEBECaZ/Mt4yZ/bP7ElkIiGcpb/aFy+gsQeFoMP6Ulu8m
vBuJDzdKFt/XcmMEsUS3pZk9nEry5gW/m5pX+4TDu37lmRp7OIWpZu3rNa0ffSnD
4T/p9JdC48ktz+ufSn2nBHJmoEwglwMS0+zba5PcrMDVi5mUdSU62/MM1U0VYv55
T79oEhHn/XjvWveMb+QwAc/zr9ZnYO+RRCYmlw+PFSbCbB5gxTAXxHlsvRbgsDtL
hiJC2kY91os3XOFSP4qhJ7AvecMadRtFiE+EUyqf133csiTeVw7KQnr0p89GduTw
9JvKk9AG8MtgS8h5FxBw7KghP17oXfpvtF+Q2plOrqcBHg+Hwdu7h0Lq2PioICA+
jFV1DWgwOlvk2YZtg1D32AyPdWeOX8D8GLxUqQqm5T5AOznexGLEaUv/iiWsrVgK
s+Ovmeh00fMK6bEjuRNKdh/DjDCMi7KPj4pp7hFwAekxb140XLzOFMFjfFyJlO0z
nTPPaKtSvPgrWswezVbnKQQ2pyW1nCI3EsT4bejr90dIQD3F01Js+ma1CzDAkDHm
c6G/eNy8KDpcNP7GOtuy08HiUG78FSZTbWYtXALdtP0bFEEz/5NMOfaAZwO9BHpV
K+p29nh4hv/yqJBTkt6pMKKPgKOWfYF729ZVpw2oAltd5aJoDThOuj0MnqVp/tIJ
b2sE8jBndotiiWQFJ5PwojMlUAW9Yo4XbzaLJzbAQA2HntFVP7yRrZMtE9ML/O3q
9qWkC5XnMMwD1GNHzBcOcppwXoD7DuUg4xy9DSXjqGl3XmvK8HUp2Gz1dqhAqO7+
46GESIox+P+9mjyK8ozeTbmfFxEG/MgtHUEVqOGuhafwXTfiMwAyq/hwKLhtI0Qk
NzMjIpn5MUSYzbTZm6WBlQ/16lzOcMlHWm/N47BCeyufBVAJmsMj/cGvWtWbFuLZ
o2tnca+fHp9/V5CRb0KwBV0lh+MvAHkhyofbXGJeMnDOsyeuu06Y1BtzRTmvsx7F
tqcgJB5JqxboyJk1I+PzfuObbNTnjyoYKBhLCEbTcDA5RtkV6vId5yC4UsTyfjUB
IkTOuUp8cnZWNgHd+Yq14Rwj+xY5DO6GoyEEwTBPT1faz0PTo2u3WIQWnsCmgg92
VoTh8dQbAUygM1G7kGGSzeMv1cMFE0k199+qaqSLzXB93eS+qoGAR1R4zNRkA1YM
5GfzBgMNBUGN+4CEVym9wZPOThbgvUuRTZb7W1w0tHgXMS6GkEGaUGcTTz0YHAa7
c3dAKmN3dyEuqYQxc7ZlidkH8f62vFuebhY3WLiqzT9dbO25cHlfLBqFPcH5jhE6
8z52R8M2zCppxmv7MjvKxFZPwM7JfLFuaQ4fttaf4cF/FsDSTCm56NVAwTdnEjHh
JdH8wCczttOeJ10PDpvQFMmBkLhg2y6eW+1HeGjGEyUiK3dhTz7yMLj3tuadEATr
pg325bxfEfAeCwBwe8vE+REo66pO9fy0zMNJAfUDJ+erYo5os0gDeonRcrOADNJU
IpYbpd3q9VoB81mRvGBvfZi46EIeeNm+7SFpTLzLOiHYlfSj4Lh2c6tXiwB1Z6Jx
Hdp47Ff38QtotpPQlWChmK5pLZjHxukz8CXr15ioq1aMiWKyI5P0CD1Bg4U8BvVE
1cf3aHQsEexIydzT0Sg3VCcbgwvLreIKGuzq4cWMkg5WQeOiRZr34IFl4lnI/xkM
a++fMFGa4kjqnVJVI4new6oWen7tmJnHZ87Pxl/fmcoiS3aXsHmRVenjJ0dyxB4W
kU0Sg17CNYTHv5JiC0RHZ2uXowBe0+0jFPjES4BfJyJC80XrxOu6M2m/BXEmrfgn
Pq7u6ifQE/ElxPnQaBIyHXGI0waSlfAH9N5n3X2JJvpF1jE2th5nQgCP/lbkrpQA
oK4ayGqHOqZY4hQZ/pMKiS6kWrcswrE7UPt2GLCijz9l1Zyj+5bLb1dye7TuUofw
JbrUC5HD2MCqQ8USCkFYl/FZeLPuuz9meDoL5NY6yiNRlgJjD1s9cwCzvH8Bv4tH
rJPjYFL/Z8M/PLd15GUhwhUhRzISjr2vUbEDDEynXxL6+pfv4CLYAnre26NYT0Ic
iV9itAbhFzfxNhS1PnJYb1lu8P5OcSl8zYbwoELb2/GbehLTxdKrmRYUnXXvA3XX
n44IRiGI7c3nP+etvQ53du+BdZ53BxDOakZhInXRtEzpP7RjA/aLaJQ4XIo3Xw3U
/jO7fmUmFt/HQgMqFLUWzeob6claitCmCnLkL/p3I1BUqUqAiVSdo1xXoYMLvzvB
5OvjUNDk23OyrR3WXXostKsncRWYH2hBi5IrVWC/Own7PICveoAM2q8ZZDKpHhhP
bMTftfKBPqAW0Eq1YpY6RNiHik05zd1PTGgYp46/WmUV6p8SgvCgFVJXK5GV3fjP
BYceEbJhTgx8tOKvaGeL9eEtRimm1VlDAQf1uS/aHYPvbhKuaj4i9MxJOS/GO//4
D3edDknhNJ0sd8o58lAOMbxkA27cOmAmNR7ag++lwFSQOdIuN/78VKHFB1usv2Kg
PE5GofDrGIO2ULfSm6QChTXOa9En0M57RSf7kjJPWPnvL8LC6fQF1crgON3d75fZ
QiMEtvIF/cSzkzWkQFLIwLixEuUzMRMV3K9Z688MEoGXdCLspPTlnn9TWCpJUt0W
HAXzWluAUflDZ4Tck2/bQizTD8I6PCs/axnThI5KdQR0C5o9pUd8S3sOllnlGL24
SoiC80Sesw2AWncCutQsoxwfwPuo/cgkvFsYn4ES2jkHpv4ajy9wqWc2G3fOca+v
LHX1vDuam976znItkDk3XMn1+CbH7V9P4g+ef7VwcYfoggSn7uG4V96wu5ankgGK
+lgy4Eo+Pf9qAzHW940cx0AibRY7CSfVIHNge0FslH3HWvrUcIWF7AZn120tNcQ5
7AOD311uZk7ISCdaMPsD6GGLYrVWp7Ip+AAikTBfqOaqoLmvFvQDHAnotjQWi+xO
Vso1sAK+ucRFA/O07raMNj8uXUm89Y2LbSUKobsJeJpurVzxjqIR27vq8YPOxdXc
22jb4OwKcocfLG12CSGYHnvMaERxY5ph8Y6hp24T9qXIoJDBNRmSGolI/Whu+0CA
5eohIpKplsg4TFT6bZlFOCY1cK2yX0XFR21gdvkepHf/EBSkws+zggzDk17uS7yf
zNsmz1zuFqRCwKEKS9j0O029bwIqSKsqb6A8AZJ0ZNFXN3Wld03XqZruKwyDg2Vy
UCLvgJxTahM1orznexBjUXKWIiMv1Hu8gREzLgvUEMn4VwlcKzJ7A8uqtDtMp4nK
EKXg1zip2SlKbZ0+B08SL/zwRj0jy7jcLmDGz6qKTYmqIv82WHy5oA9/nlb+O3Tq
GdlhQ5b15yZtjLHe69iOfYwqaMSn399f96jRnxE7tlxf5KuKBXqxIhcJYu1gWIih
m96ikTmdm7olllc9l9rhIqL+RdTdFY/C2FH2QaRT4mBKx03KTHUJU8ja9fcjGKnV
39EB8xGOBrlA+Ng/mzKYMigZuD/X9/n55+eKDw2eznqgrmmO/jlUmW/cyWQ1H2j4
NPfvorZXfbSzTlWIeGOZI+U/xT8Lx2O+tgO8xFYhm1mu8mQ7ugN/hQcJChPwYg10
fSp4ADwC8jVyJ3bM/T7xi77GzV7wlfPlCIZ58vCM2caA+1EzuWpGf1QKfu+oaPYy
/8oV5DicQZB7PlxhYl3yTCwgOPa1w46oGGl1hmqS1U2AXOI22MAOeOJw9Qe/9oyD
au963fiV9090x37mP4uKGXvwi0lbFIMvoaDU/CR73YZpiOsN+1OS+GBDUNxjQymz
Obx9yJ9UwP/FabsqaW7r3YIqlJR5qm3nHEBTyp62/xP/9qwNB6e3XJc4Ap91R/8V
CVsOn6hvGzZyV6UMmewvTd9tjSZ6y8RylkE1226iZXKrB49eohXeGGWJwiTIObhC
cNx5EwyknmJb6ZkcLiDa6RKhR/FThfjl4rb1I9XZ0hQ0kB51gfWY9ZJdByv0axZ/
+4EoI9rq1kxqoRRfCa7FO6lLbyWTRc4+pSA9cxiFQzDS1lgEB+Kk0JRPBrAvv2U2
RJ+o2VWPCCSuc7Exk9snyvxJyXC3QVD6X1Zujw9+pd6HcIZoDxW+9/qvrbKD53K2
uNGMWHAVEsbosYar0JOi5ydrvjpcWOdBc+QQ5dKzcUrcGR+oUR2uCgxXGznInXKw
4iZ5kMTmGuZuSVU5ipwTlgpcFG7LzM59DgC+K2yd5Mt+J9/gPbEPj6xtTty4N5fQ
NfBVYzKASQT5TMsT5nGUlnWjiBLcs9+Mya8BRO7feSgWsPzABPXxYta6mUvdWHyS
ArmNKKyubdT15bTK78LnBNRT4D8oyu10x/ZJdq3XnQHkffDLOjgSJJeSdT2QXFPf
iDFBwqeGHwU8pTbPbnaF5xDrTrpRFF5n7WixAsZxR629KKaKO+7/7bAtkJfPvsU2
wwzX0YQRxD0UxmLrojJ+h5Vyr81nQFUrujv7feHROC7+UmJYQSxXN1ZMbs+4PdRf
CCJ5x+JeXFiA7lTKEndPgM/uInMbQiPsAM/17RSCHfvBMxH0ubPwXsbp1ujqhUIK
NmSkTAj5QKZc4q8yXLNcqksDp7UEsxqRO5HysNXq1ZTckq6AqR+PVwMvoBs54ruS
LHU1AnEvDbXYcXv4YOESXZ3tNza/k+aOHkcRRVN02KUypwUxpk9ujTr8N5KklYle
N5/W2EUjy9kBYsAQ3OFlLVcbP/3qy/KDckzfmLiuQ8VdCqKOtmCvpoV/dm3C5zpw
syYmfFckqXz9LiCOEQqiJk1SKacVpKbp6Ah94AmRWMpr0mABkPRmJWnj67Ue/tmh
NI27wfVLbSpnlJAN6ETVDismpOiEmcDQy67f5SSYFUd6YbHyl8M7MAdSIyI8C7b1
W/h0tvUbsbbM5Ozf1mc0lIK6VcHelmsx+MRS2b03hK9T4QitC5xBF9WOiY6A77VU
hFufSfyx44XiqiLhJfqATppH1FNDODjnho8wlQsedKdQzuBBQIAbOnttVIWmGlfY
8n6T1hI6qJr5q/T/bSSdYrbHmhIp/hqoMHJFP9Us9Rc5oNEalAm4Anu6wLi9EVeA
XzrnWiBf4rO0gi3NMBg4BO5G0UW4WGldg/Z6DO1Bj3RY+59fJIwIR8HW3UYXvzYG
+5qXEOKowkDXtgNuxLazk4H8pBhtQwIsCK2Vt/DtgcT0ZcfiYgOb30PywlXuP236
vITSn9q3LtTai24LETuTYi8aQOnqyTpwGDozpjttBNMeQhZGcFG98kJIATaxeRPx
QT2ZZrnuF2U/syy0SLNOdwtBzyZZYUc5xhPBSpZFeMy4xlKRAfj3DeYsGB0RiOa+
e95uoJ41A7s5Cf9h+AnpJ6WEhAK96qDzqgnfy/7w5T5uzWJ2G/DXoSqzNIAT36Lu
v/gsR/G/o1M98FjN5cgT4r6tLNbqj9XLTPRx1yvNPRRXdB0Sw8pkxlKVIc+CfVBj
KNWCmnnozJwUO5Hu0v+iBaQHz+z4+O2hrCCnubUZ8KcQOCqj2tYukB6XcB8Ha2lX
MTQFIlJmmPir92PLxzVBEjAqzrKnkjhfCpb0PLeeMZt38lpxTq5TtcLLr802751V
HfS+Ld1vU2dwsSGx8JJVCscGNaQEk/Z3T0Yq+1Oa1GM4TwoqyuViHRmqu5rCJKST
ClHg6wrxA3UH1QJ5R+qyPcvdY0f0XHQZkl65cDP4s5qksIecctBAFYS34U7Ywosf
pUwoGuXXlrgbxlhYSUScedsgtdMfkcOPQ5WyTkECYjuY3knnnX9NIg4rP0O2vM37
fXpt+Jgy+ipcjVmsnPGTV0y9kGKn+91rZbdVCLUBRbaHBNYCngJdaTDa8zOvrMlK
lae4y9GUYwOl05PEuBSuGmuNFXeGPP8I/yn60uD84b6yH64Dgt5wzJslUzD+379z
axo5rCVpUO9CJrifpRFqp1cWo3SltTRXC5g4OnX5g7JibOCP0qmQEYeHDt2Hb2dc
nHhx9uGE4mh+chA+DUhfmAT7K6sbuGnmmCH/B4nN87XvmB3NuDWnSM7EX8rTi+K8
6UKapjDmaIoC0dyvCJlDwZbcMvq8aWhb7dPZxcEJhw+h8DK6fANDRzi3VWzeG/7S
qSuQJe0+jIfGJh2iZclZHjh0TPaHTbDElWjStz/oUPQRj6tsAnwDt3NZyFcuScTL
5vjM3C3z5GQt54YlYvLOB7Vcq8dxA9iQAFq6WdtvopdfcjrbgXORdAjtPkSnh89Q
Ee5YaDRqadEX08U/tZrR5HibXZzXo/LCbbHe3s3frBoswnsvijOSAPm3GGCitxvL
AIMfC1DUbiN7MR1eBVhFFZap7dS/780rfOfCCP8hdCLpjzJw2TUBsXettirsxwxk
6nxfQFo7rGv7grJjdvtTe/iSC3kcfXTyG5DHQ9Hi8swrn+Hktd2mLGaHlOH0KEdr
dSo8+f2lgWMFKNxXg4c10GVFCOogTqNPA4YGViInGK7ja7WIyB9jcrWNENDpq0/q
iW1XKE7ELuCStZlG+hECHaKLv/EkRRLxNYTJiAQmEM7fw44f5QAh1AbrCZH7kB2s
VGSXZKMl+l13hnm48WkJBkP9SNeNrDscqbeIErtf+ewiTnoR5U+CeZX+sESTGgyy
C+9PdrBW3rCyqiNmM1RwzmIZ5QU98f0NNXKmIwc+c9R5Q/LrbfiKZYgASIqyU1aL
buY0KIcJjcE4zOI/qlx9Nup2Ff5bxkUrpyE9WBmkCylWX23HNplLT4PGdOAj4SB5
1/xCrOTEbxf34Ang0RIQHwSmQZk2szGPysbwK7Xhbmvvr9oHQM0ErdDefP9xDfOM
TCDHvVxin8OJvc3CkkxT0gR3gwE5JduMZlUUFXAp0NRHUPUOyn4j3y8leKrNCabg
SsGVzm7uWXTybN8VVDS2ydpXMeRadx79ykxMMI+6TphsYcNf+5QIk4pkjt4OfV2f
E3EbSARyYDwIipTrnbfm59oTdDEFxXA5L4iJMagv5AzY/Cys3ICUbc1H/wT3K2Pl
pLyVS/y8QY9d6e3tZiutxsQ95CdBGIJsuevMDS9I91rQWoEVzIfcr7qpjY080+uc
sMBYuyIFHpl2Im9sHfzUgwBnMHd7TvmSsKXQDypOhT0cecu5v4C0eFRpvpHWolyV
5HQCvqBv9HMHVljmndmDfdtJKOzvc+HVxHIFfMy+bF99bCimxZtN4rE0tEffNk3f
zYWlnEnOeQrSiLARtwGXUfpHa/2kL78ZABhqH5UMZee3Gu5OndwVCQRvco/IgtQ9
KzBc6GQ6VY1RE9aKZd04tqbSjTg66glCkVKy4bl9AcoAzkoskyZp0pSXJg102+Hn
RwfMjFZbkh9ojQwTW2+/LQrUccu4jm55ASlwHy2u2OfAI2Dyybbvqc34CGxUPDP6
LuqdI2EQ2euIvubvc4YFweDzeV6DKmS8o5URv8cKISJXvAeZehzSPAlgz9/5dukg
C9TX+U8ks/fb9NmkpEwqRkIyJRwq/a9CeCXgTIokjkLMFU/pwMvU7EgfcaWPiC3I
9cFrZ0swwldlX7gAl0F7nLG9yoFM7ewv3AUP/IxW9lQYRDhrvkcgUIv2+8q9qs7C
aGas/aYXNCXTsb/Ari67qMNvsd9BJ3yjQCL3SOtV4y2P213+LlazpkfVuzw6Nm4t
seeUV6lSkNXSyVoMcFEE6f4+D/wA5sYUD/nez7i+8gzqJGiNf6mvwDNGGPKwq3G5
mh1Z6hZec2UuiBrWrXh5jXtH/dU3vCmyYYXygTjq9i+kGBIYciGZWT6Vc9Q1IXl6
FTgDJZq2u4HlJfpdqAvMqWwJnWwVnuXb3lRDzH0LRTiu4v1g7TUIzxQQcUO59KHG
g5Bi9R9+b46UfiwmOOTYR3solIELpcd7anujccRfumcwh67Fe+Bp0SmGEFRqQjAB
vFk+kDzVBZ9J5LkGX85Dt+YJMHx4/r2ZNB+sxsUT1Hs3J6+8q7SeniLZrrF/qdhV
MblPYfwbey0DP9hgOverFkt1gsEr0T6jrqCUkz8pFPovQ24+RZcu90d8K2gnK4zt
yeKmvaU40y9X30+lqtBwX9BQeWk23lFhKmkdJ0HraCmZBa45SYrGgU+Nt4v56kcb
2UoNDS8/1jrKq9B4FLhqTSZJ4JvaNp/9QBmCZ4d9jQTUdT2uKnrukG1ZFGzv2WFE
gxkNnRpTgozCNMPma5CI8SrIJPdg0NmEQYuXUU0nhKqR/VR3bYmKu+hKJLj6R1L8
OJb7gNizaUwInD8ZYH9CkbsKjYCya83dlzti9JSbQOzzXPfDCJ9TiMG+rDQY7Vf3
y7SCFqDDY/oNn3Wp3h1vx+QUhnxaccveQbsNEuQyD8BhAlIK9HyegDuigW1RxOhX
xckX25QAw0yCaCrOfGIpn6Hm0LZMF4uKRBneaV+6lJqNL/nxAz15rgYpTx3kZq4V
86Ou6w6uKcswagVi9xgNKEAfURqqUNdmI9fQVRq8iqZfgFXLjYa+To/IXJdgyZna
hekRsMM2iDy6AKtezMuBL9KKTbQndc3OsFVdEyJctOuZwg1ormZiv29xUT9ImKmO
7YdHAJxYwoWjrTkD8KdveWOyu0EpijPKZCHaaVHmW0dOPMp9Afjnxi3qZfRxmpVS
WIoyJJXTw1160tTn/kD0T23W84/AXtvgK6GT+5MDA0QqxklI0ciWF+NINMkbo7y+
6bNZwyjo2QpikjDxlal0YrG/nV6QKR939wq5TnVk4YBp/BNCoMzXd03Kg5VLMDAX
SeotDSWKgBBT0zobuhEAMsMeQDjn5cFxLEs6PdaGMQZb6rhPPcbQ9dt1q7GWHngO
yPavzsU8Vztjyrn1WrHEQBJKKFbwmV3tmbztguti5hNJ2+Y1mVCnW7MF2JvKSKPv
wP0jPN3ywZ4dEh/M7tLer84tT4yybs5PBxiYjCaPQI1qTo2DWhVTLuaWLOBpXV81
Sg7ImBfPjwhodBETriRDUQ33e+T95XDQ2mlNiIXWwRm8BxtA+v2SmnDL+ZH6jFc8
JJ/XdhXWyt2go3xuaH3/fmpUfa4nYTWkcaLWcIt0yKcFRAEFy7wkZ5rHeHjUoWE/
BQyQh0y2ousLbyShoieuUOgknWHI6UcXm03ObMWgffN+az7nuc6+N7nvuQbMylMh
qPqgfsexYiqX2WbOXfbRW1jRySo3JHvAJj/l5gDHRR3cR0G2GxQxfWbeJ+4DTGpk
V22iIXDXqNtI4bjqkDRZaHiKEks6xYOMaTtwQ07QcEv0MN8Hrz1sRkbiDty3Tb2m
bhBkCCjkHEeZinsr+MwgnaeeTMTRyRErBYzahbvHTUqnAX0RXYeBf6Si9RlgMQ1O
+gLHphsRxXRlXUjK6T9TmhUrE84DjarzROC4ev2OO98t4ko3bSX2gNejYxAE/cLO
Vtk6EVQ+R9PmG1iBdF0fRqdEB4PN+bsDL6urQk4BPgX0GbI0WXHFuK2KdDRwM1sK
hI7QkV4IIeZe5/6ojuwRqUv3Edtzk6cOXKlqzMCNYoj/RFnYHvWcqvODRkNVgOQ9
p3BnifP3zo7rtVws/Awh9uR+cuAnVz+8B8vXlgNkXdWRIeAczPpTJM6eiHIiI/j1
MxTvoxoWSqMKKWO796QY5UUVmxZ3R5Alg3leFJ2gJox68m2uMJI1EcyHLL8YJX5R
gmXEBwPzqrNUolSZQaZn4c+lQ0pXXsbwU9gQOQCiXl13yWEhe9Hg6fXKScDU3lpf
8+AOb2+/NAWa8Fozi4GzUEC8CckcLYfHDH2glp6+nCwd9rgdhQ9c/n9ABvGNgXHh
JuzYLOjLwhKOzjJfUMBsIwr32XLYC9SOtbLAkXY0DF5ONe8N/CJonUizn56r/IQm
OMffYHiU8Wnkz6biqxvbQWtoFvL11SPlGmpVDNeloEpX4JLQk0F5eiLqfipVEOyH
U10fVBGf7UFrN/2Zacs8QZRmwGXf5vZ/jboza8lE6NxAAAQTstotZ7ltCqCUZ4Oh
WpCV1YynxdQAkLcAYQOC0/EuvKTfDZ9kTpHmvZoKgk1QbKu+brbgeRyZA/jw/CXM
9mA+DBQiYm3oh0KSh/MFZt1FbITYn9ClXzmpnGBI6/f5bKQ5SQxuqTG23NhJOQKB
NEoHOhFQmxkUY3I9w+Y1E99JtVeT0kJ2OYe4JKlM+7n0PPnl5E/bax0VHtWkjB6L
53v7OtKOMJRwMb8YeeKRWIfS2ls+JRhtzXoN550Rh8/pmOCsttecxXa3PiP7hwak
UMb4VIzza/Mjeu9a2537WFvNX5j9XXVYtjgid2Hcab5VnFO5+YlQiZv2nE2sr3rv
QamonoEpLwk47H7qTSbot9Og6yN6Fy2BT25yGPdUaEHHtxRLR2RfUVAQZDX9DQ/p
SEtw2B1KqMv90utUGdMFD8zltNg7WXAlPkVMp4cvkEFqq7oIbrvBHWuM9ZZ2I/Yf
2/yegrpuxyY3FkUCkTGBMMo5QKBu8hZ3C00k1g06w0mJAL+MYVdFJ9SiOCUnzgrr
bEFyMH07d589g/azoEJZSc6oS1eCGKbnnSKQmQ8nMYS8rBXZw/RLzdCDkHaFFXhJ
re4ruLoaQMM4hl2CLEGfEYja9R+yasH3iZlspUIDw3XfbI/LFEZ/bdj6t0HtPbhW
09jFU6gKhZB9XG0UdqyIe2eUHP66xjLCvmndxmcdfTJfrcnNbrC8LXWRlspY3hsN
Zt+/LHfAvWp1Ej9SkMmbr0bjYfk0lnG8cHjoUleKne7sP0HC28Z0PeEwiyNgseAo
kDeIvabvZ31UG3DmHi58y/Dy7q99+Wt5pis6lGzl89pryExbfiWArYKeP7f+2NoC
uMvKpkjsihGZugnmy57WHTMg9LmZdv4XvGTXtBj7Ra61Q6uylXU8ZUDQZDru2NaL
E3YMIp2Tmz490r7ZZqvKjufWFAsHJ09OrdshbSgSA1wTtHpjfL6pZ2q2qMjQVB60
iRnttjRQFoZ/kgtrHTq8dHqX9a4t4E/2jTnUa/CXYloiISPgut9k83eIkS8c+S4O
4ccr1s0qxEqeeOhk5UVKot5tMY/JEZyNTHA2Smv4PT+0UZslMIaMNfh8cB/5TtGe
sfZkq5lRxgeVKVcCSckn3h/3P79Wtrf0KypycsQaHKw+gfO/jb7E273tXMGLsr1Z
BVXKFOIvz088VMDHignh3GaoT7ez8SoVqEJmHBw3NiVGArWdhrhC/qD4HcGnbZQF
j8XDJJBlWXTBmdR8lw/ZcgzTLOsvPLZQ34IXhHQYk1Hvt/h5bYs2ceFQVXY0U6u7
x4zmsbrzhzvRupDVmss2qetLYm5vZYS7qzp4HperEZ8DZZwQiDxLdtMSdDx4YZkC
BSajJ7bPwwxo/gUkrgmLQTXwiGrKazKJDOWIpg4DdvH97e5lFgsQxg6IYDvt5aA0
lJg1ElhkJjGJJ7WzK5Oa26YxvgLU2RJDeO/BoXryP6s2F415c7DjhzkKUOpnLqOF
T0VDhzL/mi3iYR7N3DnDiVUuvnAguIMhppdAOY3M1GjM3kd9P+gRafQBG7heOIp3
84Re0KSgjTsiSYY4QSIYsijYM7S8l8+A60x9tTO+dkbH/BnBJBbjYoxtS7liQNJd
RV5Kf6yqPfeuL2hULcaYjO5wcGTzMkLr4EiqLK08VvzQTdgUKSOQ420QP93GIgtT
fbDteLZAauYU5A1hHFZMDh+7AxiqYVYIhoIETt/pg+dFvO8UQv7hTRNT+8EwGr+M
hzaU2PJwd435PoS2xgQmKDsibG1ZrWHqbs10rAnwMhGhpUT2qZ8bWW3/HYNOQu0d
kDOw/JwNZiYGRgqyLawSnENKyWXmNRmRR6e2RKNjft3jdYWDeN0tJzuqwNT30bSt
n3PZ/OWfNWxE1v6MEe5iyUWamRkr1zsbj3xJ7MOT5bkKS9WhG3ZXQy6M2eDnqIBK
8MX02x6QYwA5bx9SyE8MPXCGHaC1gJTE/T929e4omr9pwzLIh/XxBvZfKl9U7WSB
PVbpruWcFoB7YEOxKOx8c6agDBKK8Q8AchGjmto+kY7EJj0pbW0rZWr4scW8GhvV
RGWc+nEoeV78/J08CbUvAITk6s+0eHsTTvxP5AiIyFqlzuSA5mlaae5jtvCmK+2E
6AAk2cBmTf0kbQmwGLWJ1MD0yyAShUJ7CyWOcCg+mLDCOtfQBenQgxFubgrZOc7g
pYsDy8f28ZTUXHi3KB1qZXI7LikvjooHm83TgoEvx6O/+9kYz6bYouO4o5QqGVIk
ffK7GnbX4z//9W2kFUsuSJVRYk+1oK8C9IUrwflWyLD4NhJW8JNSOGOPo84dkt5B
HpbYLSw4a+ZlKPjKidSs4g+Y/DA4K1bY/iocaiZeQoQAoWBoL99zrbVIjdrs8+gE
j+0pZHrqxioILTbalDPkgtdR6bsd/NIwwP6cm4U7cQuduFkWXnNYiRlmOi7VCIr+
PTjiqU6lQp6CNFFqF+LUo3ufFPr1VgemUG1CZ+648om3E1vXEiEhoMlLOhFNMyc+
RtpsrKao2ikCL/pG7fOCdmaS3BpEI2bHwOpixNKp4mwH5UggWle3xKepp80V/NNk
mlQTBf6KT+rPAJjgDJHHeg9pLQonW4wCB+cPF3dKcp00aMgwdFVei9gPBU+qUkPR
awJwvx9tjA7zf2Yo7Usfav1EAC54Kwu9/zXyBe6aELsgiye3DwMjn8mmkt86J234
6o6M06Xe9eLwGC5glaEXWXwNPJfLuATDklZFKAHYe2KbCuKdTDcdMPOM83GVByBt
0HGmoILI41td4raLggR5waQeETKuECV30Edljh5oyChDTsRBkL8dy4fehRwFC6h6
c8beJ4t2DaxdRaU5/KzFm4EqWSeRBFoH5I6VKkbgBOS7sOlolElfTgG0eVWKxx+R
v7Hd1B66ZucuhZveyLHnilGO5IVjMfgBwswypTkNtAYSQzZYcfCQ8iSaWe7Hufra
CpZUOYWWTRvCUi+zxWO9HBUYeo4P4MQ/vgooYYJ8u7AwdWB2+Y0IyWJi/1SmIpOA
hYESxJoV/uqp+8BoIXq0V3CCJGR14eE6QJL2QOLxyRvgf54c38OumarPKnYRNADN
HYIn0xMzK7ElIOh/CZUEbaNrXosi+X0p+Gi0Kv3yCNt78GGXzfzDftmYKC1h60ct
SZiWbkTbrV8qocDQhPWBKe/uQAUa5iSt6mUsffSRfAYenexgxG4OBiluzfA/E+pQ
0AwmaCLwJCQqDnnuvVLU3lKxbeQKCn+i8SNGPt3EtM76/w+LzjqgQUlWe3kG7rSX
3ekjdcK7WKlKl2s+GDX1mqYg4+d2pnD63S3Fni30xC9Ob2C7clunW3B7pyQQOQ7z
R0bdjuKBAxtT/ST8BvGj/HJu8G54P2DB+zHUnSvuPU7Unnl/2fAyhpdki0dlh+Mr
UcjFI/s1DRs0Yo07xngk4kgr4Hf9M8ctd1LdGkHiydX9BZPIBXabkheV6F2i2C4F
9l1CJSdjYm5U4DZv+Ri/ah+AYFTEZ+TQBjJF4JQ/eRN0ZCfsaz/VnfIBItCGFTNm
7uXXKVkzMM34PKosinarhB0I1a9bOYqA4E8r0WDCPG68VeZ521YXP5GJJ5UdUVKK
Zw1feuhd0qZO553bGuqpR6Ky8u43ZSPccp7QwfO3ZZkmg5NmIZGU6jlOwRXHnc7X
2oSp1I2x2seG1MVdChWX0//VBfZY1XwgBNwrvXTyrCzAoMf8oJDQ2haQ/xyyLET5
A3XC23h4A+lLdYiDiij9s92FqiuAA2l54flZN054Bo5mrBf208A+Ne3qg2eaSfLO
haoKB+OHRup/YnzeJoU+i5omSks44L+rxw9jxA0yzmRhy/UPgZE8ra4RWZLPj8Ln
s4LM0U6jmc9SuYYSShpHLULFHPrI130v6A5inRMsWIvyJVmvQhPTD2qcRJy2Sf7C
LKmBMbTZ/EG34ufyyBfTBv5l4wIHBp2Aj5ONimOu6VDjUd97GT/4yu4n54XPVkf/
U+PRFjcwSGPj0Sp66GEI89/0ezYBjIKASHZsunJ911ClyhgrFyIMyuSw/utossgk
0WK88iR8FS7SNjmpf8O1YVakdmgxyFpwcxMytODFfbeFszS67AsClbWTEb6vOcDG
iL58yPnC8TfmGUPE5Hw4fkg9c/ykJ+S5/5nsG5vAsGLsxBFzF3otIN9RyY22RXup
I3Nd1/xFKYR5oFjui/Uv8WvxUosxg0dEb+RELMoYxMbcDI9jy1wy0WYm+KgC8mu+
ZazfSMafKrbhfhDfV9PuovccADpvVnS5w/Z71aCeCZp2oBMV3DxkuILerWfNLVoh
vliNZ4mrysaj/vTA1O/04ElL6FGFzfK+cXS4NLcrqqWzPYNwlwO89PcfHt5HuGs3
Lts8bkjYvz/UFalMvEEdObehQs+lDdFMHT41oTlG/ziIqb128ifIv5R1T8grjwfX
uya956FJfAUb+Xrkf/VxR4XdUF10jjaQ7CB2rK5AFhPCDPplyrL/Kg8hr7KxZpKH
VDpIjh5J4BfPU50BLabdHCwZIMPmxT9sRTjG5J8ySbxzOJ/p1xwk6uW0D3paDcFD
xABwp+DymlD9M61J8aEjealESddtBn/iiSDNS4gZzrKRr8hGMu5SQJUK3SirRiaH
Fq202cAc0dPlL3SMl2PC025UcLaEIddEMRYymKaplrjjO6naiMoTeUQMp+OTFFY0
t4I5JLGQSZhlHNpG55JQOYOlAzBjNAjMVxwT4DF0Pri4JF816bJoo1DrfGWauw0f
S+dzKDYgt6u3m5qH14nfTy/d5yUJcDwwzQt4wvU4bzbWoMthkE0mPD3Vto2f3yPR
ze6viYflAaG2+YwZY9LwMI8PdG10pfj5dcfZYm21cS0OEmzp3mjmMrM0SMz/5QY0
h+3IRY5ZaJel89fIVbMqMDq8r41sbd69kQrBMYNCuzmUY1bZ625YuT0mix+Ygjvl
FrSKSzB4reUkeiqISOk0SO4XVoiWIpCWQ3gp0UISzZny+cl9uVikH/hXwSwa+x+P
sruaKp3RYJQQ9R2Yr0awvF4B2CEZRGO48khN9faEz9g0BSCCnWjaqoZAlNqcEc8u
T8okqi5nADKLwZwjdDrKTDSrtMNOHyqKS4/c9KT7jR03XZzXQX6kYCoxCF7uJ0pn
zigah7mTfBMJiRGxr+w53knVFecTwzpL6IlzoNByOQVGqyRh+STAtH/iZLqxz2J3
rFbwoZA9JtVG6cAkTOVhzqYdGUxvNPh+SSd3RM+3VvnBxaLXN0c7hR2bAWSJOIwu
4nFLY9dVfiReBBhMyDyI89O0KbGqp/YYPap6Oa9Jd9NGp8+d6Ww7eL0haDYzDNo/
+n4NcKVYzYqT5TNGHAbbOX4g7P/elGO+vfq0mUf6A0PI1W+LuwRRXuqFSRybu98j
+m7YRNYCUW1vBSzSwx4N58qpnaQm8lB2kqqYsr7YA+fdDVAbDwXWdV1ATVzL2iKL
rC3NkmoufPPT2qFSdsFqhNlIIGcPdcatj7U1HmSWFiFbDnTtuDuXkPseLpUNnH9k
aOAlYS8nDnU2VZxxURlRU15BCv+UJWW9IhKCTx0BZwnpacDPL3p+/O7XjKBWgFaR
Eu9LgfQ7t8E1appXNHyHHuHPrqBuVyLxJzL9q3IySZuMZeqPgGHLzTHdgz7kjmu9
9z+gcBvsGDdOnAZLJaoJRmHlYoILEAwKE1mOg3/wZoeIJNNgiaNmXPCqxiGYoCtC
QsOVKUE6oTx/qbfxiQ5GuqonZQFZgSkoAL5W0Frj+eSGnh3IUDifjE2QdaqsE6fP
QJDbA11/LOSmIeiNgb+wuXRpDoS1AQ5pRyWFieK6hFHg4bEJujfltjkT7AioPgF3
JycKlgj0f0925OgjKYCBMQ5e0/BoTu0b6ToVVY+1VoNgMQr4OColxqBSzt/ESWPq
tZDIDtKIobUSswNfh05BqHPMYAoq+zGnK769hb5lKlhy0DqaJlGHNwe+vXEMZuFQ
3+YpPHRRwKIgI3pAhvy4OcqDR0WjAkDaOtSOcYSh6zPMO18r2KOMDKxtbtU2k1q7
EdKT5B5ZMPs/bN3oARbDg3lUixts3uWJ7rPMnEEPoYdqd2ZIyOuRnbF8ouRczf7g
5kTKcOi/NwXSWx9ZACf75DLZMoJtuPIyoSced5ps7a3HZxLhbQtM39b3231Wqz/H
l73ku2txqlQOJF/0pQYZa8+lXj5db1Uhh8uiSNSmu2CFDnBhV9l/MgtCaMfqWGl1
BWf6unuwegGTu9vXZPZZ3N75pzPCIOoKBcsIF9SkAPLVk1qGIxH0zWBpgHxVe+jO
9uValefShs9roTkezjXZYxfRZnN7DiiX0TJC/uoB8XzFsLtjPhUE+FOwRPdiwMT0
qFGODF3c51yP5yG3ezmN+JV8z/mVDFVJRca/AMNL0ZC0g8yjvnPyYh59UyFJR+IA
GxTuUGL3VwzUhFIrSIr3Q9JM01VyHF/lj/LclatBsRSg4COgLMyBMNmk0RgITFWu
pDVNKjM+DDEICWJ+qGvYnzqYYLFNetBE4lWbx/5wE6hCdhNtapurFcNUFQcGNFSq
2T658VaEmUUWRLqtdKYeblfPSLVSMMrN8c+7eNR9Qybt1S0UP7Qq67tqDh+cW05i
Oq5LAKgxmOJYRVhuoi5dgwtWrceoSjDjJIy48GC/Dt1zGJfZko1CKLIcKPqEOP9B
n3jb6EccmvbtUJSqe8I51okHad/NHTnrfUA/nh0ZfQhv+s9qDRC0pc/scBK+MSG4
3C5fOJM6cr7iwAUpAxOi+E66Q7EvLmVuOkUABsEAdsHp0gLiTahpTA+tBCVy4ihT
moBxyJlksi3n4U5T/D9/s/8qfvj44B5gHvS2NkOEXEmwS5qgZDEDKjQWxbCyDKbG
1EI582jII+hqdWXkrZLJ/JdfU+7fphm7calxcfef4WDS1YiYPoqA07tfexf4hzjR
QNYexSyMpdH+oRA+Afs1ENTkFCV2Dz2k8fkFGZIVqOXUKMy4IkYYM64tX6IlPIf0
WLCzdYxRfVl9ZJ4seke2e/4+xX0CYd5U1258DDb4qT0kw7TY1CVAeHnvrjTeef1P
mOdNRhAuFF16j7w8igYk3gTxG3dcNJzmhwpr69fXim0CNX5B0c8uIaP0l7ltF21k
FvcHAJ4/w8iYBsZgAxXdsGvwVuI5BTUU7WDxMhTl7/xTteS52PBBzDA1/DgT3yyp
vjBVoIrIWFbg7w5axPYpfsx84EQub2c3oD1FTP8AyZAL93C0TJtEgmVRyoGgnDt0
G7BR+mR0tBHUbk4aQS3AybXHv4TdrGN+mws3UgUkb4hlGX7qcKkQn+HdRg/mKuhs
msNH8Dg88FbBLUXbcxmE/CAGUIn1a8jZ3K6/5jfQsnDami0odbhcNqodOn+cEeDT
eBM4Bcl6tXfGIrzofvTmiDm0v2RkSKub/QN1xDTVeKjMMyb0rq+88UzKb7IVvsBm
eOpNYC/Y3orlb6WJpWf5bv+8bcPhqHfpcUchp/qLiY057/ELl/KN0G3F0mWB29+s
c28yAaR8pgdL2Zziqe844BfFRCIe0WTyzKGKX7pG1NvbJK5dTRy35GkY8mEaNhC3
1YObxkeR9Nc8tWNkz9hDSiGx9apwTCb9MABl0aWXPpkgPLUwuTZNgtcQ88QMpqQs
nQ/HjlrfuKX6aldDUWToJpcnC9xmfxXxlY6RhYbjm3z0HFWb48fiNAvaTBaSwT8+
Vr0QNL0Zq/KLroacMYDKuyDu1tEg4twJbi/b5uwMWvmBdfcvBVhZ9PGAR69G3dtk
jIxsiyAgEZJKtpvaGjEZ2Q51OPweOTOgedXkFy+T0QD2y8IEDFunoKZC9416q3It
RHh7vNxydPK/NpX7Rhv6lYqUpHtbwv2u8DOWqE6f9d6SsYYUTnfzqdSW6FulD/3M
LOgx26g5WcwTrcheXz1nzohQ4a3+wqK0QojbpZ5Qi5PUX45EYcES4xrWNpxMUKrI
5Y9udMiDxmdLQWefmaqIseqJtYWsilQCitkbU0wExXx0rB039F6nmSvtVvA+xfMU
DgYjcJBuJbuFOPxGK/Df5t/aWkwJ2HPZKg4iDFYo9Z5M0k63TMYFML/Ob/2QrGjV
EZ5DkXDkCirgyrErOAtDmhjJ/BgThlPB41gnSbip8xt2ArISwI1luKllHjeGrNAC
QNLuqdEhGzUqXORxUrS11CcXDYMuf8Iy0Rpm1vcXHIDikXCHXVxck6i8naGh2t/m
CX4A1kJBjLzfeYWF15ml7LA9HNvgu04KpO8TKs7Ghz179pSVSMAqXlCZJO+ZvuGP
7lOukfU08AwbOSXByM5MAIF809U6yLFdBFOZDZOSUv6KFC8ho+nmRlioI7SD8eEq
fW4lYTzAFf1A6ftOCyibED0nHJERpiq8tICEbGpBnj8a7PVQJp6Ibn1jAtcT0+Nw
CKFUVA1MlZzRRWuXZqABSiBJNE8+ujiy6HGc9yta24EplLq/LivJcgi69dt94Wdb
Pmu1Q43G6J7yShsHzb/47dcmMlYOeY6ZENp3RVFbDaCf0PeurWAOcplvGCkwP+XN
inYqkWYIZe+ZTjK4/2ocAYRw/c4MBnd2bpG48kEQhGgpYyaSCZpSaaAOJnHEGXcb
BwfH+0AGD0iSytGWnayldCUCxg1WzRBYBclGkmT2eYPIqCoN7xGgMhTInWu5e4NI
5xIJJsCb5M0gn0BYzxv7g/UaDGUURWUM9GmsTcA8FtPb1rEmPtAdnyhlTHWdm0Mr
hsvwU7XKoiYrDCwHuBGvoS61UidJ1mHfu7FzJ+fIaVbBovwmztNCxGjm0DIfND9t
iDIsUWcCdhVREuT/Pd3k5hhO09YjAjVBpSkQXbvMY7m8gBqFl9voXl8DU9UaufjE
fOLCraUgkd5RkvF4GytddS7vs8gRghrg9FnVUW2UpLS9aKfTVdO7KSaCG8OpRTiT
EwG7u1fHZc5ixK/57JXGQTOX+b6S3SWZD5XgueFWLAYktiC1k5UrXw6tSjF4b3FJ
L3vLsbbOSGKEhYEA/x8ocNBVY3OexpdlFfPQxtLS+zG23z1s5iW04DQNKfd8kBMb
Fe13AHY8tRrHiSu0emCwcrVG2PzbtknYvGf4o9jwLyjtNpKXwyRkHO/Vr4joRE+L
Q3sJBSMKrrcThZ1/KV+ygBwFLjTVxu0LmpQgicuGkuLgOXJjIcvip4IodGlYVZZe
5GpvABxnBEBFcy2lrbaBraBf53eBZLiJx+/9LV1QuoHon+p26gdNAeHNXW2PHru0
CmNxRAJlE/AxN88+qNXVT9J4hXW0SBNXJVcfy/5VXiCpS6O7OzdaN6ljN+mMX5ww
ViIQSXR/F8pY7Te4NUNuwkqhhro0CIke4qbAMDKVVs3wc0djdkkCCQaAKYRj1yah
Nw2FrpSkaNtDcqxkeqqvDxQhoFJJfxQ68lufilG3MfvmePABHwJZhd1JxILJ6dH0
qtGwjXLoLzjpXuSYDn1EujMeXQvdhnDSUMFAeetkdHZQajm+K8Hetum4VIR7cI+t
P3x4GpibVqxVa+vB4D+NAQT60K98y6TnX61tZfWdQ/JdzglELrzgbE/uW9irE2Uc
ZA+K9VCFuN1Zv8Jf80/XLs+9hdSXGRHDX1WfRop9EbFmuAYPhU/Z+KAXpIxkzPKN
3KL3jrImGrE8uvH8TnWzDey9BeoYLAaaoMC8mNG21axeZ1d5TNCNO0ZTeNda4uXs
alrFcn1vswq+pfniRTYTyVhLWpTR5KfyyYlaBAWw7yrJPUdE09Ko0Pip7/IMo6hO
jBiWl7W0zxqeDJzo46CGVaDiH9AM6jg8x+VVSWy/Ce+q4VdvS09i18QTu5K8naSa
D98C8WQXK/+me06152qYt0bLJ6OOLS/51/1sXJoqMZIfagPk+CAF5moZki7EB4/t
F7Vpv2Klg7a9IxU8GaGOP9i7XBZZL5g2d2F+e+VfRK/sBgPjVPC7yPMAADwj4ujV
Y1Mb58ridyJXHyThFAbILfats3v1ZkBQxmpc3BytMEZOD9sUR+/ZK4N7yYycMfYL
gUn2QxzMlmqV7Sv6ltGs/C3+3UZkAI3jvb2tmsYszHJCXE3lBOyo51QERSgNxRpQ
lz6EDnm7+V3srTzkOjxNIsnM+3KMKlVqvcmWHq3rlOLVeZHF52hWxnBhHDqxj8Kz
+h0vDCGuxt5ejBYkrd+Y0M4AT9XSl2wz2F6BDO92LOQx35HtvSRmGvggWNSvGxST
U5h68WadZOz9ePudgu+Xf7kc+mIxwacwjn1pfrDpXsT6+bDsRSW7LV7MCL8kcSlp
CvhdhczelW6nmNSqnXe/+db3pxu5fkTXYZodSnU7O8BxGUSPQYgAycgn+5pBdXzB
ClJ7nosmNwOG5PSjImh8FJP4SfAMVlRBNl2sG+Egk1OLfSNEsDp64XrOk3ufwth2
eYM7HJP5IfYd5uD2T5binozwAp2i1uN6ltZ/MeLgUFRwREU1vH/dNqYoKUh7ITcS
BQxUCNbohb5L9HYZg0Gu+3EMsNIfcIY0VuylfzbNJdKmuPq71veuJkD4zJgMdr8M
eMkTY7mAJw7KIWoPeNjoW2wArBV0xhRZ7bLq0yM7h+YerU/4BbEQfVJ9BX3PBUGn
NpEKMvoSYOOZuVu9gMmTvFlLrTRQNXoRuAnsFhfgu6Du84n+2USHV0VG14twCnca
+M4np3c9xQ60GTdfNhOtp3meV6ob9adgKt4Q6FlWfnJIqq623QaK7aH9whiSAO/a
fElsVtA8brsk4sr6wPk3w0jcJY4BdY5U5m6dySp2KkLxpzcxQHtcVji8z+Xex/m0
Iwfh5QAxIu7F7wCNcKcVUcsJ2jQRkFrlIGaqZf6pM8O73rnRn1hYXGXNydBnfrJH
68sK/pCB1Q34V1oxacjU9gxPhp4lGLBnpZlSQvGAsktyZqS878Gy7poHo7SYZm/c
BS6Q5L2SSaSP/S6qANYG9/pGItM6gW7uFKbNJ3U4OBJ08S1Ckxw/OJvmZTDqT6jK
OedLz3pQ20FTvCGxkCZ3RF0vbb/ZiluoVgPt7nyM93HjKOBU3ea/w59uMQ0sFRVA
rrt8c9lAGsHUI+gwDbIEfFVoYnPiplanPL2uYIDm32gPv0Q2zayER+DFBcPtC+mA
KTK47gJS3GOo6e2iZ6nlqH4csepWQ5CpbLqzyickFrvRl8zmWCRF8uYRT8JhAPaB
5jE1QzRWxTdCrt+w6je3cv/52ZCnT+bX6w/ORC1aqyWbx3SAmzKEerEqWmo08tUn
FUliM0gwNLhflvZM+tkf02kdED94YjjL+1zJeAq0CxUcwGTPv551gQ8FTc8X5Fp8
Gv0vY/UBlk8+LRxS8w2AqQB6eNnn4HjTJhrdOEn2rzxiUYx8kvoDCHrsWM14k4uN
pXCgvGH9PKU+ku8RnFG0H9rrYHeX4HCgBK4bXZ6WObk4484BNZ9lHc4T8ok3Ak3e
4iqNX9x1eS/yaA3gYRUn7GgGLMFmOUE416CN7CjjXfmXNvmXAc/5hUCNvTIZ+sNZ
mrTQFnReb2GyRrk5NK4TFZ+Rs0rLIQ0VG0FmDVAbfUKRfl/CGBZ27bZJGLQGulsO
1fxeLsKSHoJ5eubkW0cZEV7XahrEbPZmlM5mnZxMWJxJduSX6AuXUaaOQ/GNrNlW
aQ+dCyWUy/KXErk53mcrVrlb52LgGGggqa6g/BlwUlK3iRefDJnqROh3JXpMfI0Z
U0Yn/8tbhFTuX0iFgLPFRMx0xpsFfRdJNgFyFi87BQGyrebqB73PC49/wuVE7JEe
UtUUxnHyTmJBo+s4Izfq4tBUX+pVa+C3sMXDBtPYjxpPFMZBJCZMX97Mu8NcQTnS
6wxc5ViGV+ZmAs1YExrGdv6htqo/SQjsjMjBdvLEOmkCiAzrmi210Qm5fyigUrCT
E88y7mdutDBCtI5+6k2YevFxL/zeEqOORKruNVoJL8FZRpnzHXJYptPEiPj1JsK8
QnlWUkQw4CXL6rW02R47T/ED0eFW6wucMlL/Y+zCy5l3UoRXbgRJS4fVeuajlgp5
S9HhEbiqpJ68DR6iniAx1BaYNQveLSzkMnU5NYEGy+IGqxzwDTsSKIN5w3s5lku5
g1XPIhSPeS+BGf8ZrXo5M5+3jmn3wnfHHTDw7zQMM48iUDJycamAXf9v+Ms9PDVq
S0aJ4JbKU8KBGdTwL42j92jhiFCNBD3bw7gIHtKBLF4bGciNSzI/aEnCvBLrcLVt
Mo2U5x8mjBO6woG4wDCQ3ARXBmzA05F3v8De590evDb3ph9HvRs2/OIWQ7dinI6R
9VgDhYhT2uu9bFCLvroqpm/Lhd23kv5bGyFdnjlYyBP7aH6UPUMvuZdVgBk0n8XL
AF2d3849byZVpTtqtQSHz4/aFWAnLPqpS2g9UL5hyzykvyu9y5A3NCGr9qL2laoM
080HUQbJhT5LyMJ28svLc3WxiztGp4hVKxkB+aah8KMqhtys88WgMQbcjC0rBaW9
QVjJqtxTyWqcogIvGmNSYwS+sh5SKGWOZAHRruWi+4oTcMZ5KpPKQYy32j7t5DNi
bfSm5vG+xRFCR7T3FAXwIUfqaZgsxUsdt5Y1A52ZrO9D2+q8xJsg257dHyZaM5X7
Qan3asMhGGau+OybOtsbXTWB1KAJGHp1lCeqUch7ljxDBbYkzr++RbGgFXXMgqQs
IgkKmFdj5HfI5P+QQ+5+kYxhgkQigfIlYgsGGL/KQv9DQUjlNbx+XF0XYgwnDq+D
yRvuAbqFJJKIvbwuTn2NAYsxvYtEeIi4a3Uk3ViikyzKgtprDYOnLeTu6ld02a17
32sASK7MYrregYjSopfHeJxz705U0AOocTXFJUagTfz4hBzixEs1ldRcAAHuezPH
ygLlMttMh/epTDQCvEXiG+Ykx05EFKBLCqoi8VWfnDoehPinK7yrGxmZnZLuIWZF
gBg3ihlcfQvC5330kKPck0KeF3HDYHeapsh9fV1iNj4rk+eVA6GlDOQPrYwMksHl
OfP2N4TK10/P+wis4D5imuD9It+cVsFCBsmTZCbXUVRMXT4HU4c2hHXQK1wRSl6P
utC/2Ad+cyw/wu/RU4Qh7t2ouCw5KurY+XP8d/B/tBZaRErN0xSQrwAxjiEPhUEN
Zgoq+vPuk1Lj9R5bBMHDeiGrJf78WhrWVoRZWm/mBXojpRycTP+9wNz2Ti+85aGg
nXHGHK5y2Fds8+1zwi0WIvEsgmdcN6fdTN5F25mbvCD4D2nVe+UR08/zk62YllYV
QGnFA88Z5bmADGGwXwv25rFwaYyE+B3W4nmlQ7EAyC/FZd9N1sA+TZUvdjGfu73F
F4WKAwx8eGOrMVkUwVrjK2Nk/YHsB+N9v9r4XRaqFZPs8806GDOQbGzHGwvCb3Ue
YFg+4caJ2xN0PmlAXPoyj/DiZtTNujZxmfuiYlaUgAIyLByOEYXgDe7x5m1EnlBs
gerrGcA4DY4pW+FIRspmXqBGLoj2pzElKoq3DgtOPNscfSmw8S7jtUQWYnTmeU9u
+Kwyqbp/ldcdalOQKsBFtCrdIzeJXhpfxripIedkuNU/pJ1DRv1THDGgN5VkaUob
dwf36ijhaajLH8bdBb0bbgBGt3Dht0zrMI0ajsyUZotwCAyPWTUMJ4xN2aVsS5zs
rJPw7L8n1SsE37thQTc1l/vlEu+ZRsoQEtP9EB1LcEvdC0YIdX3XzEA46XMaDzpQ
ouoMdnFhXQkZSH0jve6WNB7sF2Ci9lau5BgSymsoTt6GcMEa85kXMFgE0qgGnwx+
VjA9JhxbjF+MLeXWJPWtXWG8GTxV6D2FU3nlwkVpmJJSdA83ydswZ21AL6rZtkZX
XJq2QYGo3SKotMw33/1rrFo8ciF34zuiN1qZTZaefZi/sPU/xdKyL3HZl36XDwfu
G5Uk5djT4ejCuzGH/paoG4fmDlSPu4MIuM/joQn5rQ1JPi1E73GNWj89FJfLv0YO
vA2uvIIVZMbHbanAxQIJ/tOjJsyPBOlThSmdJkpLHiI8uyE8cYs5awbi59Zv2jVd
2vza2XAKQ3ywJjfWdi3bWUEJV/NjC4kv2RssmoTAWrm30R0RmKwzSHVKWF2NrDx1
X6W7yAWNaIbpuKa9rBEq4WM+JdKYQIQo7ZvqTHDiLmAwHjzpQBIUq20OaxbalgdF
qXR5+fbFZlrYeHwlOkQiVPJRT5I/ssD39bxRoMItSjOH5VeivUSKgutIEOmF97E8
etCYGaLVoEhJU62cIkblO8TjGVO40gNERs8lUHPELQbaN7JXzy2EjoAxGGGLZzgb
vALF9xKZ7f9Q4VWs+TTvZhzpMgDFJg5R7B/VD4LNnYYqJmDRH8hlJBLzDpXWyv8o
tpCu5YXoYCNhgus1pKX/YTNWrpS793fgtGHf0cYr/Q3qpWgJ8I1MBPbyR0x7Cy63
d9xwYGh9eLPGWTw8D09ryX0/7N1ifPAxLF37igONZ/Pu6WAuUisyIJ0niYvo8y98
DFdMs5WWXvLuOeIe6qLpzlJyg5IzFt9H60FrviqJ6dp5F1EgxlTNeuIFjTTix2WP
LZlUiEIGY+pYNcFzwDVSm+kEKiy7656c2jHec5AJb3KW87rSFGxIVY+vPfpfmJBC
wE+gRkUZUXfds3KgdlETrfxJFk50qezb2F7mIGML+LfK5eTPMcgXs61FhfXPTNEu
0fUlBGXXdeQQuo8F41mJxxpV81f1jE4KHNw1WKjRwej5SgEtMM6N+a1a26Ra1jDQ
y3Jdc+x53sxyWu10xbM8x3jM1AIvB1VerIkdkBumDPZVynfpYFw2MKPF+nq1pSK0
G108cBkBpL83qNDP+KhRRWm33j5/YVflcbFAwQmcVvXQB5+EcZVVARaCpkIgfH5q
5mJoEtL5NGr8LcTmBJee/S9CR8+Mwpeq+h+btp0S39q5b+3OFZ3StEIhZ++GN3ej
WkZBEAgPoLP+JxNTAeABbDoYVdKRsFxhUVL3VRKJfLNKtV1/2iULt48jkSRmijXl
vXICxX0+FOquLCiZRfFfW1MuxJc6P4etmtcJ7A/QhBJvGzYTpsQrO/L8IFFJnNbs
okmk276DAwlGRqC1YKNvVCccSZM3kGBcoB4zKzqVWA10UtvTMCU+1NVQNKiNnb6H
AbgD7RnzCzTgx6kAzM3IWZcSU8INDqv2gXMZ9vWrDGrK/KtoBJlSnEWcg2HbGfJ9
v+ZQYjlho/Qtgh8Pk8LX7UrkanZ70o0u1z1lMy02Nc2jHZ6aaBB28YRKBjNhE+mi
1bhU1aWkbMES4FvJpnijlnptL6sbaWb+HJPDi7tZzouwfSypgmVQLEEkUhpmLSsZ
6yb81xbx6B2wghKIKToK+daczwEtc+iUV7VL7GWusMzb7ak2ieWEIfjV8vxYan60
LylJ6fM0hI9FD5ixTQfXNVqGRXDrS8WzRvI1baWLdE/rFEG3khQmLYlpoMMBUkmk
qPOyYl005ZDuchu6CytA3CoQQjpWGpBpk5NbJAQyxUp8Pz74lrDF47F/QJZHMXAn
Ysl6EO0fP1twzzUIoxPO3IaOPc/62AaqFQLYEXhkMPwNHP7EzXRD9b+9YvXMmUn+
caSFvn+/fJCVcp5DpV4Vse9nu8HuRrkF0OtcUcxJWfnV/JOvhm3x7dQvFVlJaCw4
CqAPW3UqwymLnx3Yw9GRfWAZFeFL6AZBTUDuspzpzQfWgoswWH68IdFemCdYKAu7
xHMcEP3NJ4tvAnp9CbpyuRB9GrtydqOi7llsHft6LSMKyCIr2bUgf3SyKZxD8Lt5
7TgaoGq1Fful8S/qOKyhoMl2xwwSY3D3lBQEMXQps85tXWvOUKscs4DyqTTAWwJl
xHk5doAMkxUE/0zO4wbnlSLLc8x5+e/oK7OEZyi4RtqeVji7RVqLQUr05FZ2xGyd
erCdoomcCIs9q0n4ykTLkZykDDD0HzTMf8FQgx7JoJ2XsC9+SdK2IwQ+Dn3HDUlM
kcaA+gOfazG+9YWO/LwZ8Mt9jTwlVA+0vlEu3B5n/uVYFVb2TwM2U7lQYJ77Rxgs
5hRvvMrEm91vD/dzguPsnBVEo0voBlf+Hdta/AEYJ5lZRlP1S2Vrmm5HmFUVIPlE
QGKraLg9tamYoFkjMorV/087VztxjhGpSaxhqYh5hbtqmrelOFynXj4nwJthpkrN
Uil+ojwL6GSXEHy9r5gaafXYAZaDaSWGdrv+otKLCnOtVlfikAACPm/9l3qaQehd
/4qxq4HUYr1p7kyu6U4HY0oDiRF+ZBQASYn0Or+AMAIL/JkTkJG93BaO4CimsTOX
FrvA6DqRfoLFaAzSYWA7Y8YGYzPBipI2vZQFYvEU4uQoh4UBDDA+L+KGlDCW7hXZ
LkVmd9PHf328WIS78KZcb9mZ0oxwDpPke5308eb+EU7zx6+deoF0KX3zHB1JbucC
s0AwbNJTg30LLTMVOb5zOE3AiPtNdmBM9vKefIJg4tRyUO7ZxkSGXTfsCVyTDa5Z
L1IHxTU3jzAlUKMvAqiWKGR4/9Y49oUD38Eua4FCwSe9ONULXnG9ISw1LcxA8L+c
xAmnQiEA25EaTJKyX1Ac2BM3Qz4YCpys8gudwNRgDJrZpyZc39sWJJBOZ3zbXZCJ
zO1OizkY9CYUZeLnkEFAm8ZVadF5EoCvesis3hnJflJmLYWNd+7TNHpjH/K0PE0G
9Ylrfl9lBVWMXKgXb7PrqeUjrLAz7k0zjdX8nof35CsuzGONiiz0+p+YUtEwMpNT
sLuwEhgvZS0HiMP6IhhksIjRESNjwqFuE7W/Y3emLhy8qHCCZOBj61SMAka87vmh
be2YzI7SMLaJC3QdnToOyR9wEBe5wEvrPYWvhhGOKRCm7O0sG8PHJ3mF1e8CgzV2
T0xkZzR4ts+wwH7FDtxHpK66lYknk3PE2RpXcIM14CHA/wyePiegiddiFUiB9PyS
7QKTWek4WFPt7fId5FR5SAOVhPRPWpFBcTdvsLvDRXPeLsp096M71EW3e3utVrod
j8Rln7b/wNpB3PuGMtYFLEMKPSi1uAC3J5WhKd4YXACsaK4+T/XQdrpBCytp3tse
6i3jqt4szr1l2jHjnayhpoERKlrOn0PwGVH+9MZc8r9kvhgOEDqcxQhQuUQEIPuR
5+/Eo8ekOSfD3rucM8PJeF5me8Uqb3opOFARuQAwtkFgWh7Ku38ZEFi8lre7OCF2
E/d57MfCHO2cZYP19Ar9sg4XfX/Gf/xlMr+Th7L057n0pWcT9Wgyf16qkXlhCa4N
6gsHyp02CtLflDLguy8x1rhqfo8udECpgmgZjceme/EF2IfJ2LuEnrrBOxCl3lxt
3FIO4+Aco0GdXDEquxxbABvLMnfNSqwiSjkQfpJBppDGWFyRtTRVXp9JDODgsgbW
yw16+lF+/VYm/GcYZjlHUZym2xlffRSBwv3/Fyx+Z2SCMJs/7q/8fHMR3RmutA/I
5Bfvr3Xt1qIbnXSj9n1m8aEuYA3MA5bBb950bp6B9sbmQ1zovuOYKPp/+CCr7E3H
NgdyAfXaRRHTewjAP+oRCt/a3evCb8axY8aU8kq0OinYdQZI1xsk4bz9cqLPi57x
OehsJ3FTaHOT3Uw8QSLL7lHTx37towV4uGnayOXrSWhjLvDQmC3qghtSErsa9AHU
VqjiU+beUvjRpdqZwTLoQOifW8irPNbtnCCxLNnGlmoDm2/GmpyNPs9TbQHwylKE
VULahcV9w1tdsEU3AKVW3NigIQdUgWpgXC2/a0vNBmwhNHYk1cCaofx4T1bPZEDW
kWfxoalmUskCa6IXjsP3i5oDx58Kw22B4F6AqPr75WclqlRdIl77dZwde4O2ZejN
C3BcJa1yS4qpx50yY5T8QzMdTO8WJdlENSgpBmyw6nnv5wdKfC/MBOUuCBVpsWj5
SYmi8r4Jrg4ofFb6YBoq+osFuF8BsZy2oNTyzmI/arZsSkOaLoH2eo4Al0puqNna
u5uuCQGqOPG+sqgWp6iGv1k2RyHlpZNC3gZH/HJ9ZToIj37wIamta0JbONPTWXyq
FbV2FdfwsPBbzlxeva+ysjHI2BGYO8+YIUkfia1AWGgwV2A6voO8kOlda64joZqJ
b3j8DmYUhOgdb/wrL5qUQgo0K3yyjko9UWMGwMvjDbCLhTT8RoC3eoymjCaiWU5g
LO2zmeWWSP6+HtrUcIO0btjTRfCM/PG0e+tWXE9uCgLkAmdkY2GyWBlVOOA8v/kO
nbqoxvATlaKqGuvuqgbT90RlMG91pOBetZtL2/6CGfyx8wz6ikmhZsBQETmi3NdJ
rT3oRXpdBJBvxOKFxgd9AqmKHu9D8p+aNu2xSkKydpWWsoxspLvfC6EYVOZVt1cp
uDTpG6FeAwt+9kgrr04wwCAfIx1nvrrm9yLbHiWQ4j7EOgysxU3iRoejz6HUxcaB
koSgpZgkDDxaMIxxEqu9q0L6cNpFd3Osk+YqS6Ge1iuDHojWUKNaJ4rckOLwUWGf
xB1LolBQu/GyzmyulRzgcaKOpuDgOAb7bOJGv1lrwsnnYAlD52PGDLCYWhPLAiw5
8hzpSU53mcscvYc2I0EI00pviOX/5XVKWZqPCJXqTFprbLoy3nUUzReomjjN3/jL
lxePWV/PPuoYV5k+Aaek+zkwIvEoOTcnC7R82atBtrMlglUsNlX+8IqLSeQi1/M7
ar84Sl18z/p4Wz4v5utpYXKQjjOjjivbE7K5UEhMJPRQ9LI7omttdDzkYFUGDT2i
VxNo9yHS3f4JLIwkTH2sdJH19DecBp1s3ibkDpRBvu4qoPq1LS4NUykkhfLFW/th
2gd70CXSCVh4ljoTlqJ2NeC5o18tnMLP+oc9tHfrfFr2+bjA25QoznZnVeQIT/3A
WxxKc9VmE3uDGagadVg7cX+zmoR7K0sRMQUu4f12ctzFtOieCUgZ+S99CR2FK4Ht
QagZaNsnrSCmLmgTldmPfMSE/e+D3BRNUYZOtCDCMIdSRUuBV93/yTCg7s4cz9Hs
bNHpFJi4kBt1xxUhVGuDOygIutmPngIdYqOwheOmVr+Nn0Ke5qenpSWwZ1em0SVn
SVEgjzUiXkgbjXBKVYT1NbZXP8Vm/ttCMknpA0p9LNT+aXcu50IP5jHl8i5jiASI
i1jNVMShW/1/OiiYw5uGl/lrpBOWoiJHtJ1HqX+BUv/r6+AN8hrZXG1oHdfuRVYk
NGdOgg00TyWrgPxRnPHeeFTIqPOa/sG68NDr2+1b/5DB2oEokqihoolF2xSP1SIU
fq+RBv/JLblm7NN8xXTqxXf8g4enoOIXEnBke0pEpfxCevHID9J82iRozYd60O9J
ir3tEPTylNuPBdQDMHMRwXxCBjiCGfEo2X2vH7Bfn8LbtpD5YG4Oq5frx9Nh78a5
6kjqdZ0w+YubJ8z6tnxZ/iEbz2gjNr7doXzV1pffl4Xm0rh6ItkVJ9KWhTIwQZMe
ErAd9RZ7uf+8f8iFf416SQR736vXL/Zd3/j3Bl9X0zTBA6f26AaPbloiw7TcAD+E
z2JLTkh2hEGpYmpHl97Qz56JhlPR9hkCCDMc542eSOb7d3ImOVKIfb0pHr5HPO/T
FDTcBZ8oP+J1RayodRePpg/xmbdRGntFfk4OmmcIZ9G+4u799UErebeObSD4bJ4m
dyO2ftGAeL03c1y7EIXdXmxp9dNnMyWeQVRlhX/LJnPrmAXPFpdHFbwKaGUrt22d
jixdt/CmANsGConQRR0mZBJG61J7YrxaeC1hQWXrARzm2Tpto1KB5gESAgtcWSPK
xhCetn9pxH5l653kLXLvSPyBudnZ+f8wvKmDrCSAAy6E7siKvhzMfO6iDGk+RUwx
pDzwt1nMrBUWI3/zAygmGVfrTUEJarRGTNWBHEfyYIoCqWTApn/7/HsAnb2j+/uI
On7/HGzTrI0PSciS3lmBlr5x27OcjMiPms1c0PsM16vdAhw8BIuo6v9LYMQmUTiO
gTfIFIo6Lgl6y6mRzEYvNot8i7davR87nfYyu2jFtkCHenhqRkpo+TIhvtJLD5ww
eu9CGh06ODNa2CsWYZcW1ezToktGxTXO5OJreBX8zKrpRjgoOzZY7bI6gIpHySXe
OR1CmFzrUBwnLmpk8dB+Fus/rZws26KH5vzenglW2rqOCjPcCnX/Irf+LsOSbC61
oF+vx2A2Ora5d+McK6rV8YKDXxFLFeWMcxgI+bXqzLGMirv2PJe6OejOIAhRLrZE
LsLNeE+p+ySu1Sitrnm+4TbjPsuPpHnj7yUAKHDq42CvIDu9Af7v06TQYC9F7DuS
vJuhN7qO+OqGbqufHLXqh6ccfpsWjd4edr28p6wwiM9TpYc+ySNuAey1sZoKBj5C
uW6XjfEalpSuvKuc8a6JUE8K+BGhKSs8SH/FOicUeftn6SaIC0+xwOzdKLCrdMsg
4w+c6tWXpEwZiTCBbwfGTpujbJjPLP0p295KFldYlB0nQsh8Ezm7ZUpwUdSoC7Gu
xeianOdd1k/QL6hAG80hMM+O1YJikbS3+tNa/BLUv/G8OVL9ouebJ0QNtyf6FGWs
YRuRMXqCgxjXrv4a0E7P5PDEbz4AcVIDaRTJLnaej2uOhLx+Sse6EDPE5ydfwUJk
tIBnjM6P0sU3DjWO0XDwEZcZsxg7FmmuiIiSBuwmrjSjhrx4dZ5PbfCAAEUEiwHJ
QxAm+2UOcVDy8UPk9vKSQ3FkinjYTzoWWi2QG+3AN17vTQU1YabK5eP19s3Vi4/f
xTh+L9cbln31NpRSInLevW3jwVvORMP71dRfFHeZ6tE+mGuQA7aWnHLiHf+5dKJy
R6uDL9SyF2uKo8OfUNJNR/NoZ7MONZRAxxdYMHvJzuUweXVbKj56y+tWPtcJBmI7
in+z75pOYlpwOAct6jW5glk7Re4WWrfA/4ZxnUdacJRWMgjGrJQYlN2u9BAFTRrP
l3d87Nsrm2/dmgEcxj9KXOvkAWBs5WCyfoQvgn9IFeB9t966GbSb1mxpsODX2EUJ
MvHjgXsV2AuPfyPHOWV5hRhL+uPXgmd3968eAz/0LVFdXwUJwfln+cK1bu/vZGZ1
H1P6aZHgp/JfdYhRZ4zXS3hFv8DIWoH/J5rhVi1IKwizfMssaWtqgQDue9gbItud
Drjk88pXuuyIaGzRGhFxcumHW0ScZdC8Aa2luVyiv4TYSxttjZVIl26OaGtA2Yy7
zO//350ROjCTLKOvo8wMPaMRsymE8VkgC2HKCFtErN5fx+lwVvbSJLcqfI4jMf2b
NCuOZljLeC5gvigplQ23pDtHKQQTPsPeVVmErkvgtZDZhpbCwWL0IuRWwW8g7cTk
0nsEB0AplPl+Zra4TF8tMJsLBsL1K20gTdE8JWqG0d0z/Cb1bTvGcu4WRw0iHSX8
hR5g17E1BfNoSLE5atnkyNqylOPjbfjpVds0c/DJkcqfp9F22f9a/V0+aHmmpfBL
hvtEoY8Zym4JMWEwY0bVSU6+EPjO2EpwSCLNPw10z9oe1N2dGnP335PjDGa3ROdo
F0zP7kOplLwKGfoRMa/0NRdHzCPUTgGRLl0Nl6+TXmoPpp4+lEVIKZKD6DUfykcb
QcRiST3+MIylaBoszSSprZ04mZC3qsQLekt3Vo5T10S+tyW+nSAKbZLXOjQH/6TV
McmS56kAmdLox7D+r1FXlO7jsRPApZPBllyGPCXgV4Zi3FRk3I6eAYGXJSRIgAh6
UUpxsc81K5xtLR6Y3jNSSow1nCbPtFi+0U5x1Vx8GwakrCZJXEfaxtQ9aB5eh57R
ichEg5mfi4RBq4cJBX4mKcU0Wquy1i/oVV35aL/X/0AFRFzjsS/r4gXhcm27cAyF
4tF6DmbTuBiCDvVa1QjLXRhmkOvtw+BwYdE7qwd8I4LzqOu9cjPwpH0WjcntRi+M
LLU5alkmJnFFD7lAeRZcEOjy4u8BfHj6f1UdN8/dUK1TrPjB28pa3m9uPJ5K1Xag
gh0Vdx4E5K+yKs/MSe3+G2PXqgtAO4NgbZSKiwhWuuP4ScLMTSJSLq8JEXc+wHWt
ENLHuDbhhoxGy+zN+WB5WS4lwhLmSlXt9D3S878aeyYnUBOlPU+D8VJxFoUq15EO
QLsdJHD8r9p8hZHgN/sEYqc3cTDPLBJR5O2Nb2ER5QOKOwxVevzdeK0Llio+szRU
GRfrDLzw1NNTJl3XByxEjx71xTLjg3mg951PoTaCFdg9AzO8zWq+jnSWLmd4V+Fy
5u6wem40TNHgmVUC3Kxt65yH8hmxOUAsG+XGIL2n0z5yRojrn61HEVilkUqnHxcK
p2uiQAOcFvVe5tOr12lGYbg2g3dS18NOvG1+NmmkgUyOx8wl3RDCUJZp4F0sJ+bj
uElGaxT0yV1aDehf8EDoo13ZtqQBdj/ZnBuVLEGfVG6ELiEsco0if0mZtffaCXog
BEohXMM0EdqIsFTus4uSYQr2hYaYQvVtwU9U16zf2S1Rmmo7lRwMvtkEbDdqp0w7
ftgll0o8c4ZjXk15jP6noGLosHn7S8l534LJ57et2tmBYEDrXXG9JCtfnzYAZ05D
5c+R6JdpnzGB3HJ8OQ4gePAC3NI/TufhjfIvRctam0U1ueZ951nsCJr00ZxAX8Ne
D8NSx7B2+mW7F4ChOs4JMbrdnxvSal4zBO03XAd/3faA4B6DUqkzR0E2wMWIuUyZ
ExVAN8vvS5rHFTUo7TN9qb5PUAj9CknXIJyhIWBxc4UW6EQ7tTmbXzamU4X3xT41
Dv2z20m/c7ebDdSqQ+yAf/UN/oQyTSATpA5AW3UKf423XXL33hWbYTT4ggpA3kSE
FNp+6W5uYXOrLhHLLtSh3pI9H6hXQ6mSrC77/oy3qrbolp+4jh8UhTGegCmjmZxk
yfMKrEU0JmfDnBn7rycyde0JekoYvG11LudFuK7Z8Mu5a4NswCDp2abh1GFaBvti
90vg+hAz49rB9Rau7a5R58Y4eVrhaWG9GlzGOgAeNRhoMxcrKcuUVbtdD7O9xeoH
dzbaEuu+jnxGX7o6XBeM/6+mqTKp4GFooQf4g66KTCoWLZBdkbzlxvpasd2eFC8E
Sz3xqBB3ypSYquJQFrbdY6byiiz6tTEsnY2vOVHQXzOImw0749ur2F77OXgZnpil
6DurzUXXmUBZQo0pVpPUhAzOErvq37/+pUlERrvf0QxcS7cM/647nU1AEWs5fOba
YsN4m4wwBIZB5OD+k1D7gZ3t3ZrltFu/YRTcyE9mLe5BEo95F8FK8WZ/BMKGIUJP
TcbC3Bucqeid/VWtFuBc3cJ09is4GkVJJeC+xx7Ij2+id8CqXtFtfqKV5n+7GSDu
aR/25HBtFynR4H9K/dMtTVMqGoIuP5hnNwGUnYkMpWbJ0HeWlsKRobKSSwrsg2gL
l4tcjIXLybgpnCJJnt8uiY303hpt14FD06UrQ5PPZRzXkcb2PmjwVw5fUY5clmIi
K4SPKRlLmu9/xBodyxohSLg4OZr6MkV9bg+kz8rwK4q0mxswJutesfAqmY/V9QP1
EQzeMQrNbIeYE0SxRZdZiV/2q2s3E1M4YjfTZchch0WhB6O5VNMPpDPxsdF6qpsW
6FZm0U1OfH0kN3TDaTpLJlRH2iD1ibhDJSgfwiX+zoJGUWU84cyFGJniPVFvWY68
4ZbRX/xKXNxbSkEkuDmz7+j09AMvFwnseM6vcnSto+rkVwReS3fmgLBRy204ZxRK
xVweICJiD1ld7kZ6aBO6lFDVCvCtFWINMmqTzQUxNSHSpIcSEZjBihjd+URrBfqg
zxacjCM3VO3RVoMJBCAtPUN5oqJuQpQPr+maQsZxgiyr/rTyNhxpKKjwq6SZNRl/
+nthCHDs9ViS6NDZNUHUVfG2qRgSiSY8C5jdyJOeuE0avbsRpK1yDxK/xnoKT6Gr
DYqijRPOO/XFoDq+N4G0r59rLAYbmjKOYZ2+lmLYjjL4yVGMxkV/aoK6g7jjKGSh
XjL2DyIjvBsJ1uYc15ORMOwCdTXcLf6IjSAoTW6zFSphxMXjBP/JD5BtPyA+bjlA
R8Hyi/r+ssieLc1pSf7XT2L6Qk/VSXZzwuKPlpgrp25N9gsmMdMVdPJ3KWTXXS20
/4v9MjHmRv/De34WVXwg1kVvFrmdeOywfG2zKCKQHJCPGJKoa8snUcZlRqSsJQLZ
HzpjWW+JJPZlUs1Q2q/vXjqnOq5fcHIGykOqoXMiZ2y6uEgzkfJ8YcFML/gMKPgI
WLviIzba3QoxI3lk3prRMWD9zbwbof4nKkL9UiOUHJRE3+jD+BwlmrTWYN5akhc/
vidtAE5ZJpazrMR9zL3HS9bUBrwXe+ofFMr/dsM+FvbDGHYFD0MINBs0TV7jLZdS
XiLb9eLjT4OarjiujfxjlAgPjz+MsFLkBR7x+NgLAxDejtz+jJZEUc8/5Tl+b04J
AiAHV7I7a11PoYhvy1+voq45AjL2qZkjS7guZGqUP8Y/2bUYqYueQL2vN5OzrIg3
ro2dC6eaPS/tArSkCMOvkmbTZY+SutOzxpS7adHhwZNt7kHuMiC4LN59j0P2JSxy
HsIQxzMQNvpi3HgJWmySpvjUE0t+GrgQ6HbwSI9Ut4Txr9B1Z0Zd0Kx3/euZTeNp
4JTKJjRgm60twyKNOXxy6TKEsOK6wCRzLb/nAOp8bs868FtoDysqbNziAO9BP7HK
moDIHo5Pv+YqelWF4U2EpBe3KSKwDHkBtvv6Z9rTTzRPaAy36S5HNkqBEgEAwxtP
pyJNJj2m7n2MttOdMbwxq4AZzNI9XOV8f5tkQuamWv8mgKzYg/+DjiLX2eH5//2X
hKnu8fXnNB5z4XYAaOOwOUVwXOURsZbJumYGJ2Pf54yh4cRfYv8vVPQvfj0ZJ/Gx
Siog/JQOLBoa0C2WZfn2z1tJGGX23PtTV86zCMV4nJTQuow13llDD4vU/kD0FHgw
pHpEAsFWpm1GYjb5Pf5waTR2LQuyM+s1MLmAqgy2MfwI4EnxvyN7O7nTWk3ppbS7
H8LkZ/A+e20ZHVPD1Jp2Rpv8eT9bcqZVNbU4dED3BsEyiGP3wglA1P7lVzhvQWCs
aZmwlURG0FbxNvPLrv9VzMZBDG7n+xQ8i5G1HmMDhrJ3D/PvXyiW245Ep8y/tX4+
OYKxzBAeG9B+6tNc9XILMI/EYk/Mxyl5XsoSng+53QCL7nzk615v8RxZUZ1mc8Ea
71AsFr749NAkhzPKT5ctQpWT/NQ+aTJi/2bwA7GjdvLMNSp8BHtZNsOqVAarmK9H
0SdlZTX/RasATIhhCis2wL0ah7cdvZzuUh2BhniZyuU88hxDpXGHa55vJazNcjN8
OO5IqZg+fPW4nuIMY9tjkF2XPlod6hiqx+3xoEh6EdfXwekbLGJB7s/SCM/WfDaP
DfM+OgAuDBVxWZutRlng+eCXHZUIOww1ghGJa81Cjzg1pGKX+1p9cwxl/TiSRuqm
0BHklbSQkgZexPV0sJ/jZ64ynhaSZMxTYOz+uipd/iTcTtZuh+9e241bbKdPTzPn
OIa3kz6lumCcR2ymv7dNxbGN6eQcfDD+oIOySrYe4Den7P6GEfvqwkPFUZ5QOheo
dQ4b/cJFyDcvZNOK/UGnPvEOhu5LIiRPX6ABcbY05K7SBWVqh1faHZuuda0CpfHy
hrAgIgiwpVPsv5Fw4XK/BLPK3KCI+lQ7ZrEm7gW3333EipVQlzBv/as1PZPOb72Y
mN1cLvO434qSYDnn4I0WJfIBLf22zXzLtc5jsLdEM0ZmlEzlYcJ+41Y74N3ocZaX
b+Sl/cKeFyxn2NIwA1GR1rMYWLWtAJjB75HSc0ChngN+QqOA4O3yBgVsmbWu7u9J
zR6shQ5Pqxr6w3zN7qFhW6piD3+sAjJF2CTyD51aVpNMZZcB6cGBigddGeaI2L3Q
CU521Qr2Cx2SrBhWZuXYrJR82jo+uZz05MxlYQFgIOyBROowsP9M/wAWf00u64KQ
7nOpq0enjtDgfAG35ItUbglpkV6g4L7UeEp1mZxm0UwpEm1H9EYWkG2QYX+Bw8U1
1FVN5JM+CCFZB+PPBL5yxmxv9rk6+u81rMPkDisFGaVaESESMLGOhnCCuGg0SPQ6
hnT0Xpf2PUZeNVGWqlkkhQYDh/0semSipJlqQ9KG7cGYnRYViNL1SpKQmVlwKtPs
o5WK+1DrYAbUxOkK5ALY9FKSH0nAynpH7RxM+9hHw/Isp2zW8wEjkVK2OvJTp7D9
5GbijGBK21lA+KOFSWQgTM9sEs6BfG7K7UwWCgNAQp3kY6VNTjLlAFCwB64SQXAj
fOZM2OmIRqXYEHJ3tWq4qT+myYdo6VWMK5eJxcJvpJfeVna6d0qtS9w0oVdOXBjk
lclw/PDmvMN69YGXLN+L1TYQHyfbv3kLwImiIw6ne4w4/lRHl6or0GHq5P1bv0cx
OFNftz8vwEPXVTGkF3f41CFWoSSpGvaV0Rqlr8jRLZ69ndsyFQTTOdI+mFFTppg8
t/hn0nhJGlAKGIHUKO/mDr5Eeno9V/3dXMvnW2d99Tgedgj3wvv5EBacgzl9z4xr
MMRFugOsIKG0KUdbNIHbvu1N2nL7MBqLPS2ws3Mj2qg3WiOGRCD7KKFCwwjAW1bd
AEiJzRLQBhQiMNE9m7iMTuRPAQMrknajZuql7r2Ue3QpHkdrPBXRF2jp2DkBKUf1
ISGlRrpwHKAq2hrG4qvoXS4Gm2Xy5sQXqs3dh+052DkVrPMNVe0HwYpbJPJO+l7i
jV4/p5tWR/c49fIOiKmBj8m2zilVrD5NwhctJuoyaXz+w7gamUu38iVEy/J4Jiac
l5WfuV9W4JNzbRYb793ekVmw7PmYXnLrE942zDOnMfsqrNO4wKY6M4BAGadgGDQ6
0qdfmZ4ERlJ2MRNJukwG0/63wp4mC5QnmlnO+IZgwEm6msuMqN+k5a+87tJo+M6s
oDSRFAEkaqo3267NYuKI0E3TAwSpiKPgj6acMPuGkmlPB7NhYMq3qPeHmWSYW6Ta
//cn3eFxI4TU4SNT7QVehu4A4K6CeWwys6qz+FCLeZ+Hlc2ag6NSswDlHduhKGwU
MTOyn5+NVr9ZHYuvz9bueOF5L3cn7X+YwihYqTWUkc0zQar/fmWWU68OJTK/yzPC
tpmyJ7oXuDkkdqHsqsP1k0yYXrWmu2eGMzdhq+Hx8GHlPSKP1w6hqV1nRWGzKEDB
d8N90v7QS7w3fRZIDEksTlbUk4R/TaQEYdifMBDSyDTf04vTwA4E21IQqpA8IPWJ
yq4WwaPS9J4X8QjVyYkWP+nyo+8kTYkvnlRgC5IGJoWB576v8tT/y/vMKGTHkHk5
KQCjszQmW5vMSzuAL0MRHFGcAi5P6yvLWajJhiFZp/VMeGMyHLje740nNbvntOnt
6wi+tZPwC+mOcHmCVsQhPsq0BhD9iamp7uQIirP9Q9CiW3CLdBWhYjQXjylKxvZ2
N/4sq1I/L49ZFqeIRz8clNPdYjjazE+yZfXZpkfLI7KycGC4iMFCsIAKcf9Cz8T1
T46+cHKjS6LvVASKsUhylf8euC+lWn2Jx04PqXzAKm1tFeKMO8jC7HIeIW4ve3/9
n4Q4vd4fbsFpa7sDxsT8KAjG8d0k/ORbD80hcMK/f4KmUANGdObs+J6+bDcHmEJC
jJjMna5Yh4KaXWGOPvGo01UaM2jNtSq5sFP3wlo1ZJlqljC0TyF1cXqWC4eQ9Gim
3HRL1eBivVIANCEVsV4A/Az+B9AQVhRtAma/GBluqyrFYrs5qfIFy0tC3o6NLZ8f
d35OtrNf2keRQqdOdWLa+RGO6gLqZWi0rCFvJzxBPQHWmBptq4B6LY8x51C/nniR
eEaHqjhJxVgu/w2r2lRwcoN/8Mf/h7vkFGkPNtQvWxYAGtgbLyqszh5JeHRWRH0n
Y8g5ZDBP5yLRliJb93RQavD69mX8Ub8lBB6AgZfmjA1Rk82JMMMp/3VoZRodggJU
LnsoUtYonMauheOVgw3ZHbibg5343Nc6tYtCINklZGNDobcFNVOxd8oqxyx8BO/d
FB8dsaLCX4UnzO12uvP8WhwNGAW1fzkO68rULaavIeNj0G4lv1ubWk2B3MBAo9mX
QblW+F0yTJAYsn4qcYB0XtiryRqzC12RQBpDRXH2koNYp2FP8n77mG/jMy751JtE
GCgLmVaqRVCErY8ZZ8v3kXT8HYEqZ2BHj0a38mjI5n+9Ui27ry2Y339Z/ELefqBa
d8EPypmri53+O4pXyA3v1EvMTqhq1QU28zpS/2yP49wDSjPa7znEKrGh3mzShUzS
xIqGOAhhYLm+g0AV23jNu+66gdKfLGwCfdhlzdfKkOoJtvu7O2ARoeRMFSCDz9fy
7tXw1FJKJwOew1zLatu8/LhUltp8Mh+ZgphStUgPvq2P9bCam36odTzR8SvdssyV
DiPHFmlGn5tGouYzZkaE3ihJum1512yzqsTDmhlpjn9g+gnlNhqOTrZ3q0DxzmlO
xt+Wy6/TsIl/O94IdPJDKfbnR+i0m5/ABVTf/T4fcH1scfPW6DdlpMbXL1VjXRrb
vOLt7egpYVtmev7+BTj34Ntz1RSShZRGonxCa8qnRIgv9KXkLUX/LFLQ4LvDacNL
G4mqPMC4ao5BbdheI3OF5mTtOIdi6vmf6mVveFZ8rC1If0SEhcBEWWY9/1WFaRiF
xI+P+pOhRXAZsd4UlsfDbWvYaJsIBoY9PG9L3RXY7/Dx7cKI1PDeO9xU2zGjhTdm
MoKhuPn/XrBCxo86cs3+kQfU9FQw5BUp6D2sDxnvhXgPFyU0l7AwECcOFr6G6oO7
7hAPq1XC0v74Nnv0gIdiANhWWb74YHE4c+5tB4h/y87gCWqwfKIUIHx1gNsBntcl
XeRFDWZj+yjdbOwRkrzxJxSk/F0cIP1v3NPf5PeM2KR7Pn/D2lozK4SFK5TpvATX
vhmsJNh7dxElgBFpa1Ft8CpTgP6Uzcip/jF0q4ssghU2NTxBXxmqqTMEUv3SfP37
c+UHjrdvOAa5M9CFD5RdHVvm/sFD0JNKdvObcVDSXYjQLSec9nyH5G6GL1I6lFzd
bGM14u99po/DYSyfODtYN/FITN3tEc/t19FT/MQygrUVXNIE71K8zp3GyhdbcX5V
QUM0n8hK+olu2hSzfAftveSheRg0TVEw4LkokwmPmRmXvBiosm/O0Mlu0rHbHHie
/VRXiFiQJ8kr0L5/4BP0M+r2vObjJmR4e4X5Fokqz7Y3fpnaQV9FqivIDGBli1c4
1UbCfGYqV3FBRSbDyRZBSBYFIDhHfl/LzZrvNLVjTAgIQ/8S6dgIXoyZgOumZ2za
bzXHzbS6THPOic6VP4jo+NGSVchi+ZNqB8U79nOo3I3zJLrw6ocDlSdGTt2OpXl5
8ooBBpvzqR/tUo6a/EWqesEEz3Fws0hAKL6SB56aR5aqVNiBGScdRXqY+rpkMWTR
OjOSGKr/RjNXfm7EzkBUly8JDwafBe35SnGhnOeCN3QXMG1tXLISuaNeHbEJcQ/9
afHQ0fOC21nWvmgZbk5vblc4smaumyul88uM01yGkU/v4T3nMN7wLm03ndNNTAoc
7KcsrpZ6OFzep/Ulu+Lc4riaORyARaeJXllmEIknSR9Hz1hE7eDfTcKHx3S2IScd
wjv/NFb6PJb2PLTlMeBYilMIHxRY3cI3dob0IOYhG9sBzC+Q5viGuyvhjQTRm4OD
W/HuWgxdn0DpG1nj6ek6nb0CXyrzvxedZZVzfbjYOZ6PqzEvzWU/AL0BISmLExUu
v/tzLUEWF3nUi4aeHsHEyYGRJZtQLVPdj5hIq/IU2eihwFa4oukCx6LGyIMTjgYZ
AyE84LJ8fAPn6Ore6022AtLwnqi9idZcS/U6CATi92setq1qmHuLlnpt/4afTogf
gePfefj7p3k/8hijE2isnh90AjpOzRYvgE/J+hyYxKwXqh5TiqRpyOcFWBna6udB
KVa7AcOGjfm1Ew64EY7d1ntGEX/khS+ncrlYnlI2lJy82gn+ROmBm8MMGa7wHXKL
IEJbBekLdGTM8tjG2MRVtEKM6isxmLTtmGb1X+si34L5TENaRr0pVrHZmhHP+0Bz
ACT2K0qUd9n/lVTq2ZS+L8rQAwgdPfeBUY2XjE7ELrdRtZe2kSodR0TYAKRxG98y
RGJM5R1bIOZhdPYl7lpvBSxZc+eNWr5Ka3ig2LB/np8PO9Q/N6BM4JvBT86nCUZG
PIgNpOWCu/AW3V+npwlTI0pB9AaymvmIPvT1MjXYk7ZbgoWL9TziG+uOUtzsupVq
ju8XAt+2EjHjvMFM/l8yhv9dqPdcsgpS5FZITt5AbRipJfd7TPL99zrnBAaTIS+i
OoBIApSzn1EuoJ4RoR3twqhWAJZro/xmHbsZ6y+HMNwoztCBzleqmnG720EPWFD9
Ln1PIYTCOfuhJcYTUJlF3N8iI3Fyqe2nAUolhE9kwNP2u2aF4QVCKb2j6Xzs6uS5
O/UMldZ26jE7rFEAYPxAWBBFfiv0Pr7GyzIKR/115xx8IN+NtdiHLLWw9mkbokLA
KPTiMaYQ+UfccDT64kRS4AQr8uyCFWZAhdGNXz+OvH7m/6K02OWRgtg3n3gXOX8V
No/abPl5Z8X08CcCRhfxTk9ky0eepInofLl+MJ6EnUXA75pdINOrUUdDHIYF+qCl
tmlyus5XzmGPh11k9flPbY9afm8lt9owIqF58bR/sxy/t92JubrcF283S6emOf+L
kAhlIEdy61vE0+nx1x4dRfEClG3WPXcd0+Sw4DpCWrFFTyQPknPaQIrUVQNblKs6
XzmblnAqtqYsqGTDWO4jDaxKQfvbuIbTsUQLH9M8R3nTEDq/fHAy9Jn67imWUS+8
+1P2e/+RGU6ZsIkn6/kisEoHa//2/GdunMR1sSxIH7DA6YObPAr8jq5Zl4qkvX+W
gZtPrIeZM+WNPjAs9rFs7i8JiNeaDDU4bjiar7Ky2HaI1tA6K+Gu0kjvveE1/9MG
/gY8qV2SH9X0TpoIVDiw8UlWoUFI1H46Eu0P9Hmi8MXZIrHXV6BQ9vYcMEUA1Gcs
JgFLeBYqEnNxJH5uRfmzDkz2b6MhaO5C0NRhoVOKybDP84Nf4+zgBwbF206u1yva
W3cZBgwwfm42BbYl9UgUH8ppfsf/ttayHCw2sowbtjfoIr8n3JvzQvxTk/IkhrSQ
RvPOXgm3jbv/nLmOTMYuZWsnJBXKkjSo3XETtEV/F84of+IP8+/NfEsCXIMYc0QY
m7f3Q5FItHSrrxlQOpfYiC26ARJxtm8y1PYA/zD0yaFyYmSaNXLC+hI4D6Y5xFvb
nbCceCzKROVuYJJh++wYvgUfEYWIGVc5mFqT122sb/2HDU70p+R0W+Gcp7tKNqMH
KZj8j7mfBGoQApqPH77UMiaWTOa8zECle8g3DL44pDD3tzDfWZmCo/WS6fZdtWTh
OQqQC1dBUCcmYyDXeq+fJHwYMOfykHoXcFSo8Fn0VX0W2dqLMRIbWCaUYG8MxJOb
kbkGUuGdCvkdvkkq6KBbESpZnpDIiLUcaa4E3acST2xX6Ej4PjlCFlr6QhEK7J8Q
bdXW3JiHwXIO2dQq0f2ayRUHm5MfpMAUr99VHng9vzNBFlxZnKlM5EvHsw3TJrW2
zruG6cjrgFV/4Qw/w6GnRNr4W+dV1suk1L3vLoNs7QnN8DSzsVIWJzXgJ+A3ZrET
5RYP/spBytiYGdjm4C6A0hHbIB+eACBz/iMlgJtJCl/CE7nAEoSm8pFxfhdc9w1J
sWzlxtd8pJTdClfZ5MlM/L83dVY3pM8YtAwTJGCZoRBL6Gp9ZHRFNt26sEM1F2tA
wyzb7AdZp4A+7krdcp9F2hiJZctdLNqEq/lFiMsxdZKZ5gBQ+6DHVyb/1NThND37
Z3ON9v2vQmN6VwHx8qgBaLH1Mm+rD9nIIb6krkIdbEu9i+0xg495WfevdF9IhKev
o2sQW8pWhd/iWtXvOrl4UNPI6wUn02qrLGsNunSZ8tmK/y/lxPkxNjQXYM/hkf57
c3KDGx5kj4sWwmPSN39b8tzTK8+N8uWQcKRrBbwmq942d/2sTJKl+4bhhvm2hWxR
o5M5yDfHonDwtRuzy+dvwPDLkNkgkxfQjxThsdUmviyT+VyuAQPcRACeZE4ePX2c
520vzJS5/72RP8PxwbXxjh2bXaSgH1Cwcqy0uZesCXACtDImNQbFx+YwTefqLnv4
3jeGz5mLFePaG+2exB0HCOe0nz0vAK+XWxdEiOYJveKUFuxuwEy46AoIfbRPrIIJ
sTnKivT0vHTN/KUcUB65MBlk2jNgvIgC5Gq1lSWyHz/ISW6lBtFCSP8dzpOxudWj
gMNnD6ZsUHZOKEnkJj9E2zjCgLnDtQYotTfnRVSOAOpOolzc/ofvksFyuUT2S5x9
PiZnDJbpEUlju9Hc4+1aqBs+VccnB5QV9t31dtiBkuFjgxpasPx3I5TLagw1U9KK
MYnUQZAv8B0cXIatTJcW5cGwL6g89ECJKCc6EmX9pu2NcfGHNePPOuSpaSn5B5tO
w26F37RFSkFSiKXKJoutvoeiAAD9dUAiKj+My26h0TB26GpnC2Utp2ZHHB5gHOhD
FQY7Q0rwW1pCSmmMM8kmCGufJ2r9ZjqEr4Fa/QO2pU9g9XFATVWjVN7MXQj6htHV
0yJXIEUvCUzYz1uSqKLbw7f+dE658a0aFtX1+g9K0nJ18YlPrWPep6sTFTr/+kMl
x6FFiEIKxWhiYpGhFaKnGMrvwFGpSxrlNjt7G35i6pmca8hezIlm3XQdEkGSC4MY
UnAonk3vGqHk8RAsvLw7p4zpqNUUjEiU2dq79A9qiIrhwMnYe+gvK6au5QzQ+akk
1ULtrdIVcew+C/sMOGmCacjqkJUeluMY6ESgcy+lfchKTy3cldIBm6VCtW8khEn5
ZR4qr0Rlpg1CvWfzgFPLQ/WpW4ZaXfFlNGp9hpCuBrUXo62Y0BEIaNIPwZSGSvJ2
ApkF851U9fWZZQ43A867IbnhTue0ULO1BOMaPs5tzQcRx5GZn548JC6pl+y1M42R
As6AmBc0gdJB5Go4zmgUHRnW6u8oKxDl/WingJRg3jTibofirFsqSeFLDj6eZQde
dcayMEYHb4tHbrtZfUWyCxhhQdJanRyChE6ho1YJtmR37IIW3/JUjJHN5qax7Jvf
kfccK30Zeq/z6i152Dug9runk0MyzX2/JNYh8BXsp9OB74+i2PlzRqdvdGxBU1ai
UbFzeoUc0TqlZi4bLaxFAbdUGpH3++TD3XW+wHZqa+DPm4ZDv5t02r5MRBejqKTx
k7FrtRcEkHE5em6bfvkoEq4avNSomj6lYB6B69Dn52rHIEIEwpYALlZbhLV8Pz1z
pyNNyQHgDkDMYP7DC2rlgxmYbW2qD2eTn68IvwlVq+6k1TsCVHRnIzuTQAO5pEKD
LJF1D3Aw3yL0O+DQXCug671SnsDd2Q6bdisa/kB7rI/RNa72UJ25K/1cQlKjrMHs
ziPDBgcPHttI+kULh2uqCqrf9mYPPqY9UbkmqApcEhPGnZI6q+wAP7MSzDusJZvB
44nevrUodmafSyBYsM1QkYB5wju3d5YhddT/ChjTYv+M8MyjovuempWhgCtUCr+D
u4TKIOJSd78Dr+Q27g6fUIMZg5XFz72jvcCZpfGYdg/a/InxbQqJ8N9YSUokPdAa
HhZKY1b+BaIqNrrsK8c0zyqrZck93TsqD0rr4Sh+mEuI7JTiRZdeZ63ZBjXktZfc
+2tEsHr0KJX4ALY6WSBeDc43C5+/8oiho9ZimfqvG1ASkSV30xiQcaUlHM5uF4IO
L01ZQOceSlFli5M52OybH0XhLYbrdWnqeRw91O3jB8r32uPs61uubtmpWlkdsuXI
Sak3MoxuV99sC89YHj/RISpvCnoFRC1vHeXKme7z9Bf+7b+s6gXHxXievHv4xwAl
OaJ2sc5HF0tFLXh+YWqr8ul7BCP++SHLD3Ca5EuHkWpvRHJBQN3GfOIe8Lq9Wvha
IrQfr5uWr6JY355QcgxQniuH7JlL14tHfDR/UHGm+DsZmkHqk57BaAO//oCImB3h
kXw8D/VXZD2tEIDwOSgB7eKBQVgvmOtp1v+lUBHPGpivvDSJJB30W/irEVRTIniR
Rodb0rsHOotg5vdmh2qDi6RUoVyV+1DB1XVFYEeeCqxr8lRNGdGHl2jtMIAAWmuS
ya9BXbiR6PufdB/IU01A5dlkrVzKVvOGF8wHRtJl2zbamEIr74sj2D2MbdFt0jj+
fRkcYMJjNpFuxmMxBXsnsajEfSHJ9IYIy1eVClVHnKjjuO/Q9x2cCGHaezxo/32a
jxqVrzXkho7rp8QL/InUDpvQX5RGfFFVLv/N7pHrmIYhNyxMPGRnftAHh/HvsTXA
zOond1t3xxkJ520SCVbsGUxSL9i7PEC+NI0GMwai4EcHeMzDCRB/lTcS5KUzal9M
aw3DyXX+t8xKy50JfMS1in1VYMcOIC5Hf7Hmsv/nGsriSiBJAbxX6Twqm+x6YY+r
vnoTRnLJ7O/nCb7tEXmZyf2cWMioxheaqleobzaMBwOoz/fnCtQPaEVluB6ino8c
HupYgWy36I+xAU06L+hePsmEm+0ICKQ6E/ALYbQmZ8QP8+CLh+N/3Zyrgfc/9UUI
U1+2/PzT8N992NGipW0IFimVDMYIadwPvOi7i+aH+hBcNmTDrmsZ5OFKfAyhb/Ul
63sSa2fxImGYCMb7QGVSWq9iTT7sGb3oLf/EJvsex6CV5g7OW8akQWEy2k4Q87b8
ob0orSJJ11m1f2oK37d/vRsPSOZPsl0PRGO7f7fBvzZAUiR8A6L99Cb0K/pS1xFc
PmWzKf91mn0ugTAUjeAw8b8eWfffPa4546B4Lu8F3FZofUqd6wFTuj4rBu8SDa8A
I5b8VNqzmG2A2WiLOelDBNMJ/QNP5GEuVW1ux2l9//6S8cqNAxdNbn5X2LyMnFz2
CHzienuIqkIpYOFjRwHOZ4CmnccbTKegX6GNVaqqVU32eRL+MjND0lIvv8/KnMLf
XmdJVtIKPU9AzMhxP6Y+g4ZCAKRHvEhV6iblP2+ObsQm18J9e+eDa709ibaTiv5f
KOIKJ5SUNK3QbkxeJ5ESDL7yfp0D/JaFSBZap6SsgA1gqDTACes5b9Eb7MX5rPYc
evdj9Z6sXEu388TUeujX399BawGbz9HfVMgFpSIKJibWEWMCg1S9NhCijq6d6KuQ
kBxNDjbr567Hp6HCyaDduO+ceEx+UqPTNuDZJWWcNRUJGYqrteEtSis80B0tdu0M
Q+xDMrb3Ww+SUIkF9yDEs1kJzgq9zLlUie0JKdXyEnxeDNK4FCPTh2pdtrBMuIW2
3hP/+S3ugV7975rmVJNGLtKSN4MOQYApcQOO0x1wrWC0Epdc0+eAGuG1F8eeO1nM
N1PKMvQCaYP/PBk52Q66PfLAkbobO7eUSNCBwi2eMy2VkSS+7XJAGFFU5CDYeY8P
1YWezhOa9buvm31VFHVJLbXA/6fmZht1W/MuycsWpiR4DVoeQY1vqUI7F4mDcbu3
TZTCwfcnWqvNB1Q9T6WEQRq4MXTiWeRG4hCbrfWfv+copXamqzNhHdATZHKbFDJ3
g2aODtXVWOBZj5QpGTOC69g3XHmhGozwaMAh8oMz6yj621JIQz0NY+glSvQTkrBV
lVhO8rA6JMx9cluh610nTaQBaOJpYcRR0ThgRJd+MfYrdvY4pxc1mwhqKclFgC3M
F7/wQsvRtlghB/yMMTA1GynPoFeKN4+yiUdTY8XkgA6Y1WxvOPOL4YlS3anxqjNn
LomCtybzNtISX62CF2xse+OEP5HNX3Jrb5ULHxnN+yGRAhHzxovg40KkYfurPAWB
Lnr4VuOmO50L/jW03Ff/+NomAOWqgQZa3OE4EYcuIQvqHXu4ArIMaSn7kJlOaAz7
91LqdnO4OIWgyMYBQm4siNavBqpU8f8lc8NxKaW99CN6TJ4OjLycyZWIPYMzcP8d
5BxDYtCDQflY0JGQ/fC0aYdRjDazbkkwExsVUJE0GNYC2bVBBSvN6IpP3hvy9z4t
fqGAUl8QIGkRteEGSt/Wddv5o6H3JZ3mdNkZBB3kwM3fmczdJ7u5o7J+LpIQVc3R
YvMz49YSUvd5z+CUSzDGKQtcvWYJZLTYGJlOdLyOvXwqWQ7QraG8fBhMk2TQqldj
ZhGKUwWunTJVY92CIanBjCM2z0yt3GJOpxdhMcUX7c26eC1AY9uHSRuXkdVBS8hy
YofwSZVwKFuJizfkWcJTp27uMl21XQHD2buzcY6jUijsoZxPdg0CNJJljbzu0Jvm
2tWBHj8UVskKZyxoTGOFH9xC7lkL5+BdPaJ9zWrkuZwlPj4F6nngqxQNZWEG/SAD
OrZAD+VdmdSdQdYmFTUCvhg5YjPVxVgxrW+B/D95mPbPuNG54qeSIHYxznFVfrZI
mrqXNZMJKUA2tnUVOjpp8hlOljAaCsa/mQkGbQU/QFJycWMmE6EMDiWjNyzZ5QfS
tiMTpumqJeZgA0AFc0Oj45XJSEZz2IUYjVjp9jaXBsKAKi2bS5JqLf0bw+I+JsiQ
F/DiwrATTdiurz4D7WB3CwuQ2fKsxJhUPuyLOf+HLdwlzbD31vPCF9WxQRB7rI4Z
7993/gtLPnd414mx9ED+OfSqM3XM91aKtOwBibhQ7WQGjClAjmF5gCgAxze0ok7w
tz2nGfql7bIeeT/WIZkjC/Hh9kKbgg+z51oVVyu2MFadv8VZsmOKeyfwv0HIhRck
lrFf14Rb0k04dTGpos0qT07DtyZeQwAIAHdoc2+FcoinlQpzfTEdNrneQ5NhPwFE
PFmTdy6hTGCT90aj0jDJAHmcuraitzxg31If+cxpL2tyj8pFnhhDPAqbxM1Mu7yr
h+6Iw3yEYOy8ekf84y3jG1Wpo1NVjpZ/YzwoGG0joBu0cKsAOpxZOmTiypfpsg6o
PE+Bnf0M4W8bNBo4r5vYB9WhjoPaptT4Q6ReCBser2HOMrSp0dkFIitRuQtL8Qwd
0ffeV06b2G1ntrow/MKRQ7WKUUQkCuI0RW9I4AeYm88/kGwNFuE3dvRo2d9WLlr4
kLtbA11Mu0VuFKMQlLjWsfxiv6RIMRHpTVUisEO6XyR6IjPH1EKJe/BvgqXshcWs
KF+0QxFHB+Hl9m1y3sZHe+eUvp+vFnp/K3V7LxWUY2LGxRwGBZ5qRSCfo54VQTLQ
SXoq1DxpbvCRCuQpxKSWhfielD0u66WkT+FpcvYUmLU5iL91eABrTFUeqX1uh28e
caan5bAeRlj6M4nzMFkByTn22gck/cTq7GYbM9eDHLnDRgaRjQgEl6o5LE0evZxF
pxz+aBk1VswXiO9QbR+MlNUDPeidh+kPpvJ1LgQW1eT+n73xjhNZFekHrNsdOGzE
0cwdkIQ+OXaH7YaBq0tn5FUFBl9YL8lqJ80JP97E9/rcoQe8nhA6nOgsFCq2lT2D
pNlwmPck2JdxVOwSD1lJf+dh2fdpi5Ul3OoQpHJlOLCoy14W46qsckRxzK+bOAgn
FlaYIQ2ApnagpVdv0jbe/ujJIHZ44CHClhU3Iy4o6h23riwj43cnUuRncmReaTSk
Y142BlYutqOED7by3qGFvoJbF1J6uCbzFU3/wSEoW1MpjSJ8YIc5V6tZPO6LW3PT
wuYEo/LiS1dTLyEWDq7RBPf9Su2GhwgEAL2cFx7sYDG3SXB7zc6mXu/kmu48Kdya
JxgeVXcJt/4E23m34n5t8kaWuRPep3H0H5UKMe6nmmCIMpSW53GJFpfduT/894AV
KTHMMvlTD2ODj1INgmZIsuX8ltV/VPaKlmYRZPZ/D1aGrpIDKwUIwAF/mB/iFr6l
CcSZvVl5SHhWtSMfkizIgcSuVNVISRuYVgmAmsU6IdBplsPg2YGz47CrIghLWT7C
4QyEXJzlRp7lGJOfMW1F/PJmBiFKnwaY0vCLXXqKC9oN2aUg2LX3F9BcMXTV7/3h
K/lPlZCJRPjqSGl+z//ZmS6SOmow4a7dSItknFVWPMAi7//WTixoekONtpSQRhGu
90Se0djDxv3VadmQZBupTsftU5QmRQCv8NZAEhe4mjPqGiMbCLJsNNzIo32NiL8i
n28Li0K8bESbyoSSRUjt5pkYXbMTLrrTHxSsG/+RSIkTEJnHXx4IwqHDfWcndAMP
qulysKjMF3XSNePEpucBkJwY+f5lRkCVXTqEHjpO5T37Lm3XwvtUJCuvCQRv7Bmz
uroSof8skhTiqeBzSRNv98eUNCk5C1biFc6L3Hrb89XxoSFF3gfrMAT/p1kj4C1z
6MCse60iyxwNIZEUcna0xbShV0FcxiDvPVdUOx4w3F/p4pxeBL/5/JbqaawMl4aJ
8BC16cdvkCtknWjkehAzB/OW2NrBnoGhHStytYq69Y3X7hNd1TB1PqpEexwK7vSE
vtUBvWUdm0jTj3vCNoPDRKgs5vUAjF8sIdJrqhFvqfSAfI7w2qXbS7jsn3ksxO9o
L81NXkkViZwsI+3GoneTFN40WUgeBfVQcJtzMOhAXOzep5WjBVS9PsLegLmOQBFZ
twqNGUAnDKkevETFXrwL4CMDRMB55IGj/izuUdAvGUka4gMK+SQjJ9Gtv4S5HOfR
V1WWbDhWXphFL4VZLcxK0Wo91HHSWJGk4Ww8YLJUmQUGWpqmvbTK5ZxucbYSuW6f
9MleURWH8ZIOaklX2eZg3KEAWwh5pne2uGNQ/X0X9JXaAQIZFDyJKU+anqITWJ5q
aCPyVPuBuMUXI5NMMkbm1HQbg+51zSbxlf/p/HLmMCtdABYANxqaFFfCN/53oQgX
qdRS+v1tSBCNjHD/YdS/lWnq/naQdqg8UQLwdlEGzms7wYvZQpjMj0d5Q2JmKH/X
p5QcJcxdFh7/cONrWmrAHKag6lcK6ekTSU5CYztZfWr+AzAJ/K34xdws/Kp0PTlF
B/SrAyibSWBqyQqokQHuY4oL/0jfzbxWw2033ay3LQWO+bQD4+9lFVxLYCxhbag7
fu54eUo23B7d9/I66K66tlTio8ilu/ScCJtgjkrRicpKLJsDn4cNxveVyvxRydw+
zIoRcGh57ec5ENx7lz3gd5LVhTmCV++2Mu98GL9v/2Yl2ZNNA7R+u2xnbglcNvvy
cc3zZFeTNQwbyPd2qXVYi5K3EK+rtbeyMtdV3WfIN19NMlG5JSqGSi44CBpB/Ypl
9Jxt+/VMfGoYaliDnbZCUk/Kqm9DWJ2f5QTVZo7pqHjrBKHxTyHfbPzZ+tIST5sB
ceP/Wxgp8PuiTlIZikgrjdhYU1WFjRv92CApaDl3SCon0+RsTPWNhZjxal4RrWJh
dWdlFQEYXXfX/7Hd0CcabtVJ0H+0Ocn8nfDHLviQGy8HxXcBQQcFU4/gc9ZKvC/t
lDGAMgsl2OL1IOlYugSR2+aRUqFvdD7Y8wVTghnMiB2MKj83tPK8ZRsyn/P/YVAg
TmrR//1l0VkgbCJrabZ6l8h683V7ITMe6rU4Q8vycRU+TUba0WNgXG6hUo4WKG+L
OXv8U6b2+69NM5ONroXatuWc26ttaPAI4l/nLuA+94FL/llt3fOCJMyd3tgynpFF
sNTXrOSgpyzVnhXH3NaHP6t/KelGnaFhe8LZW/5wbbUvB2Y3XhrhsM3ZhXPJQRXL
s43Sm6jE1wXeeh+CqoNmSX86UNW3My1DO3lv2AyAL03OtUT411015JtRQJWda3JG
YCaZZMlu3IOJWRJXUx/UbdKYxCBcrhlsYRKWFlzGYwWLq3B7CQqFqJnl2RO7I8/o
gy1OGuJGH2oqXQX2TeeNwt4QmpwcgAdp5vmngsmLQ0UE5Os7YgeVvEOtu/nREwtc
7uDcCSoOxqByAVdP0mKjGSu2AVNwK73hrm0xI3iE7aazud1rVQBlZnWXHoyH6Wxv
xJSZazn1C0YyP5keXc4B6HCcR8HFnmQqvTCizcpUvtE4it4/rQQUh8EZfqokCWzZ
EVMBzaHP0KJCZUwrIUYqSL3sv45nw7yvvbjAhB66QrghchfUzcX3hKyX2VbhEvCe
/uybQmBXTgrdJNKepQy8MrtKaiaO3Ut/34xCCkqMnVRyQn/ka72AertbfvVWizwD
w9oP61HRqnDX7hQSgALvhrIiK9OnAQEum37ebT9d3TndwUYK6qfY3UqNPhcTLXmM
UKWubDUCRQHywJkJfeFajNkg76GgW2iOdt45nxfnx9D0fmaqBA7kxVY90zsjf2Xy
YhqAS7AlOpBudrWakCRS5qohVjSj8VAXbsYcU3TK5qvfUYkr3NyOZ5y1GBHjzbTA
6iAzqUmSMPkVT6K7aznc9UjlUuQVHjHgPfNdtoFA96rR97he6zJhAITRawivQbAK
a0QFQXPUcN1W7YpYtDIgADCddPzs7W2msoGJwiczf9L/IuURGiL9h5j2tq+9WBZR
AWMepNBAS8eajxayOxqKlxYXH8+GS9M3BpI0q4HvdJWq3uHGduma4BGw850HpSmm
IbY5gX+SejdRAvjOKn03MR7CyAQU0IMI9z1I1MUWYDM/aLrvRoIAis3cg8GDuS1W
/OlatOp0ZOwUc3T9xPO5QEnmgqKDeTeQLvzVFT6zFIk4Rw9ZOD8WSefi/UcuHlhE
t98YK7sLDk8boJx9rEOXvCHsZD/p5B6AcR8o8dYMwgTsjebSOFjatHP/XvI9FVyy
l9oyzBdJf/MlG4hclYn7zZQigYGSybmcd+CB4g4TRW7MMYLK8JsmVnr5rB31lkam
gMCatawwJ+7aC2rDqZ6PQlf9E7FObl2WGzlbp2HeTEgsg81fuXPC7OLoKuNRiEcj
dLa7lAeh4ashGIPE4wSF6JTOUV3+YIXueknxVW7VDMI94xIiqtneZ8mCRQFsHudC
T5ciCH1D/NK26MCm/1OXwHjb7w+FPzSvxc+FF+imUsxowgcYHbdfP8HinoGMfwCj
fAk4qy5yG0xBAmTkqil1oidL9Sz1yZQ39NXsznzMnR3X6qxb0kapXtrV87+FuvRm
HVIHUBknumySnMD+db7tsmefRavDSFfGC8w2B2UHgBJ0m3cXsAfP6ttouS4YjyFe
8P4G9rRy0JhB8MGMRPU2D950BddemsPqx2nkn8pu44j1McOXMVxnkxKa/HT7px6Q
Ja+KxjP58tmyHIUfysq46uRrHOgcgOXckOfTmXLEt4sH/JYuj1jN57Em7ej3Jcza
lcgwt3h9a7/OHeFRdELnfNbNQMUgOyOA/YM8NYfhalG8BZe+qhfqT5jN+hwQrUnM
ik6Ju6pxL2LVfFK98uDahZDowV5AyzCsZQ5UAD/d40Awi5kQX9TPzaW/8c16O3CK
GgMWSxccohEgNeVsDHPc4RQNNtRJXX3Ho/Pb9da01RyWWr+0VQLc5sO/vw0Qq5X2
uDftlooDzyJPmQlx6CrUeTzUeS+XZR2uJiIzedeIz7EGSauzhUCtB4ybI6kOp/VR
xNUSZHxj9v9jIRzvLBnT5RMWPsCzriGh8vSG84KMXcqsNpCrd4ewLAkPyNOh9Zqt
N9Ve59ZBtwgksvAs2NBmWLX1zigZ3jpFJ/VJwYTOEdfHP13ZnyX8HwhE27JPS5Zs
IwVltCR+IeOo7R9XdK/dW8OwSJSVflgM6m+1NeqILy5rrk8rC/NDHYscxh0e9mEN
1u9a9mz7rFHwZ4ektztnAY6AE6i3ZGIlftwsF4OeAiH8Dyg9qcp3QXUKAyfUpHZl
CiK+tcKZmuDi7rxNrvnoJrVzU3viPAeeqD9+BgIaUnIVmplfga/pssLW6gKHOeX5
6JiWY413Z4aHMUN0rwYh0lICyDwkNKorZp9BXhhBEvZbtWqME+vzmlLA3QHdfDgn
ZVKw51XDUP1G97EJiz3S/CFk2kQZatoWXnYlbvuFI3O/8x34xqGCgX+khnlJDHkI
ySjJcbgOxzt+57RHHEWOlIiOIfrA4MlIFcUgTzsxSXTrD+pQLxNxj98gIzSP7VgU
RPMPHixAm3DBFPNLiS549Ompd3QF1JYNfQqJITHuB5ReZr/HLl4RYUE9NzXVnnte
Z+GkC2hsYIbAkjWtJWGqeeHb+sPTucEWT6/0x1vha/X+7/xxKDDwzyUqiuEx/Z5S
WFATv5KeIRV7zSh6LiMTqEI8EAP8SUxoIAaW/3ZAqZBDRQ1oDGoaIfAeWar78hK4
s5hBDsO9qi/ETkQdnwzON8KpV+Wkcsi8w5O4QmxGEq1p3fzw/m5abABzEuV816tA
fGLbTWxZV51RMhZeLxqSpZnTrnR4p9s5ngG006ZTSygBaZdOeWS5UkGeCxxo7CBf
UkL7KCiJtaMnIAcMZ0a1YJ7dtUIcxgcnF7pGSD90w8ndJNqZpZMHYhzQVbE/zR5U
w1kUYGqYwa9X2aZNNjQgFK+MlXI1PFoXr7bOd702BOdCd/NSuN4HCOaWZ9z12HX5
jq0Enbled+pX//fA27Riw7/k77jGdF1TorNld+knyBCWT3y33Tmu4V4bUGbiG75v
LOY2x4xtPaPuicMzXVTWNiwS4vV34DJDYVqtkjv/E/NgdqLOtWTVg2oLDTjiQYJi
8olqQgVDTczk1j4kBxmhaMeRlDNBhVXb93b08UlgibGeJ6Wrf6fMSQI+7UqkQXW3
W6esXpBleSRYcDCElU3QH6gGftIk1Jx36uzRD2ECjXXuDWGnVfD/4OUrjKVmsJQg
i8iS0dqHk5J2IKn7wthp/wZoxAsTgRYlF5nStoeUU6eU88J1gpT5WbmGf5KWFh9r
B8ZAZGSIkKzqz7dd/9oTa/GAQDiUOE+10RcJCg5J9kwp2AbxeJPM8iBqDBSgQgE2
tWzqRp8JSIPgEMsARjsr8p5iJEdAImv5pXnTT23XMWpVBC9rI/bmSybfeYC2entn
ps/qDS98VQpSbiWmeOCtiKDg64WDZDoTgPzMEaM/Vd7Eg1Vxk7w/ixGArjf93Ft3
BOoA58Yre443kltdSqiY4BeWZ0nC4S+yuRNXEw0fA4jYYM0XL7ZwSrl2TNguFDd7
hzCThp/NRctU1mDkuRrYm9LRuQdNM9w8hB9cfE4yzlwB6S+C/gDMs2MMOpXnesvO
pam6PL/bRrEOSO67H9JiBE6C0kpcYuH4A8RDOHnS8USnHaI7VeIWi4TntOH82YpU
IQpBMqDFeQYM+MvdANxESdB5uyz8TdUsANzdhvCmJYEefgnZ80GEo8ufl07zp15r
Kwc4+luC6uJmtC7Dq69jrUzXyhADIBGpGDwNxD1lHveWgeh6dP4FqP5Uh+Ddt6je
9ZW22F82VG4XG0hXpSAo2Na/+yYO+a4CptHv53ijEG1R5GXPpNRu2Gm/IIp7+lRf
rbdZlf9CV/eva69I4vQMGTp02GZkrETbAzaMB8pZyGG9TSRjk7MFkLJ3V7xDRcGB
h6YsMoWuGXxnbocSbadTT+LUxVyyZKpergCGXLhPMBa4ZWPUlwPmN0VHGl9jQwIM
ccD7FvDW6MjjPXHJDmKZ2OuEZT0SyTpPkMjy3ypvZ22Paj1pFYUJ3VP7pnv4f3JL
SX/Km3Nm15rAUQ9leNBRXywwv22Xgbf0Nvg22P58FwTbd3uRSz+WuUAwWLi8Od4t
N3RMhxvVU0cQvjMmhjZJsp4pxKKQQmuWP+fYdfEYky6mrvX/sxfexBgQ3i0bifkI
qqZcA3N3lyCsxxwEw5+EqxFCBIKsGvli5BIAL1wRQPLYC6GW24YfeLYdv+4JtaGj
m1ExrG2fZu5UQ4x8iyVwaubLIRFrqAd6cWzaFZpgplnfCfngBps4WFFlmAy1NNvi
eW4uLFB6f35TXDGDAZTOA4m/7ACqOYFLPgr9LgvZ6kumpKUoug80+PDYrNqswPH3
PR8aUtfCbUpFw9eqk085AIkRioaVajj7KzfU/meWWOfTmEt3jF79mybdgeHsvrRF
Rc/1BID9RNtqAOb3sUc9F4tjxPCzzTveQ7V+tehw+Y4yVTqfUnqN8AbSSXyHz4eA
5JTIMx/fEG6aulmnz0YdUFeU/lytlQnLxwiqgyBtGWtQkga/bouuvqqZNXjz3cKz
2HNdSlKlbPH6J+ElK0/Tbua03upmkc8Cit9nIQ8Zga28Dj9Deg8R1HOmHD+CotMX
87sVJtgVeBuW2nc4AqGAwLMIARY+nJyzhpC+cSahhpp2Wju2NafJ9RiB15gJahvA
P76YQ0mzD3ov7GaubVAVD5SWhGSIwsJ0Q9STke2ZJVUqnXfsneVtsRblXJy6udzo
L56mkdLU9dSFUnajwszVQ03US9LrWnxAeiXvQVI1X2ct+z+qLhT3XbVmOXJ+tZSS
m0+3ffIGq92q2WiX4AuEyurl708EPv+IplzfWdDOgHQTAh9DonDERO2nLV8cEryL
65G46NjfO02mFqvRO16vnLVDYo3bCgkwRHS0piokStKxfGEF8vyb5b3JQtCTdTLR
wVO6i7YtgnMU9WPW5t0nP0JhbQHqpa3ikmeMdEWcW7CXYTuHS/7JkOvkGgANfTKn
H+ZygwOOLZiHfkNC+Cf8cJV9TPH3SBNrJpqa6KlY8PFQH2bVEBr9dukQu4Xfon9R
jnttJ/XAS8erfZMbbxR9CA/FJG56e3eTMfUtsKB3krq8HD4Cu2VdXo4nvvIGv/is
TeKo40f5PArKhND6UIXCKrGb2nGIOxXSaxoKFEQw7Wme3wYtbrnaS5pnbsxg3sYX
+IkKc1LjEGtpZ56yK5qd43b4BMYQ13NDvj6hHtsf65z+zeIJg1L1JlElUw+wYYlR
LNczOktrNzclqDohgd4Q4J2KvlnGPFjtx1F1jcLGqz1psNFB+YPynIASIjx+XLlN
NBrDPlTvz9opZ97iYI2yqSVv7eMtBIsGR25FYBnxFp1BdLiR1wXdQAIes4SHIX90
iOybLqpQnepnZnGCU1FaPsohkgpCUO5/HGLtgsx3bjCsxKwjnFh2SEAkJfqfyKD9
i1FcQtDxv/SAXXbvCLI5uThKJ/uclJiKI6ik7PieGdaCTs+k98ByvQ2030PToZxz
5QrQOmHqGT+MB2EvQBOkLSNZAaxmwpfT175BNUSgqOwx3G9gEhDar3i9tPDLNIVK
IDBbWsND2qsyoY8Gr22AhnP4ttXSAWAZJxxxI/uh53zX2xCFF5Gg/C1MlW51hkyT
IlOslc/OjSFv4AtStfBM6h2zDOJU7ZDTGDkq723uw/69wky3Arg6N8tFhJc3E5g4
Dp01lTMIrYLEQkr0Pfa9qUZ6KJ6f+hzs1p1AbD6VAxaGwiNzjDR29l+Ynxd5xc+T
811xlVsjMRGQSLK8FVRkR+7hQDUsK8U7b0FisZLYh8U4zERh4+cGIkkFltRHBNZV
2rZpYEmcVaVYBEW3Z4X+/G+5plAgtIoiA4G6TqwapfRoO8UmNBDkadXz2FtyhY7W
Pr8vJFj5oSe+o1j1jMUl3a3qprcapo8/Kn9/ZKlYYA1e7C9XDQ8PVZCTpzEIAAIW
8tCQI/xo5dOTEi3emoCV35UI4Q/JHFnVMcyHNLlPMrg2xy5wT7AtpD5mZH0FQ0AO
R/IbrYQlW1au20WTrNMyAcybcBJc7fLDZLNvNwgXlJPAKRwV39u+qTP3nY7gnZPy
q3HlIsSM3xGV6/bQ6lWKo+Ryg1UBgrjArrdTOIoXcnMxU2NLWNuR/lGYgbrMlVLY
ro6pbyqZPRAog2H1OQEpB6BzYekCJwKe/SehdzTVuzijwN4j3jlOoerzAfGn0Np8
uqRzo0T80wcIAxx5RKanup4Q/F44cFjixje0D24wpicJa6MQQWz1PoXxoSBaQK/4
uwz75ETCNn+dPhgmZo++ewIYhAjSbxPN80u5VzLSswyhvYZuU7A1LNP3JlaGgaB/
zqE4XWAi+yBKfmtEBi+zuyIhcEs/EEJa9YXmgYojmt5j4FpGORitHYl7N7IpKAPf
V4HzQ2d0HSqs9KB3pkMFosub5PypGyEvtXkiOac3eD0FXldp9zcxfYeNhb+uiLAe
67m6MlcI+cwID91WIfRhLk76Q9Ef5oNvuM0Cr4iiOtjS/oVK25TYIBhja5Eas8ik
cqt/b5WQJynSE3uKUQ7XgjvNSdhbRWvwecz7bPh8jBMGTKLiBN6ujUgGdBwAHu4e
/jMTFdoLfZKDOZiZ5Sdns04vu4O2Z8r33XY3JbkLUBnVohf1sZXAmPPeDs7e4ZNB
LPEceVVqXVZYRWiRp095e/lPh1aZU5oiuA45bBmM4eKPWnj5ibn9fv8M47PSrE4Z
r1HNhRlxnwyS8RJ+xMRT97g93LA6FgYDlChEWHMz/ufbI3l6JxsVE+pWPysKkvX0
IlFrM/1ME+d14eQ7Q4iG/jmyAGQk+AU1zxqAtD3DOUKfV2QSJtWWgP+bulYSOOMg
hcw2ZN65iEx5ku2ZlwsXusXG60lXmWGoNMKtD8TkcLDdBxmHR+4DkOt7EqwIv11G
YvIgiD9FUou8KcnyBSD0jQsIRf3Bj/tjRCMN5/WW/HngXNzBhKs4pN7xLgOoDppZ
6uGl8EUzyApJ6L0wGaLP5eBz54gMjBM7bZLOrlLcTGV0Ym40Dw5AmpcrSz+zV/Pk
YKsFUfHjfi9w/HhGZVIiyuyB7Al/Rj42jA1/ZKS4S9YpwDGhS7A/JQ6x6i0tn6Xt
+KtDiuyRC0YwGWuUJmIkSgRfZ+s5FEkxWZTvc5I8HFGPGHo+GIzHAhYiBA4fRfZO
Uu4cprn03RYgqsbx8DqdPY3bjSp8leMqgeYmPMNE5bOpQYdua4lYTa6Tx1L5vcYD
eHUyCwbkBjZteB2Re6ZUHZZoh7JNc/OJ+uJSd9qNONXjUvuqW8BGpXWtKzc7BxKt
k4tQh0purlI3Lo+MF1nt0AvtbQ51HAw8qsKE4C5S3LaZKocjCgddiqCQSWiveWA3
ViYsLdr7y/lGLYkKos9U5omslZLjwwV2A6kDIC6tsMh598gngLpT0sLORhyqwZ32
bGlJqmcKdZ6rgSyxs/FoISalka/BL5BMW/Q5zRLqU0XtTxw3t6DgyrXdpTfQTfdT
wsz8X3p6UABQleemLeT8qqQfNL2QkUbm5EvpcQq4O++5KxXgCG1T2a6LY5WYVU6r
RrjDkMi6guYZpmv1b7AbKIWyWqGG19/ZxdKd1lHWN/cDVre2XQ+FwbYizr9okhOn
v7cmVqJCxCrh038ug0WKvcsM9pDhMeYcCNY7jAmuerwS8JfCUXQfdQ+wauTSSvQl
NfR+Q3ShngHCGJPqaNosxtY44J6qzrpPDyGJQ47LCnIobtAEI3g2kNGbJU/Bbmxo
VCYeXkMARecOE1ctEY2aeeNPHHad8MdwjTHCC4gWGxRYNFOcNUTPss3vwyJdUGQW
2yJaD6b3JU8PPZFpaMcsjO3MCd1yHlSbEIG9Un63jzQ1v/KvoLSU93DYC8xYFdxJ
an9q/aFqBAcBKhzp0/Un/pnmjx8ktZLOI9toVjdRVaKEuafVXcm1s5WdfYtjfjtF
tPGyuuVE8p2V4vJ93mc9D5maTcvlWdaVjy+qo2qSHyNHsw37ymVrPlfdXIeNalJK
+3CYvaBVdolaekWSsMzltFSeZ6zrCtr/cBcg5hs77MvhZdXS4lzyQ9gUWP9o8pqm
Hm1Fe7JvnExyRRDur2+FXH6if3A0JvydZFkYx9O6iV4A6Pu4xUZ5qZgc8glDKqeh
JzJoU9ZWe0tiSude4o0sSmkTIE17ypAqIEgCoh2MOc01WkCQuUQ5Q4DnKJz8MQ5p
A+RMSiwHpGfMBsJFZrAUN94g+WgAL2rBynSmSKjd4WjC7B0qiFY0glQs7+TyLnfF
Qs6RjDpTwXNZHNsvnXDbS2BXTGrZLkiG3W9MooMJcAAssqKEh4kkqlH0G+NpWipb
M5TocE4Nlr1nYC7o77yPISi3CdHdEEadiWUVY6AIWQQ2AFiG+PENOSNjDX7yqdbO
Z5vPKmotmvYJ08Y07tGNTeOzKoLJC+7dOHov/9eqNd6nd8hD0wcKmKWBsvJCYgV9
xGhzLHq1GEe2ZW4zbFkYDjZiG5XRd+LBcMMeIMi/O/kE5a2LytOffu69ppEy7pWM
FruwKX3l14k77f9VlH9GaqFdOluiQg15xP/QjOeVIw9HAitlp0ymUnQLLy9Djwbq
ww4YISYwMTIhmnxbKvF4z0vww4gsvtowai3a8HoNNxtBSChb9fMkKPAwbLmoekmC
O/OnN0BpsCGXZ6mcyN+3aPFe+dWOIYA7Xiy4T4zE69J9vRpKmEnBY1yXPZ0DAvtJ
ycKuJEH/7asHHiuPfNwBdOJLKHahCfKyamSI6nJ8AbcQTEOIJ+F3w2xEF/VY1Wpa
wAbGTYNDX7f2EHeMRhLFXMRtUFQFTUdy5XzPIMRkVKYUlSgNN1bB7SLvvPQzzAMG
2g7TVbVrR+ASDX4AV7tqEN/navZhiKTMTL11fcWURkgi88MxUazr7Lg1tP4yzCnb
pqTGQrV2OlK2NVFMqO93sX846tUFeG3872k64xkl+OiDymvRlmXgo91t0ZnTpycL
8a1V2E4NJD6ZlLOWi6A/NDtkRfvg6M88N7ZeojBdG7pi7QofcIf2QTLWjCT6uwIB
IHAABpgnKAH/rZrGlDt2i0xJ5jClt6iDOn9apTfDEAvg+QoNcp9zOUWwOT4PV6lh
LR4pVQYOJXq/LICdwoe1ZE3KAeY71CDpIxnVupkqvP+f2KgqYq1nzASGj/EKAoMe
o0VJDHrbrXxM8kmdntcBuVEITwyiYAmma7WxPYmsVm27dpvi/u/Z9ZJZFt0uDkSW
yzvQMtKK3u3QCqfM2cVwg9IWNX8rc9/SgOdX8rpDhIKPWbroSv8Xy4OOrFs8OXLB
JN8rDGGsTEJbELxtpAk2miNIOjFQ8P8R71wy0rjw5p5HDvwqAWSrtZsI4b4jjY3s
gXxvEFi9KFITTinxyQzD1Vk0rgJ1CqZiwno4q/JhZ2xj6oN63o0HffphZx1nPtqw
Nnm2tZuJZK26InEnGynr0jlBl/ENElPq7jHU73vCWQoM0cYBMvpw6fbXtqtDQY0t
FeflbGbQFG74pPc3lsp2IcnLqX6xT6XUo+C9NPB2PrXgyUriXeRT9diHfy6Yf2PN
Qx+fdt69cGAwoyp52C7hrYd0468CEd3WVPWz2qj6dhUUiS4RG1Rz+U6ihZQZnXb2
ZlV4T37ClExoQwclX1uZ7uCgKr9j8BwzEQiG9D6dnTIdrTuTTYmScs/QXXBtk8CN
d0BVPJXTuDYUJtSZ5MJzGBnD900WJK136TPNJ5hV4GdioadacMyod1wXIjdXhuWH
v/ijaXQgSPF1Hc3hzDXFhMxuWYDF1TQnIfKHNNph1NyFlzcKWf4b2oJjbF6jt3Ll
Wi0NqnxopYklJNx483NrN5n8meDVQO8U4nToDmvgRM+NuasxNDNl+TYVfZ1n53Vw
WtxMijpsMMw6RifUOnOp9z39HvzeEix0LXSCZf6atgCwZ2az+ms3djftJ1CJfPKD
qGhDhtI3eTQpf6L5R9/be82eVbxnHuEZoyh6QalAz0MHaHq7eizcbGxMKyjC0zKY
Q0u7bOL/+0HWw3FIhtPGRd0QKXP5yPqfQQJ2KWqYi8/T22Jhz2JjdpfDlTY8ktuz
5OxcTvE6cXTYk/FWnOggXLGaYfdTGRtqetB9inkRGgWgIod3EzQw3fK+Ip8E2zX/
Uuni0YrS9VPTDtLsms8LuzCDCW2UsDe/iK9mZF1z/A7MC1XvsEnvLrqvwaU0GNBC
tgeryR+wGt1ckqcrId6b+7KsMk9qA1NIaAurXK1hNzcRl1d+cCmvJoOiAzFUtEk4
Ke7Ow2f4C2B0rxkdoAtbMc44IPvgWr4KclgrkOuwc4/hCg+4c0sYGN2OLsvpb8Ew
E/QuNWp8JvvlAw61VMSVCsk7i4tYIf+b8DtwNB6RiLMiSRvl57m23h43ao3Fi6nY
Oh8Z+IQw1TorZSWRWFBVloZHy3/sy1mhASvZ5NEQC98rG48JT9a7FTbASwfOT0ZI
AEka6khwzRjd+QVCANaJeaXb7Nk+j92Bq+V80KOzkMymQ5laQ1dJGHXGNhL/zbtI
DI1gsORgNPWZcDCfXiBXGqAe0jFbOrOqOId+yyAwsQJ9uRpv/N/i9I2A+SSbfk/V
qfjeO812RXyVvMSkmAcBQRmXsWY5fkEpbRAyYGJVFOtFMokBxz3oDBkQQG2ANNTo
0+H4Fyp++Cz1069CeztMtRYWHJ9eTIqLehW/cR4QT/Jli3GAH9bVnLsqgHlaFAcg
MmTpsg4jQxpLvQ3tC0gpt0UcEhYYxes/cvmkRL6ZhcwQt6jYYDxNV3g5WHdPO6cC
gMAjKOURcAgqsHhUlDUTYkEOhqZrsa0bGM35rlbPdGp0VUz69JOWwGQiceYgysl1
Vs+cgJAH/22cv1h/UJVrnNUz9iebBXbQ8csPz1lo//dnfyY4wvQx+LXeD5ieX3ds
ZgEOeKC5qv/OZoL0fqR3KkQezEJoLLEaRwGJ+oUFrkYQRIr4RiyKgMor0PZqKdJ1
zZQLlTHXn0NBieOrdE4z0LQ7ov14wlgFw46afmGnWwNIZjF1S+KRfysIhP1sHaON
YZhv+fhceNKd5ug+kM+g41M/J73euKLiipSzjEiFa2/9X47B/CZAPkhwCAZNuqhh
wv7n2FtCmde+4Fp1XdUT6nc4A/UbVo3Hg18r3L44d9Ob7K/mKUopMRVPArnc9bgk
VQRUiZsZrj+jgGK15SoVblkx1EauriOOPpRMbqQmLpDJ/svgINiY/DBo3Vmfw8sN
qe1W5O/l0AE/KO5fo7KkbVmZQRg9x9HKaZh1ajkuBHBniYrbtuCXgxSvv1veou2r
teIYXrRNGf/m90ND0e+sEe46iZH27q0ajzc2ckzyJSkcsuvAit2GakhjSdl+u9cD
tbI9jqWHuAnlQr3E38PvP/gG55Rtn01nlvy1BIWUj+1V4C2I4RIIGRQB0P48trfN
7Bno0skSFfic1n6uXdzgswETzW6qqaobdtxkd7K+VWIe90ts7033KghXik1eGoJy
6w7XHEbY14Y2ehBSqXOQtddvMT/i7EbRI0s36WkkUGmKglY9LrT0k7paa8pbgL38
sr8W9qX7+lUntQACMElCYZdR/0VtiORwcDtt58faR6KXbIiAuAih4NoF1RrceDsB
PPzAl9vNSjaXWSTJhb4x4+uEMU2KUcFHD2r5BFvfNXAqs5Do6kIJtAqeX9kdiSMD
4ej2B+yWcdtk5BcvU0PPkSID8v5jpAd7M5+XxvMa755oBq8aJyouYnFtEuLIRjxd
rybiw4v5KcdB5GmIQU6LFQaIr1m0YrnyK/BDfcJ3a8bxsj/C+c8Cra7h6XKy939C
WeOLH9GYMO9I4WMwiC+Fyr6HVll2BDdiYSPNVcIltBJyJevc1yada7AJxQUKGLp7
7GhZMhkl+1v5mEw+E9JWzKI6pECaD/nugUIT09+dd7MUBouxd/dXIc3/bzAhUko9
66wtVftEFUNiDln+Rm18QzeVZcDF2iKkS4lS7z1K19XYBY6UvvPzNmKM/8gArZs1
hpiRslpmh97nMgfmQYngRbL8XJhY/smzvrp4497LZ3t9v03EFZjdS3EbNu6s6q3b
sf6tDymy9c+MoxENhkqOzuG1RsdahqBlEdZM+tOb1/W6fiCTPLGKmH07vWq3UzfP
U+gj97+dPXUye9aBlQL7NRJkEnANyxerb/D/8Tjgy2HQMmQfQJyNwyAVEpRzXrZ3
IYH8u2FeGpuO5/RVlKaEBZAXvFqCBPxqvjDAraieO7pBgSCi6puOfBY4Rv2FluGM
93gAhq2/VvD3yU7Xd73imPVr6I0hYErwIzQyAqkrxwauEEYMvL2qqk/I49ij/JPF
7wNXp36U+ELP7woJY/NyTyBNwrp+PInymMHbsvU4eoXfxhB/gsVj4nf7t0LOygIM
aLHRsIOjQWjPBrKxSaFL/9gL6AtXcETcrsqTzljw/mFWsCCwmJvYQnr/4i2+F+Yy
+1Srn0Z+0khu9IYcxKYMVnXK8iC7gZdNYxXpEgbm30opbglWXS7HmtPV9ZYZb1mq
99O6pbGnrACdP040lYLJqN/wtDGLLlpfh8ltKksU5FKC081oZgaHOc9SCBKhpFva
F+SPw2uIu0157M6A2ddVLOdb3Taxl4dzc/3iInwQYDumhH338ckDaKDro9EVcfRH
mfjvKrEKLtql/XBq3sQN1WW6G9n1LrPg/vwsL7wozDTgY+Zlo+DldHqIGBr8Pb9n
Qo4v1XNsBVG85IYQjDE2gs2Hv05fR8wSX57nJgU7fomfqL6NSzQZdRyJgeRpRO/6
UbxjRL7zxprTj/6kDLnEysvjG0KPMGWSK/2GWIe2NuJoMlRgmD50bCf/a80VLCye
W/X1MUoY9VEL3Vyewd0MzrOo8wYGp7408zP682KLblJFHqPV0PyNUtTXiXTDp4G9
iDq9sS3YCOwX1IRGxhsairMrtkwoHFtNmwVwXqg2lKrpHHYSpLTJ6YlRtO/NnYKB
gIBWrPGxzUsJRX+kXJ/7eFYdkn9h8sYGndaLRCOT0/AP4uF+QA8jnrJeNRpgLxL9
MQDnzm4FXMzx+YdGt0KBfkAAFTTCi3Vj6CfTNVCC/8CLIbusQz2CvK0BL2aB0bmH
TBiD7hwiFp433ZfNftF02QOaQF13xmmjOuobeFcVdXvzZW+Y/acbvZMbrsBPn2FM
EhSdQ1+mJTPoZmzQ99gaVksz/gfmh8eG3dTC2AmbVEXBDxQHj7HtCUo7EpZeQWbA
5mkHb8Xl0QC3UDLFmAmlRVoVw+CgeK06n9jyl3QJJ/oy9wI0oREitxuAo9wdT4RJ
99dbtEvGQczdrj6Kuvd5WSw9qyyaok+nl8CxTo0aMcglWRKcY/qSUXD+LVjcEck2
2GV99OoZVMufuZIwyaxa1iSee8GtqJ711EZ/50pxZhMVHbjCpO93k+484Sb4HMN4
07dU2xRG88cET9XoNKkoR+wrrpRIDblHjEGrutt0hLWcFTDCrd52LqLXiQCQWi8J
l/PzCY+XDvI4HuSFMn2r1vqaqJlyiRXAzGoyl4l0UU7pRrLmUBZBB7OuLiowp72a
9dmsbupaOLT+IqbIVcG9bT8ElKmqqtO0jqE2DhaESi0NgJxPADdIiN5C0cOAksbZ
Oq8I8QM9NT7P+e1zX69qLR8ZlVaAUINg2u2f+nw0TatWEwa9LzTqEWz4VVNz7FIi
kO+v8agLzpdbkCG9lj8S1gOwcfl6r7wclxbdLiThlglWWBMPnhDxaBBNhV9AWj2b
urB2w2bkOgUcfCjraXg/mydVWA782xP2+F7jg3JKhiX768It+pl5M+te6aZePICu
rXXeaqW+TgAflZG4ZmImcOpFnELW5doqwcFDsb0fk7tdulU0UColB7TbcfPoxOPm
gWCZvepFCrkLsvV2QCYWiS56VX7VkrRZUPZD92RvPU4eEC7ty+m+jDzqYR4tY1QI
DFBc10vXzOoXklzyUcIGAabNrwfC7HCTfA2HsNcQjGa8dCnaA0N3BuSZS3mIKnkO
wxR4Y4oGG3ekIVs7lTy4hhCbQ9puibMGCtBAxPiwfCoGpeTqQU8SXWuoKCiXTJxO
9Ewwm2leiGxPdeOiH3sz36zFXY0XuQ/sBTBj15pRB9os+lS6HZ2YycLMAPgINK34
RxvhxiXjzn7/7fFXtfGckdxoZECmaeUOK7h9PhG4RyvCjV/yhMp3aai5n1lQTdd7
CM12mAF9lJfkDb8Fz3RiQjL6TnQoWdlWgqbrGCm2dhkQvct+lZohB0Obpq3Rq+AL
mpMDmkEZmHuwytPzW8GemVhfxxP0eomQPwRa+vcKEBtLpC3pMsGc95cohWDUu7iF
xNWQ6kZt4E+mu66n862zFxUa1mbVoIEAeZETGgHLDImv/hsBZffOscKFgQPLNJ1q
HRGSvOh0eye/mugUofgfDQ+Fj2SMR6qI3h/gfMhtygTTz4kHNeql8HYjWNL7cOfc
fRhw7w6IqSbsqZFcx2bMgLlqCs172pS+UppNEXYdgz8PblY49u3Ns6P6PHABi1fA
Ws8ZK1RcI+hPamKCdB2iP8S5ov7zoqk/AYJOPmtzy5yNZx60/AKcwiLwHfXktUEl
LkQMMqU9cIgfL0ipMS9hBfGA5ErfOwWZPUqHldBXuzgUU8FPCZQ+kqfg37elBWsc
Mgko8itGIkSNm74vB9NiBIFaASmJJlitgpL0F2FC+Ca96LZ/Kpb0LkC1W5WyjJag
6+K3UEVi0eD5DtjecsNDYSot5xR1X8g5fk7bQdbfi5X2E5JD3MKb57jYb/xXW3o9
5atlaDjsYJca3ad+3pOL7uyrqNU5R0sQjztUuAg4HuVVgmAuAAO29Xig6WlmO8+A
LBi2HQi3Pa+3X9mo0DmrTQy2bZfPajgmuKuxh0dMez3GSuX7Ja4Vxj8zMailQlB7
dJgo8tiBt3DQjrLTLy5TZI32ORqeqCfE4VmGw6QwIRBPOzDpk2A1XziNQHtJ7/Oj
010vrF9FnqLFtej79V/FN8OoDyFj9GKZkxfXgUAqJ1aI6gCpYioy3rM8Xdwmc5Lr
dJ3PJVyNTKp+jpJBRmVeMCEo22sWlo4QDAMSv2kfzk+iBFrdz6SgsNDdlJnqdBsP
JDbLeBfNNxd/wosATlVBEiTef0MQNrKdbnTQSoAjnuo3HtbUL9X+612wyFvUf64S
YDikSFbdE0aOCi9i1l0ALSptxuWDn8/dzb6RN5UZ0OZfxkpCdC4/6ZQwl1pIkyo4
rmHEy1AehvjqPzUOMEyaV4j0s7vxWc/5YoXTN3GFHkCVy/tqVgMoBHlfD55qrB5y
PbcvwjQSbOYDADMCeOVwNUgHgEwLFuAGjEXP8Kv3p6/c49Rnwm/hvifRw2MD4twy
fa63KWXCnGHrZG69aDGxuJp/KGYEsPMt04TsJQJ5qNLTEeSGcB3Wdo926FpLlN5M
0MBepLYBSI4967XXiQs5LxRB8L7kaLTVb/tN2bLVGzEdm2PqE8vaOi0iK7PYutk9
1P79Vnk9+dLPFAZkWUjmeAnLjoqagvmBVw17jvY4ZHn9o//5aaPb/LxfeD2J00Oq
Dk3Yy34Zg1bb8vCO+eBmY9Z2jNOV8dstfAnRfukVmQDEkj1CvMc9AUGZ60VHxE4m
RisVV28VJE3grodup3KL9l8adeLdHW2/sDM+J/Z4Qx2rO1TXgUWV/LacrFVvw8xf
+1swI0KYOpKMqJyK9hzxSJQcEB4z/2PDyR21jMkUN8Hq3XyuN6SGAkNTd8E1P0nm
STy5N1potBTKeZ3vH9Afeygb9FITZGZa5/tSfFoOUvA3fpcdLNyUJ6sMSet5iON9
J6LtfrAR0CVVTK8zAYcPA5x4fqGm5oA24T1U8faZLoGtONn+Blns3uce0zjMd35J
fw3RTU9HewFaZvOXCv+Hk2JygdWkHraAM5KTOp26QntUZLAzF+GJiWz3w1XUnQk4
bw30oTUmB587qZ72Yo4gQWfj7qOLjjDwAlfTu3SBGiR8OrI3mLwMx3r2lBL09YOy
t/atnrFBX4+l7KqssI2evOT9NZZNAcHmheSuZO3oDZUCcQy3NfRbfNZoMgo6rQxN
CaG86bqzqjFrAYZwt99Kjmltj0yOBo/zRMthg0aSzAYWsM8XzO5t+8wBAhR4b0GQ
LB/OeC+bZEKhnqAFWr08IOGeZyMusHYzs4tUru/68Sy2Iv7uovT5sT+hIl2lgUM9
dYU0P35Yvdy1fF3znNbejJOHWeDttl8WMbRRPRShxjJspsXXOYLYo7998tBI3qzP
Ip2Ip+uWMmmjGhn/x+KYK1fEGnmFiOhly1dTDMo7eo+helqc3QQoYxOTAAGNk2Uc
/PxAmagSrLiZRVbGRSk1HrRuVDqzM7z05/N8+U4fzFkoKsp7wOtyfafd+IzVhRKb
x6Jun0LLS2M1uj4VXkJCkgtLOMHzazpI2jz0d5t/nnGzsKz1jhNoe/XSly2jtKq+
jB50pMX+qOrbXhrJow5Mp+DNuzu3yUu/cGyxqNNR7KR6tWTGqv2qEeF6re3zaO4y
JRwIqQBmtfHwnZznaH9/t/uWsB9fYI4HT9iWJdszzCqZKD7OxnqB3Hs3XFRd0ltN
iKZP/mqKTI6H/vW5nyke/b9GkkHjedKtY7JUAU8bnA9w2IYXIKXMp0F7I7cu+H0m
Ee+nZoo/yMNIzVF4LUu6mdZ6gbLNIfMDJtIHSm+OWIsrC3ea4QFp7LxuPHmaW30k
ujhxovloCPJG1EFmn8sHfn2CvxfDCBvDVo3WMWI2Hw32tFEI2/9ZdTyGH2ceEYTX
tBNEW7NZY2JhrwKNDYQDiNij0cdZDPrJ5y/P0bFL3BXPir/trjjdSPJJLtyEmRKE
MH8i1veKp9ozpdClhGLYNjOR9zi5y0nQR9QO4S7CCAgrQ+HrDmf0miwtX3si/Hrf
zV9Gda/bF8MesU2hYCpc/Zjksx+73Fd1nSDYr4iPbTV1NzyNrsBSa+RL9yqMRN1b
7SVGdQXGrKRsg0jW7V4jAjWIn4xtbyX3t7CcYaIS93PfhzRJ37U8eid11BBYF2Xp
0BcfOEx9W8imZNiITbQnKQzp+3qEwPLOif9RRSW3ficPV2ZeuB7bTj+Y6L1NLuRE
z/SWfXUHHD9VAmAuxkwvpqbvD12LcKq2karGG9vYjRCEi7BnBOoxfawE3jA1gdZV
tMDdsKUCIqDbyO0cc7lPzkGQ1WS15AO7eiOGL6luWD4PRNeru06FdWxzEjuBjPid
+b+Do/i0KiLjabuykpBozoDLZObHe/GJ+pklxt3xAZXQUMZ5M4s5pTd3nu6OsD82
Ax87odJdk1NGktZPWsm3kINcI1km+Pohx0xc4I2Dmhx5M+ox25OSPt74Op4kJFEA
bFTTmUWmy8LFVnahey4UBP1dt6YW6Lui210j5WxnsUfQE3G2auX10bJmEB38SI0J
DQHeCgoX3iYDe2osGG/ePsQ5Jb37weE8mjWSUJ7axSxw6qdKKKhoaUIRiBza/PLP
ulzKkk5CZ62MLsgMrF5i5hblwAyWs7b63/v6lbd93AR+D/D3Tc1dHxbZDVYFGhE7
RRIeF9Ynn0rolyMElFAiU6L5ke3DH/eSvD7O0Fe9yrJ6Qms2XGPcJgsVgEpoGvks
r5bGc55vwBLYPl4TrIPviie8J0tSKlPN6YL/VHzhUtAEUquYNrdxLG6aNXUxjhdg
tYMD37I6DerLd0zfLM/Pw8AnK2WrMUaFjIukbuTBTt6umzywmDTbfnldb7TpEvmz
Dro+QUuQ28Iu/KhZeu0PP9Q/+sHnj8Aid0QJIXpvQjaSUToU5TlRu8q2tzeIAq9P
CU3VrUerDiL0nObdS4Y4oI3TlSCocDgC/0MmaDjKJhEg12I0Wkom4aEm/Zv31Tam
Clz9lD63AewvAj9pMzoH7jxJ0UXhNZKCyP+8JnsYlDVMG2TFd8wK8HypW5h/xSvS
kZwi4n+rmH0wK20TajLp8DZvYK7Dj4LTQcyzMGXr9Cti0jGhj7pcTMHohBK1uMcj
y1Q+I0xctel5rjpfov3bklI3/eKPcNyx6dp3tzuXXDg5vRss60LU5XtNAwtFd6if
q7SnNiVxcghGoiI0xEHaaYmm0J1Ugg60h3jxE/rDuv1cUgT4aw1a6C7w6xQHZK7L
cjeBG1DheSLNQMkd5elG7Y/GdWR48SvZsVZi4bpO3KYvDzrRCMZq1QtMJntqbf8s
ZhKhVv4P/Eul5lEEMw8PXxXKXnU1JPGegfHkL5mN9tDc+EJ8jyI02dSSj0xLwEHq
zgARWN/vtEadR+lLNiTUH9RhIrGkoIl5C0CMJKfd3ZZ/6PwsAH6ZlzOKVh/JxINm
PaOz/tINzw00vZ6xFOVspvFVCBtPhy/g2KzTbxMQvm9dj66k7I0uiQO574VvHzW8
RZNBqE4W5ozmMjnb+OH6d40HsfDTazTi9OMli7BDp0o2IUkE8sBS+9d7qc+ogJr6
1H8+RLYWY1lQq5fYU87/HHQ67sFE9KlCQGCbVpgL7LUtBx3XTQ/im7Q6aUkzYCZL
RD7dsE5RGDAy5Hv10SstslE3XbzJxtK9a6+SjtiqFWG3Od7RhUx/tlHzrwAvvpl1
YkugOQjA02KtyHPZ+MwW/QsFIlD22kUygCEu50Dz8b0PueB/bQSyaQD2v7siILF0
A/0Ez97OUvZf1WjgnUz2TNlyu1KaXaAp7751Timz3j1x9+YLJ8LEqx5clWazUmSV
UGV2x2hUZXwEFOiaBUC053JEn34TF/hH/9dfx6YWLEsZboIxd/n6mRSRinxDfjEN
d1Eh5tVxwg/V61hymb9DKwV/uK+I2suZskSxK/rCgARuuwnYPVtJ3mLlZ2yxzNYU
6Vl6QMnhzYf4EoorCpEhTVMQdi9toPnTgz85NsvyRiuhywiwD/W2RcD6G3TBBS7V
l2ioHdTCMnZjNaXzS/trGd+RnFL1NP8adYR4oXGY4scrEHGG2kF8RJoM0BoR04I3
yY1a3CTxmiSBQWpqoNQ/19OZzz5Y2ZPBh198dorkzXdwnpvpbojqq02djBOzcOt7
6Sn6aysfxxUO9uxXlSjTEez3W3qxqdecgZzGtWEKpGlflp0IhEezCM+K+5fXBKfL
6olrwsaOuFbn5aaEq83WV7IzbwYcNkHzyT1i/lQxIGhUIe+8kqCc2yV41fJDR59g
s6FL9mmUDhwdek+CzCcWl3qOLc7uFLnVkJ8EjBLUC/zz9nODUoMj27TM/9WWztSv
t0WsyRdMENWRpRfetiboqU8pbv2kXoi4Hx4R8Td0qTKH1dlG7THKHWBERJIdz8Q3
DB7j3P22y+LSETgog4Pr61KrNaYVlL+dd4k5Vv18C2yH5wUPFhJmeHBB5DlJiEja
5WTOaNOWRYmtPWiR707FSK9Te8fZ9jTvrq18sLV1mQEkzL/RGjNWtWL76wgOs86o
SCXYteeValAsNnV7wZ2KGh8oJtvkKa10m1sPuMqZ1QgFFY/jJyTWrj2X1AbUhnkw
UxTziRwu//2DFMN+5ErxocsT5/0MdWIfmt80yoB/aABJEjmelqOv7GeWwXQNEB+r
pXLY5ocTL4C6BnEKG6RQbIXYwajOpur5SD2LFGN+QYdx98l5jUim4+K2IAPFCimz
T41gsqGADKpk/AuCvI8JZN0aEeWwfNOoqSg/7cy//UYopa6gt4Udm3/swCCWaT94
E10Lhi0Ncr0FvUF5ZbQd8nY39+NtNyMR0GvPEm0nGI1/Atuv4XflZgk6bx4OQnCr
afaA8yDLM08ZE3eptiHplQpoP3nwMRcrndlQhWUy0LPrYOxFYVUOOeHRpOAzlSAz
xuTlGlo1eWc+7mfR1+bAYNhjYfPYIs9Dxpz3Y50bR9lCSWF2q0VZQTGotKwY11jX
W6kcpKqUCRAt8t+BO/wP5/oeATmGyEtktYUHZDGrwatsGd+bhU6AJ2kOoujsX3CM
nXMS+qNa2K+v0IyruMgQCoQpm/uqC/WDKoDa57tBCrBx5j5fcSwXAnEXe6yJUA8k
EOXj6g4gaIW1+QJLdjPFd1ILr5Egd5qf9p3Sp1BWquFYPVSQU/cF6qAofRmFZT9o
9PgsNcOLhQ6o6CpK5MAik10SPiQvbuHtmDVCMw/qZKo89qbudqlLqQmHaEPPACV0
Cn+REXLxVQNtCo4by5u56YbHfFXKlPZz1UCq6vzhrsQBst5r7VU07esKmyfYEbyd
jEH41y2Iow2nZfw0MphAwgQt4Jd0o4PWe+ujuQsBX+TBrig70yiEEsr+KH/uTpp0
cJMMNg33RTLU7TyeSTh3CImRRIrTV8pbRgm5FWDubXF+28oMAMZLw0QY51onCBuJ
aZPzLfjJBKSXQC78MxXqj0o/HznZtv7F5mByQYK8xyTBz8sFtEoqiisvtpoqyKDj
7bVbrmSoqYrLRFYByb++ii4agVG6gWCT0/TYKCrDd28eElQEZ9Y1DzLGxceX45xp
d6o6czMdkqF8zyleWtDZMS8qlJ7LGjF14iwJIhBazjssHCId8X9QQICTba8IMTI2
XzKUgGli4ie20wcenLkR+07JR/Qz9GrkYc9CbEIpcPkK5XyqZ0oqX1gUJEAUwpDi
oZ3UuwWn3YsrpYOtNzF3NqJrOyp0ImzWFKnd4c3k7O9HG2yqs1Ee2c6lgAR7DaVD
FG2whdHLhfahsBam+Ki1GXcSN9fyINti09Ah8eZeXbjt3tFzSY0cP7SjPvTHbRoH
fC8JR75rmyPP1ox9veDhSjsoSyWgZB1Nx805AW2qBeN11wKB8ilI9j4OES2a2zKo
h/t0fP0T2PnI4EmX2voEhRw3/fLjBuLXE9gYcjPCfpawxg9HOWuYQI6VBY766qsQ
0q9/Wc/HqUQIlDTbu96HclxXa7Txu+o3O77PowwaIjf32g/KF7AleD7vH4YOqUGS
ACU5/osbYRmm9mcNRV6EQtsWoelp952w3dDEz4xeAtg2HcgmYFrm9ndp9q4+MR+b
dre6ioWCdDxv8cUt3ekzOW0H0uQq8sqBIdJTyxfr+gFsjGYtH8htfLgOMQvzx1nu
bNYlvlUcHnkFpkRb/yNNc3U8FKwrVNvCGSjymADcxWHG5kiGRk0AImZ34alzItT8
7F5TXQKOMy+TSsYdOMolESoL+jHYH70srtLn0FRDF/SHtxGWXBc7aksBjlHEBCGY
sJTePiecAg+SweNQFuoMik0Y9G5HZoUCqMsRu2x3vXm6tq/7nmiyPaMMHLUzOK3M
mD4es0P41SHNzbPwcw2a/67b+Eno7SfeL2dbkD0dA5UoyTaX+ep19JGzKAqLIGBm
3jy2tGOosBzDdDI4JME8VYMKCGd7dcbIcn5yePyBfrdv9Ox1q8FRcHgszfZ8lxZA
8rFdNefl5R5WbwdFC/4DpPPNdFbBmB0UPll4d96IQ4SDbX5QZgR9XpwKswhXHZmB
GmkKDe/zqwcpYXm/V5Mxf1BH3/BQfzwmDyItA6r3z/Yu5myHe9LwenXK08rgupyV
Ri+il85H4q17zpotdAV8a3Ja/ZE0cQSCxniDMNJ6IOQr+PKhUI/MzBXKejjLJBmL
l5xzL8FshOOJw+NisjdhRH4i9KgyLzAFMdWWhVGwUI1lZr5opMJ7hcF09eHhAYXe
4FtVyczAPYsRimB5HPxM+t86p2YTT1UsVH7oqoyrVrN0jmKPNIKA6bTLy3cE9Yk3
H47xvyzxKqXddPQ4Y6h8xgQl1IsqDv4m0YBAjDYYEwjJIDn7HvEVTUC4X61waODU
ULQpqhG4BvsEh/dzpYcmrf8gRn7Xe9ZgxHTglxCAtKFMt+dHBit0v+fmFMpoWM/A
qvj5W0poUuCvYy4XaAOmAJBOwd6WdgvodIGTMxYDX5OHptmYkZmJFCjysYZOuAit
Fi6jSUPgxrQm7jEZgyYYof2FXnlvFLHTWOgWEw+V74KJG9QYeVVethPpl2IyFXxr
5+8n2jt6pw3gVXpjQ+1karFkcpendTz9WljQ4smkJVL/hxaNlZrWvkM//o4kzQas
kSSyYg14cWDFFdbgY+UWN37XdprPB+971VUpIBd0cM7zZmu2pkd8VJyThFEhztCl
zjoMpfMEyf4w6u0eupCzRSlm24U/2egf9sn+NG0/RXJyX2zil+vxwFBI+CXPYOZ6
kIky1RMhkYD15KpCkDjzSjsoGI9bseMK/RBEcZwmuNd2Jq1qiZfR1Er/73EBLFeh
Blvs6DzBFkSwr0gGaTasJhisy1a+bDOqjnSPTTaWiCwymLWhjI6/Hw9v5s4QvH7v
A78BKovmaW0QW/JIdxrokVvsqF7irzclV+AfteFGgcj+kh4tBkJz7zbI3A8nsuhx
zWWhxsjUIyS2+6AmkLZRZuEgQk+8nQ3K0tDEGFFEIpuUGkuCBTyK/YGvW/qxSNJ2
MWAB9y5gYH31GUKEUpl/Hn770NbCDgnzYOzOGM9u+1NXenAv7/SJB/YrMO/XGMp1
E18++jLiTYWD68LEnl8VoIQ8iooQaLv7YzWBfuQhns250kHlO+Fck5dkp8OD7YLl
niotqxMyBOZpUp8+lEEdjdnf2GAqH91S7QRTCvruJuHHg1rLEQn5qO2XXe2rk9Gd
mSnVuixTVDUv6zZkPmSBNMEKaYOssFSXWFhtrBN8zSzDNDYtt/tNg6gxOPPSHnSV
tZZC9WhKX3PGIOpcjUv5QEjX3AFT9tuSFYuVIi98l1poyMyFw4/cqmbbw3YT90oL
rzPXkBrwrfhvk1SJmH1ttH/zywFxXdU733q/I1YV4uT82Z469b+n5ayuG/56/Q/S
DHZ/1QiYEGv8mLHAss/M7JS/C1ck/thKsnJfTXPvmFbUiDoQzKKKx5okeupHMMhE
GrIRR285JL7bJPFSeB5DKNtjL3MOTFPziVWobFyATMzOEsvD8jevJa/rFO6g6Rlv
bBXS+/kX67b+281Pw4EfhWs7V6oSYA4dzppoTw/ocZurrJ0MvE6zAhEL5wXRmQGN
8SYIKrrRv6dRF9yW5kXtPeyI8Lzzuro1t7Z+mg9lMw12/NQKj9U4jBgZgB8PPJP9
LuYP+fiRPAxnqOYn4dRz084MQrLErK9iqnapzsjbNQ6I77v1dYqInKKISw0UHzYG
NTZ4o0wfBN4SYD5V6beaEq7uO2W/S8/5H2ZGAWQ5/CqwWKpsoZY7rZp1LP4TSpjj
UTpHtp0qLktVur8pwr+BiSh+xoTSJEZ9SPrRn0m5c0ByGuOSwFCz1IHgFQDFADf1
f+klG/qS0oSc5c0IFydj/UquIsN8GXEsFR/qCLr9T0jZ4Bfpj4bvgJXEceoxqZHr
1acjRJM1MYMVUYyFbHbP2/bFsBhPo9VSgHyIqYBLAFPqhQr6WCphsLmEhUYt3bhC
kb1GosgkDaTg/rIHYFPf8LzSoh3TpsPwQAUPcwJp857cELVfeUPaLp6zKBnV900I
sYKodTr7S/x3ftgE4ZmWwJIQVJd+CpApRL94V1EPN5YJyC/djKcSCyx0F9X1dRiZ
aHLrRXMFdVz9FTmKz5xUjKs8Y09v7zVi9Woo3qqsrFv0TVb79Zjrclq1kZvFsz+x
LPBuEOYQ4qWp+pfjFppJyQWtDn4b/ZSWqUv3A8ekZYsJzY1agvDGHJugsr3plP95
umSt00yYNzMOMrju/B68ndRSr8fV2DXVkJILhqJKj6c87P7oPCKVnL6LUPLCx8KF
GkaD95znWu9n7mNFFHTQydY000N8whiMHio15BsuV8Kgc/z7iZSnjChMvTc9d57F
iIuismLsLTXaMhWBQjBfEe8EplalMD3pPcdpT16bUrk1//Y6fhABFIlzzFC9gCeo
eRb4PrzxSHXTLQ0GGmtx8tD4Hd7sBTe54jEa8rsddN4G5sVbEHxTb63uqt0yqkVc
iJkqIVPg8pULQhnsF2QW5oxNx2KI30QaIJRKnWeyLSSCQFTTWSvO08YxOiuHCWhS
thWxM8aHEoSJmrIAGk99+E/+9hDaJiJBmKsi5w2LVLLIfNh5eAYhBNWJm6HtiLf3
z+uKfE/LL+rubj0Akdjmuhsjz0nwRZWrLGHFtDyuyPQIczWAFDGn/9HJL2lhCksS
melAR3TG8U4rtG5ZEwSVW2MgnMTg5fHltlFm0S3O+vOP3hzsC6pfg6h6UtbZWp+v
KVwsPKf11X1Sn0u+2Yc04EbaBDuRjYvmFp5J3G4wLjwjol1ZSFBNM3Di/rKu3Jsn
zLiZkgXzmFhx18bcnhlXQERyuSprxw1BYNm4fp6VYGAeIDRMafPmZXp+hqegNISe
7FvSo6CHIgTxQEut2qg4D+stfKg46SScs9Pf5S6Znx3IQSLGsX7YPabzude8CiO+
dchsj7hO+0YbFo5d4y/+BEGUayK5aoDggl9try44ypwfnztFuxyLfaIhGKW0NUU3
Ib7s2g1EROkNGskE8vmaktvAsQttiajeQ7aAD6WJmnRORcGu0am9qf9nbKra06nn
J4v6O5bwBafNzAvM5j6E7lR+V286L9uE1zOG5i8anj8nr6XAEMy9kiPg9moXkBq+
IsjjQuPJHvPSCcxw5C5ph9J+u87oS96+GSJhgjFFdP0oRGpv8Yx1uYmZ7eqsMCbR
108PMmOrHVfHXgnUu+fdmAUvl3TIQedqDTg+WVrSVgP5cgPlD5ny/6JkktNPAdz1
nAvDGiR5l4q5bMoTr8lbikpi/io1dUvsaaAKfMQslLFq0FqfZzh970xex1GbdoUD
tN+g26zON34bwSYA3DzkCSpEmfiQVDSfdJJo6wVUCltkOF9TPTmKuiZmBUFotpQg
cIyLooWtCO7xM/JRTfJ5AV9Iltv85sG2MrkEdi35yJpGXe/tKoT5kwkPpanXJH8s
y8+lzOGMryPS6uIJqzBxxxkXHg2wrn0I3gAkL70+ujMvbtuDeDaRbDxwKXO/ZXkO
wG1b+h5riWYRvk09Qmn8nblExCEtHIscsfY+lZJTEOmtP40amSfj0VH2bop6fj4R
MIOAC9QibxHxQBDxvPKwYkBupdP9MUMCMZzVJQn/KCudMElKK4Cgxqu27BFTTZdA
YRd7+ZdP2n7rEqYG/mSNox1k5rcEUiKVnB+Y5PkRu56u7uLCLGER3BIpowI0TjSb
6UrheEdR07UOUCsQaFec9y40ZQIU3ItPX8KFzm7Yl8Hr4Ky1zsDfSvL3GIoJIhr/
LxPW9l4OinGhg1vPOObmahWSKk8+Reaem3CkrnByXK7thyML1zeBJAdajTmbFgzX
lEdQAPbLthKosN3AHp0Avmm01cvO9iKqYEcKiJC1pH5dPx5fgQk3V4kCy3bLGsgS
qAigRVrR1dkiYXiYoRgHPjFfIaIvO9JkmCspZRScjJxvAo7uWpoMf2LtJkrPjBIj
eHfxF3eyD2JTjLwxc/QvFDogvp0EbCNJinnB1etwr5NQo7dsgnWA1DPrKYoxVY26
dDix87d3PTiGtV2yWkIpKyfniKNZgLuFSl2hG1kjTo9uSbE0TsOSzyA39Std4zc8
MjpJCHrumJgNndAca+MGYLt9rWkeY08TvjKWt0QXaWrFWY3tfQt+27kcwxnU5yvI
FouAFEoouh35faVe3fSxjRxDeiDTWlc1iE/tj++bj7N2eCIkhYSOOcOE8eA8OEYP
EEdfEpNVYxgUA5h+8dSI6PhG/yaPIMAzgNeskARtZLHt+M5pZAQHtJ4LhTENFZPh
R8TNCeCZ9EQ2q+ZxOC2lsLq+pAUiOlvSZZJmpIM9ABfle/3rxTF7yAwVYN9JsTF9
SnS8frXpiDETIzlLl92WRac3E+S0YE/nxzto84b3G8II539LrjuRhS24I14ZyWu6
SSI4/VBJBPfq4zXe4N4YkBxBUwlQB9cJ857ypDX/urSo6RxVHjhpVNzkEU3vLhwS
8gXXdtPogeP8hpCeJDAPPiUhezUlkVujZRgYe5PiE8r6moVTAmatYfsxmkzcRssT
/reJleQFnXOFZ9Da1gbikIfA118HcXHf4RhwTLT0dlR4IXNLd6Buov4izdPykiXt
vKjL34rZ8h6428jKQmH5DAFKDfIi888XliQf5Jm6ZBZYSEev28xKvjIp1gPgXzhK
z5z42dqIyzOX6MRKjIOn5BDvSTXw0yhpWOi52F/6PRNAGJXzw5NRzVnXwnAeZllv
iZNW5UH8J5K6GwbeJGKr8e9bUqqrjEvPk3He9qGzh2abCBupU1TrUesJf7PDFo+Z
j1XocWkg1he2duxp1aKLpT+eVUUdwIjVHw7rvbl1gGvqFcH7dPyaJpA/ElNTbko/
4o1cNdW8EsW210MVAIzR6eUKAQRrAoT6sdeDQ9XcH8alJwJVgJN8Kl2maaWldCtE
NHY8PndzMa4j7GRMnWMfBLmHZa3hwOZh8WvPNTSxghovss/cF3EncB+aeqV2xVmB
/ldan2O0CaLjaq8MB816HeRw6jUWYxN//KOKPWHeeRD8+IUqipqN3kd7z22FTqtZ
EFBL1sr8GEXk7s5bo/d5PX2gsUTFaZ9ae5ihoKr5YcL/k5o+FNfaet7TOX1FbOvC
w9Mmcq4dRbdejDm6PGt9TMWIIlj7gJpnLcioZZRF8OmUvtkx1gV+Qk4lQPZVxg+w
Q8MXD0wxUBOXi00moO47uZjnxz1KGN1GW8OUqLFWNF4saWrNZJhptfKjcmUzdI56
P8jUMDdZAefYtfXUoxDyp/eQfJwvsH0yaLqcod/pwU1GToHEAoM3xwYdSH0hKLUl
bRtAibG9T3u5YQMwmGj3GxeBVigjw9kMHsH3CDxUjlA3grJE9/87vQ9qFeYJbohs
y1tL02IzeFB2JdI1updvdGQWWvqwiu0wLoUL0WdRAz0lKaXyi1EhSL/eSLIEyamQ
nv4/iNyAVq5tfBlEN1LuNSkfR0/0weT3S7w1f4qLduYGsJDPeH+P7QKq/aAicBia
hs7lg3nTOlWQ93v+X5eGZUvvbDBxWj9fbAfYj0bXR8DAYvAtqO9rOX9+rJkoHDFd
I8sShwmJxhei7LmJkBWu3mNvW5A+DCN4kpPACIvQolwAmypT3heSq9XS5d6H5NBg
3yQ/loq6cE+J8pZkbc877rDd2gR8gLx5hg8uJQQPQCEk51/vZ6odCXDq/hp0XhTo
jn56vZZ+AKQ6LeeJ3fQNYTPpvc5MEG/a8BwlZGptO8vlevq23XJ8u95xWMMXEP0N
NhcIi/X0FBr/5vq/+sAJStTmHmiIiZNQV+uoVY6ZixDaOSWg2+HYL+o2zQhPuS+E
Xg2nu3bYg7aQ/6okmnqvSBIJVbXBEdeZOqf9jikFnSGGcCLIGH3TO1za5TRnDVZX
PyuYNj31oLWwZY4wA3S3F6850Kt5skhgyL8RlVmdFciDBUDp51uRTj/Gfopfdd+6
WTDEV2i1Zvl9SPuZ5PkE9obHKldkkP7bppou/jQ6lxAwtZs6E9HWWbmyFeyf9o6o
rnAM30c/nnsT1qi/OcFhiKMkKQfXOH3gEqkhXvRnHf5XU8wyjtVE0DFUVVlO/z2C
nXtX2PRL1zUmy28roBRWe+4kl+Gb0bL8FEkKv0j+GvtI8w2q1x5lNDan7a1C6FtT
nOJoPhlWUanxILvmUo/bRv3XedmBRtzarLc96x5QPq96tfFgPaapyPT7HHPUMieI
YZlLIcMvM3DhqeLp1tJjnPsLShBk80CZqPRDPXZbZSMYAJ7bIW6AbBqZyMofBJTt
x6atTtxHyk1sC62L/XBNElxnUBaerylWNZdng3cSUvRqwm3tS6QSV85pLMOeq7EH
uoz8X4ux+XJ7r1vkesB3Nq+q6F763djUYOBnbzhK0uxq0M/LNq6FXFZivuzXekfG
gQ/uUmnyXzad3gH1lPlNpShDCLItKRpR4OU+d/+D2kLKl53u9Zh0ll5kxcf4e5MK
GbXJRXKz3qH3BbM/Ofi7U3Ec9z5vKcT+ugDikPUxxqeNDw2g19noDS7d6Y+lGQpg
DzUbC8tK7E/JshaVJ8kwIcAo3Eru0oN8IhJOrLaxuICEPL9H6WM+HHV98cyp3rKO
KsJYsyT9sBQg2oxWL2DSS70tV4r27Wt7cjFpK7dlwvyUjMjAO8ulyAnWtBljBJwH
Q4cA3ZO6nPgJCnd68xTsrfFmAVIgvNhyLj5d20Z9tAzl1X9voYBkIKfnZJVPzBCi
9C7Buf2bXk5sj5fyHn95BvK+aL/YMssVMSazKEwsDXLqQ2wrdPxH1ZJD9bB07wdP
KxGWZrwr61YvezIK3U8is2aaB8A6pBf/bheBWw77k5iq++3/4nYuUbFQQbNQSmob
DEZUM+n5uGimwLrrI6pvhXazTF4Rx6dD/zD/u4iS4cv5KsLiJIIR5jeRVdnP8G9f
gE83HY3iyeosO0x1qijTA0LvHSfIkJoCUtCPLptnkzW/40+iLwBqTuSj0v/Z7J49
yDCGgp6Wf120OkbBGbAT+LXNKjROWBv0agB4L8+alHi9UazRsf//302zVPXGVUSx
LMr6+oKGelhbXcKH483iTplmWZxvP+k/zgCslb3Rovs2UVb4+Htath4lxcpuMggF
fY4ujpqCL29Ekvj6JUf9TnSjMWexmgANjb60V3G2DqHos+VFXcfMQUeLRg1uE7i4
sanKyVMClWIJv7grA89y7LIIcDiz0RwqD8/yr3LKhSlRzECuLmUWhEVUy6BrXfo/
P9jYf6kfQDOptezsWXW0fxPAsJM5MUhz6hz4ubnSX4Z84wZ8B/AQQWlqEC7/ezBG
tZUOgkS0EdcYbh/HmIWkJHrlmTQ4epAM9YzS3qBlqWUqBhIHAJKTtr2HJVY/Axs4
u5CL00wEFEtL6OBMyoqxhiUD9dsLxq225WD6QLhlnxirB0S2jImRZALexzkaR8DK
wSeZ+s4f2yQNE/gnA2gYWdLgLl0hziMT4zh7ncUeY5HTJfR2aWmT/8x+fWR4+Ig8
sK4RsqxNFcvdhtAniMcIi/pLmiPklt053RapG95/RerzGQ3zuwg1SYGmlvbAsjir
+GNW+DMOH9ziQ7QO9JrZc35qH7dGcPZmK+A1npWta8QeF+J0ZCtiewa5cntRfZcq
Qn1B9VvTQbWjtPFSWc8X01HvMKgrlkdhrl6h/6Oejm9cBrPqjDoYgM5KQ0GrdFgH
+mxVaJhTr8b8OQ9ijMBTXEoUE9wM6uWMFt3oYd7TbDyrKz3+OXoNEHNHFn588oPp
+Sr0F3sjekLgISrHPo5dY7gpeoA13wrTC3gt5YY3QjV+Udp9bZgUClUjTJZ76Gr+
w2++mLVj25JVLWUHD6WzvPKJ3oL7RZTSb6UuUFjzJzXTxb+jXXyhrEYKEs04ALf1
RZoqQSYwevsCRWIhyqPzkONMhPIyNGbDJhiz5xHeymb/yupc9hImHAxwYyWc7k6/
pMddhM6HhzaeJq+6abHbhD2CyPitdZDLkqi9yTXO7dxVaBj8BOIiPvJ49j0LUDS6
U6LBoa0oBwWO5lir3Bhzn4BAVoizwNK0gc/vKO8ekRA0RCjtjQYMzG+5Tv20dVXa
K5z6QHPwXmEl/zVc2JWMMc7+Athvrw/+VBjYMGJXoe4i/HEGIzFl9FT/f3qXi35r
Y0TMb3KlZZAyGkhDAiyiqRxcSJH32MBQ1v85eilLeNT8Dn4vxzDQ4TNbq9IORfc2
W/lpIXvMb6jwjE4jB8S4BQ2Dq99eZQrMdtxXkdf5zOyd0sO8465dH+1RhwE9V5B7
oY3qVnykqe8Vg+l1me3h1A/2GPJJ9Alm/2zsAYdN6SOtKrAMbVuzvcWRQ5EgHoJ1
426n/Vytjw9eSFHbvRTZpbxHaERL1C7xcbEezjMB15FsH/+/FRlWk7ZS3/QHXwKl
V9Uaj4rSzPS7dLkFmjXcie4BrtGgC3H7qTZYp8f+Bxr2rZjwXZ9cQBRvoA5f9F7/
eRm2UmPJt9uNVuzS26P4dUUWrm5GkvTiIgGhcmeiSgGXTinP7DT3Vr6s+jRF1s06
6Lpot2RULu9f8Kxs5BuVhi/dmSCZru9Aaz2UPmtyrpZTigsm5+fk53GTQaq0sIhq
mhVEUGSiqP+TFFd53IT59N4gHDaJd2GmJl9EtbfAw27+g2922UanwaKYsb89OoXV
cCwTM3juBrqkHlcCHkE70W4PnfCh7Z1ioxsl8htrYt1MKatgp5LhPCvV1hdVrqXp
af0EeihMEsGB3T4KN6so/eCM7Afttcx0m4kCUiQsCIhofLrVO4wTvsCM0OpctxPv
gbIdQKT82HfMw1T5V1DJYZhpqZtYltSElP9dmyHnEG4vbenJ4CbEufQrY7Tyy6Ht
uYcLlau+r/vv3UBveWIlXZJggEHXEAxCMO1jyeST49kOt11P+CjBzi1cuj4b8Dm7
IO5uAyyXebhLTYeFdyNBFEGSG8ZQN4MKXc0Yro3aR8UTlu7o1bWEAtK7UGYhuzxB
wnVRDpv/Cza5kxsoHWZyeP0ie8TWMTgaoku/ggVB08eaBku1MRYkqJIw6XKRugNi
u9YuHdF4qUwgmSrNR9hwhEQa5M9Njt9nNE0TxHggOi+tYNmmSR6idnWvS7QOzdnE
Zo/+HhbLDMZtcKGmcCCPOq2NPvLm9kIzTE6tb0ZKxu9A+8Ca6Qq9cnWw3Gg2mSlg
Uy9jE0tjrElLR70I/rYRbk1qHazf4vOCuAKV0YSXstEMi48QAe7jnfdF59+H7pjv
5lhN8ViyrDN6M5JS5H/d0bVB7XjpcWoNH260z5WuV6jpMDp/yqYTIDrdA8UIdVaL
cKAZI6d6ZJhrxAfgvVmJqdpIbGw9RhVA9vUJGA2icsZl7vu2FgikYexhyqv1QwA3
fKx515RtSJisja6mD9hNjVerK6v+FyIrBr6ykEci7ejH1VCW7mupC0dwYlxOTgpq
nO6o8yyT1BA0tgal2qhqZeFE4O4vv48dmauEgvDcrA45kJKk2gGt+PU7a1Vfatch
92DlVbjhaATM1ZYctYt8HbZvZhlL9wP1HNolgFG6YLtcGl68IIsX13uy7nXodEKq
XpeBVhNGnr0nBqQ+F+hvdV2DkKtQ6la/0V7/rlFHw2Ni2XIwpyIagEv4nae/J0oH
lWG2ru5gKFPjsRE2mR/hOtQ0j+9p80C35lKyYYeMLwdj5Fhjo47Rg3NuADeyQiqJ
iyqtdnZM92SdrzLY7IBHGJyvMPVoqVAYmBuHAGVIUly4zZLTofDVAs9wFxWwQLuE
Pdd8HCYKxDQzsQ2eRgx0ipr89Nwkak9HyPSoAqWESQ3axqCnJs14itjoXUJFdlo1
FKsC3he7fcL+WzZmM2m4um7XE7lY6DGlGIZCmtwT+Hpf8N8OfUC/uJF+C2SqQDzL
GyBH8RuVxi7S2dq515ziSD0Bhwnwo5wb7cKhPBwbIa5XEyOkeFb9vAmtsUAC5qNm
SDIDM1XlgtYMg6xqkMh4qPGJGcCVmQKTNTcl3fClCNPO6PafBXgXVzJX1mNHKPeZ
9FWkFle9bxBrX2wqrBjYJ0wEh0sfRmlmFYlFbdrWa8StYUMk7wjR4plNvWwVb5Sz
vGKS4AYXRTJ2yLmjAqVBRGm3w4hI3+JrftG6S2vd/HmrERaSso+istku3Xxnfp+S
z/wwns+pxZKO4Hdur86nbOs2GWJ1w7aWm4DQccOveQfsAD1yyxqrpqsw6TMg+qFf
UA7LSVB8YhSVIRgB2FNd9qq2S46Yn8TY29r1UjG5Xr6knfP0qbwGiLAd7pAlVrYg
HlHNc9QuTMScO6GmY0Woza2rkVolVZTTxzVR5PemQxc46dWwBUaiXZryeQLiPOds
mxpsbmqdxORLEumaskf7SkS9xigqBTJwzHmwbfCGgDVQVTXNKHmwWIy/w2uK32ka
2Cby3oTtojwXks4/ghZRolKyg8/NlZg3JsMyfCRGQW8SE1uG311bPaA4x0Thndqb
9/aqKciF/jX56xO9bDDoAhn99hOKtcB9t8v2UZr8fR/EYSbC0WNu+5VPB2Bwc/r/
/abfE7U1pPKdl94RdkiVWCY1Eqtqvp5dfL0cXTOpmZAm+ociaFaIfgQSW5N879Rg
C3K0/m67CyN5hCy/6gpmzbzqAjLzjwe6D8NTxfa7hmBl79VmcUm5pvd4NehgSM0T
DtJJJr1WBBS8AZuQa58zC89TfnO4Vd9Xue4W+hVJ4U6kYScf2JoQ73TCsUFsy6+a
5N8VKn2yRtLBYRtPTkf9BaEQQpp8ot6sxdEH/o56OtRYlR+V+CxYbiCf2ZeQvQBM
V8c0ctuBO8uCsyMB/uUFZgx08TTg2/TqYN9WlnG2jhUr5NdYrpnjZk699TLh3r2n
S7johz9Roh3T/E5oIDN6/w7syVUeCV6jTnNso1yFTNPMaZq/vEK9IdN8kr1ohnjy
TSEH5HveIenBrNoEsBFdp5H1EK76Jgo46QFflYZbzGPM0/+bZD61sRdPjI1Cywte
moREvcdpoxMbPd5LU+HwYyVa6gZx3Tgg4nHqZrlKyxVYTdgl73DLUQXD5fwlKupR
3f+WCdiwiBQ7n0kqyIb6ntpLyLABPU5s6tW2icN6Qem0qqsIx80YUBsT41yMoyni
zUY+uA+qYQp81sf7lM7e2N+4+d0TAT9P7iDQvEKy19ryXzb/mPZnmp7qmdlOXlER
Ib+UGWSbiHsNvodkqLCc9sbJE9d77H9e0Vcbqy9SllLv58daxAA0Jx30vYoAuCRx
BzCEhokyTtwWhmCnynIcw940ioHJm3NtnbfD3tMvPwl0LdfAnvXzxMgYkVaV1OCd
jahQOCkkqblYh0f9225ggzRXi2cnQ8TGJ9QcGb1ve1+WmtY02OAwlo3/EdsfS/0B
jtwcsLqoR9JkkpAnBHSNQ8HsKS7Er3gRvi73GsdPM6adbO7g6DV1CBiGep7/5yeI
H48FkUqsz2j8ICNCb4QmiWByKG/CpzeYq4f4xdmxiPzNRY3v0ubgi15/de2ReDQo
bnCiS+vUmR1U1UUY2ZwJ2RRHTW0LZSP2EilestVlGp5jQ+bm938d8dctqD7xxByb
e056iOT9IC9/nRqSUSdPrBEKQ2VvEkf4RIqTvClqGwjX/Bl+9cV/5wRSU+N+6Trt
N26JQGjRXfJU035A/rtN2jtJUPJc/v7/z+p1iMtm1A1vEZVKLmgS2IjgurEG6qM9
huK9UwhCkrgUBOnMOFtuipPgeNpBdb9HsScPrfGS7V+Nxh6oexwMyfjcH4kfudZM
E1raSnYscT71JQazgnBpmjOKju5/LuC1e1EMkBpsnoH/CAexs+/LlV6NFkgnLA4t
Hbq50zQ2hC52oNrBLCljo+910XwKklbZC+MT0rypOSfC8g3jy07UVTqvO2bd7KTO
7PjOCpYT7AG6z5KvY+9xbQ7l9awBNWC0WkFJ739/Ewp6DYhyJp9io2uorbU+iSZJ
UqkcjOGMcVxoIPjGFS2F2Whf7p182zlWIFP5NDqbaAiOBjml7ctvDxhXoxnzxxAh
I4hseu7G0teM7DB3JyTr2+TIUbhCgbrCwhoNNZ/XPN392Bl7dDOB31PfjYWAVWQS
YDVISKwGUJS4032HO6PA/FHpfhQ7lc/3ISVlGEGH9pWHe3AojXFn9W1pHlQQx/C/
Oy/2lIulwoiCyuXFxHQpyghaYy8zjd/1F55H3RygE+Nk2srsn9E4btfEuVB/FW/J
0r9uF/Fs36R1xlhbqldhLApUsm9EjoTqDtWwIOGQqxPbFoFHb0Z9hu7NGdnzR3WP
mmoaYMm31W9IXmknxTFSspwSf1vMek7vZCtTLbNNVX9CP+tHW8U/p7DsN7zLt9Yt
lG6/rEIb0H/3Rv6Vf0N7tK8PIQUchOsGV0a4zJxswjX60I/H0vLsNNbL4RL9i1g9
kx59oLZZWtljYkZGIDMYBnS9X38e7DHwXUc7D/5vFEIhDZpp/l+Z7Wl9iQMEKBMQ
qxC+qtFyPhRGaKz/X3InM1jfsJxq5ZI+2yXqCoiSIO4rHhmoBi9b2mAaYJACDbqt
mYs0b9hU72o4f0z1XCkGxhLXQljWRqi8ZqKx8qxhzdQSLMEvcY6jC1yd951lWMhx
EWnEfnRHBVHn9CMBx6I8sRTRiVp3FmxSGbX0T6ITzrX00kQWPMWZp/OSS/jcDsDo
yq35RZqU37cFoB0yoyyh6KcIctXx6tCIXhCa17M1OjklXe5V/XZN714wYOy4R5Py
4u2X3PU4URuDuA7//tYB5qqfmAkQ8qIGJAIeShI72F65Dxpx5U+RJfWq5A8qtRf8
pqAh8y9QVEpEEXlrd/tPCFJTxH+cDjDAkbZ/Ht4XZTu2M+ru/bAGvpCNqtX7U7Q+
x4sPEmv/8I8pmnSXF/etEuTJFntKeFzdGAgAXOZssdM0Fhn7CZEoLvv6HlUyxo72
+UqZ9jRF478K6o20vSpF9oomBQpi3hMLxjnAsNnlAnPPCFAXmz2UlwMVzF1gOFGl
LUMSyu6OPfBrfGzpTlt00Ebd1GEaM/BA18TDbZ+ZfrJZT6o/NsOCpKDvz6Yekk2D
EOdtOyioonp+BSCET2BasHh8TSKLNQl9r1XcJ1gXr+XZJxh1d+zxrWLcpTTnKpQO
LD5Lq5rjOaKEGpqjI5LPzdXALXsj+Va8HTyDrGFcoyHHRSbvlA+cYaVjNV5yHGQa
sgF3HE50yZANHya/TVWudVCSiIRmKxwvruPpuVZnZdP9NTQb/IJLxiugHpb9Xukr
yoPoWEcCtPZS1Y0Fr2Cmi8DFkOaTdLgMmNvMmYWjpn4aE5w4IYWFgYY/TxQtPayG
f88zhE+2JP+e/RahjWXp9Gs6c8dRf8xrWyyvEHK61TeC314BfEZ8BmmyEYLCkU6u
BOCQW/FPDmP1vM+byfnSmCGb1O7kieEhzpv9XE4dV+tVCrOQ98e941WTFZcOIPeH
mZEOStTBrGWQYzK78mlOEMTn95NWC8MCclsNc2fec9ujVyx2Cbygib0cu/5Bf0+X
wZpnDDcMLfsaQIweiDhruyRoAxQyQfZyDjFvE7mdtowqqi2mLTJWB0uTDehpvMkT
36TX7b+CLWZ0TSfAqHl1WjfLSy2Maw/En5durX9sTYDFbNDCF8kZR/wmNEEwhT7X
4LyogCHqg4XzJ77kureRghqUGvn9urRpcI6Om0FmCNTyOvIlAmlvWl/egxfnkrK3
LpZm3Q4PEWJ6BFNk1Am+iX8KujiFYYTjJvso0Zevm5UAT1Pux+rEe3FlTvRr4f5I
cTfG75/N3f8QAuYIO1ejSj+sMgP6SZe3PIYMYYnvro8iX7naXh9ke+G0vq7tcpYg
O7Ody/XDjJXTsZIbo035Hu9yXKiSgyiMr3buQIGK6qOE7pD67v3/VRy/5Nec75Nn
r6htY+yQActbFUJbwqmv3S877mBK4GvBl0e4N8728tiq/EbmCdtDeY3mVnt7hRYZ
L9iwKDR3OyoXgQchqUU958J+1ACiduBeHwhBMHnjYlS5hJhaNcWX+eS/j8JYTeNc
sKXSjYoxxjcMF+EgcFFv/aAjykUlWSUACjvg5xX6bLCNtvSxwJHgc2gHAkf9OqBy
qAYZj9xovpoiDVmbnWqOqiZKWZz7Ws2xkYMqoBLLviwkhSLLu32geUlJj3yg9psb
6cpijsSIUEARBcr/H89M9UyxB8G+VT18RgMIy+5u5BX0GYEqaHSspuIgZvaLsvB7
xNpocIoO84b4QrZuPC93usYeU3NrJwuSuwMqMAlMKWln0tbWeghLi3Takq7kJsWF
GNLadoV03OhmupSLbmk+Pa/7RT2Gd3k0OZYsfXH34kjFRjRKxShW+vy9uYKld5ft
BG8EfSnngvRlr6TFCn0IsQipaTz2LlPi0o8PHZpILgvTz1WudPNC/PFoeRKKTSTA
RiSjmGMbO3BPAgztXgtCYrJKIZfXp9RYNwd6AEaTLyq3I8HowZ3XnfMnAb6mnNci
+mUQYJiz+Fc0bS1ImN145hfxXUCiNP63eyu/lxHKX4wyUZ1ibkVOnDLkl9Zmco2t
cBUdIWWp7sMqpzYz+Z4uXnTVDyOFrpWZGccTjRjj5A3KAAqnthVNB6qqIg+cQMIo
NNlbvmGq3yqXpZ4a9deSsbRpCuPbfLqPmNUgcKCJtb02nwNtv+OrvBY1Zc31MxvU
JOLSp9KoioIPFsDgSlnf88CJlF5lyndVUt2tiwAqtOGmiLu3xvasAOS02+MBeJOs
2tAOji3tS/BfJf95dOGPt8Expj0pJWTdeVy+nJNb87l6xsWi/KDCUyNUe6QJfzGv
UoM/ef7Avc1k4YO9JdHdJGQWLSv5FeNw9jS8GyNzb86Wdz9vaCWojJAAv2odXU4k
lNnWvapM2dUfy8QDPnigfBmmto8C3TQdobOx5fqZZGyN4mnhZ7KbCv+ASheSKqYH
Htzmi1Axn361lsNfqFDSChKYBBdVv5miDDHo5pgoYTPfrPWy+vYwJBMcA/5KRdy8
u7YBWkpKz2BGqVZhk9Y0RWC83Ui63l25bcAKR594oTYKyuf6cNWHrjHDsCkTBjZC
9ENqmorwByhTodiM1dU0NA4jO/ZPZcxfWfRA4Tq7DJVPSq1TtWaPviulIVpv6cA/
YbOIL2muzZ7exOFigyfviGeJc5Sbb39TOZBQM9EDjdlwHXa2ltGBnJQbE7OH4HNu
LZAmE1rZYydH8I5srTbnkazmK7N0tqb/oCa2r5yE8328Zs+DGFKuPZIOa3J3+G55
hjyF2bUABqnN+gG823v4iGNR0lLXivtG4kpjDyrar0oLzowK3LJYgke9c3InPrFf
wNNtxr4g1x6Ji6grhzs4GtwGp2U+Obhj50ACOgXhUDVtswU1ZzoFoJYywhzJmRSf
RzJo8ip2qgEJdSkxFcyhDmaqJCmhFWCPVsTGsKiQhCPG50vz3eN79zsR9i+OhCmw
3kggM+IOHDJs4zt2T+tXXgYaMfD8oS54VpxFo2U3wxC3mW5WaOOPCVig62NVufcO
OLlUTuUjV2RLmdSZmVmZFiJP6yMfhuvsQ3S/6GYdujwqnsD6O7MmPnf2zjt/Emas
bXmG0zu3Mfe3E2nzW52WErbPC7Mbl6VgqFhdWZMyHorqv7TMsmDAI81jZPL80ObW
iyCqwu3mxUjXubYPSEchabsCzbRM0999N2jBQLDPMoS58mwEdwsbS1Il+6Ypo5/8
2O57vXHuz8o7qtMYBrgnE+1iPvtHML2ydu5Hqo9sVLcbPbifFPVJBp/LlZVy0OmI
73kFGcrf5prmri+mYllBCmfIUcDmPTt5fgRF6SQMCv+9+MF/tf7YimUREPjfpRWz
LOIWjUlz30d+CpW9moXNRtruoeLY9Bg6L0dqwGB6I2M9hGZhxvvhVNV7xvUNvsIa
c8GmBl1ofV29hhvb9zP1rNRT54ChlT9TFW2mJqguYKZ6fJORR/McUBv+2h6U9SOq
jKVdK/am+W3wvCpOJwFJ5qh8qxtiD9KurIbtPlN4xj4y1+COkjI6yTVpG3HuqaEM
iyfYpMzcvxp8oN+2em66B12LFByqRfQvGxkwoDs2T+D0L22X73WSQAtVX3khjrO0
6v1uQ2E4pK5YTqA0+5Q0rzPnFxCOAC2zvDU9eq6ZhsmInJx0T26zFq15b4JMq6im
YUsaUglpiBqolibTyfzolPSJrTmXROIyteJbkE78k3yGdzF2NZqKIWWf4KSKbpRk
8vJi7RzxO98I8kJSGmlqZbcCxUhIRhSH+FpyH5w7tHeRN7e6peJOTVXCOZQghf6S
LhitGiJOdZ6bUFHml9aM1w8it4tI+Q38jW4QsiIdEr/kCrNdtr3uRnoIGsTRTxI7
UG1fXzhZeXQ+88xcNEdzxBCOKtze3qQpeVPCnN85h6WLTU6KqZLgGe4WYr9m2Paz
NUAc19W7F046xr+e1DqAkU/Zj/Y/Pq+WDxNdu07upEHvxYVMxTCiDoo8hYybLwoP
mxS2/iVsNxTQfLuawtHstOyws779sfUSNGYjW4En4LcN5w6V0NwO+NBMsutXuaUI
XSHYEJlKjBvGijSEPCI8eYcsoYhJwW5Xy6MbSvkcxk+91s2I5gF38MVKTkE0ff/v
qMuIe2ceSJ38jKvfwxFE4IbUrycPdzPNMgBqkTQbUquuyCyFxOUgEUBjVdQAjBqf
ksjO3AlD1lK4yuUVpSGQCaf2gg9gdXn1XXXWu1lYDUVXfecgRQixAbPsgs2vCQsl
KvnhZ2TKYe1DfT+6mp3omZF0JBu6ta7+4QhPcTAbZThwXQhJkWkB0pG3j0RShbP7
Rb8binkEhgz8ZJ1FNN2PVCTefMJbHPZptn0kqfoe3Jp1DT+zi+BJPPB2AFlNKZ+l
lesUbIP9oofSU2dQqQ1z2xiZobF03AJJ4NjNG4tv6ENvClQd7BNlQES0nBNK85x4
bUzh+F6LeZ7XmA5rggowPtrIT1m+bQQ6QPflIu/56bDC/AlZwa+37kpp8E2awPQY
0ZVNuwGqN52tFHiSpge83WWCKUbbNiLvz2+gI7+Fbccpjgr3UyynGkhR3uxQ8jay
2gxCB/kM+usKpSo3zfhO2VN+L3EjmutUSStKK96R1KMxBULnyx+U1i9sseNqno39
139p+w96av/HJi2YzU1Yxd2xEEoaD92p1VpohbLKIprmMDYcqBgp57MAuwA+uP//
gl48PT6EqSejuhKCqzcu/hJtV9mMQPB6Pv3Az4+bSVbQJw+wJUqQIytYZsp0lKsq
r0b7XedoDNB0m/pRMu9USIXbyP69KpZ3/7NFoEJ0qymH3UKS8553Yuosb8AKf5Ie
OhrgQe4ViRE/4W+yVWUNgdOY33kHdZ6BtC8kR1Bb/iQdDySdgrkhlTEfQKLtqF0o
HOmLSdljGL/ADlL192FWFYrzUV+RyxmNDCgRR561R48c6mkcuPRIWSM/A7Wedl6b
sE14ma0tc/UQ9p17FNk+1kj3xzjYUMnHGl01+pb0OYxAmfcFFenq+OGozTYMqC2h
sEvUYuIThmCquOYgGJUEcx2ew4vniN6uXhe9IfU0E2cj8IUHsor5zFFyfl6B8k1r
pOcvP0uS/ueLwSIMMFJ97Y41/dFE6RcqiwxUa/dGW+h2Z48nUKmajStW4QExePFc
vfowA3B48aOzZOzid0xdN4aeoA9aTRB1EBFhevdOy1mVAXDYfLqbIddUywr+ox1U
0tazOsIb8vF/KEFtMQbp8JOoHEWusCeXsOaB4cWwq8FJfwYbGGS6xX29P6CRdK6e
lhB5Q0rnJjK4oauOvhHcVQ7nu/fao1r5K7OX+DG1R2VjKxdxC9Y3/dmIeUQn+BBp
McN9+eg93lXHL5VBxDB4HB3fj7VTrLU3n2CXeC7epryI4YKZPkQ4ZDYpi7+Zq8+P
HO+0MbOU9KC3JzzzwPL3LJp5PTfyx3C+ZwYPeyVKm7+7dSQxPtwbYs3jvR2qtjRs
h2xB82TkdSJO4kssi9uwney8AJ8P/ptbX8rkHKp2FQjHVF7Xv/Un2tL+aHRigksN
kRzaR0IC1wouW5dYrJ4pRhV4TrUk5K9N50yo6wKEY7nFHBoWl+qTTr9+ncqXB1i3
58bwuGGb86UsDERPz1UxtunVVHCOTHh3HR0gJVzuol7UKTDwbb8aj94/ytL4oYWt
DjS7JnH2e1JEsU4DcCVtpWNSoam/m8IdXDNtfKnTU+5BswIeJ6byiTJPaMHtSqvB
Mw+TIb9vQg/bKaC0zqDVCToeRGkaix52bOYSRNz+Y88cPQ54VrbM2xPAsLC68KWD
2IyAIcuKEDWcm5VeuLXOzEpbOW7IUeYNDXO9nZvUKn4JRWvbcb+F5ng1xp56jzut
fA+yplqj6dhsVGasvLkEtS3S9Z8QGTvejnydlaiwKlC3mr1vDfPzXfqJ/wFVckfZ
8/uNErJrqXLvGHji0qwKRUPXmOoOdcL3novHxyzCWCGBeLxIYlMeT6v2B4Q5H5qf
6p8GWpioxsQ6rfhelbL8C5ZmhXYt167O+nElmG6lOgxAc8PwMYO+ZetPo3m5wYAj
yNumR65rNZosKz4Vhb6d3RyP+qqV/g9zrZVEMWA6h21st+mwvuWD/gMZlWPSMmbh
+GLJoEidEGfiH65XgmdhSlIfVYg8E/CEIl2dZgcG43nILyEwTnKod/+cXAZ7a2xL
5EN9/aamZN3IBJqgJR5eWHtSJR3OSsE5/xWS5uZb8H3hN0dxvA8paYbBBabq5zRx
d2gWpb97st+LFhB8DdGxzQiJ6A+R1++S/RmYSPLI/V0VPcdEhrAoiZsPfezTVd9I
qCmwP/gJvXzwa4vSHkQSjvoXKwsDDqy84RVRDApz+LPN1GiRzQetjqjiIePJZxOk
SqPR9d9n/mDmc8VFhnqaFHnDzHmWP+YReKkSL5OzdrSHR6Got0dvFp2d+zP4svf/
aJgzWQV2oxM3Dijb3oDYuBT7d0Q6341ikWeOmZv+xMOhXud9tFIr1mFO9vUYSp37
8yUjhVZ+Celg+SG+/sXnCKZXswuaGrG2TZC79e93lVTSUx2diqLQUSWRw1Zj46Mt
VwfRmZxtovn+wkm/IoVcLdIsqK9avx/EH71Lhv/VBtS6/cEQW3ZiuYqSIvN9s8B+
ctNq/tcX0/wSJ6N524NNFGSDSPlPezUKKAgJELCOqgEsKz14+llnurB+rc8QAmUv
UTtUJBykM5IbpE1oS3+10xu6quZJkG5sE3wCS1O9GZgPW9ROVzMK5Yk1QlqBmEfE
H+WGkectnOa52mXeCUL9/vwP7I38myFUoMH8pzDeOImahifg+GIkBQn+W/mPiaMl
YG0v6iswvirz8NoC5ByKf4Wl6rLGJd25HevqGEz9VRmOjYqmXPRCGlsGvVOMA4K1
ieDvvNjTL5hYJRVNn++7gmyM+dCN/ZKuQsIXH4CxkKx1iZodWHvYcXjp/51mAuze
aEssIR6961IoTOsWrIOS4ZGUZAa/0wAvhfZCqy5pDi7A9gquTUgHSep2QnDiAq76
L02gnnRT0OCrIaz3ZL0QCGkCVN9GpEkZSRYlzcczLfYUXXcatZjiYwNVwWiIfaek
tHWkKkvbbu7qW/2f5Dwjh/2eumYPC/9OFD1GfEaDPMVXAdDXFJPlkZEk6LmLeShb
dA0wRQe3BCkiZLHKhqY1JdM+WfYjp8sP09FRqIwUzSzXMvi54lzAsKjMxCJv+lkd
ppkCbWvyPfKuhKhPVJpea9r1f9Q1V1DttVs3DQnx4I2NU9FNLPon6D3hQUtZEjeK
GDHEofHYqiK2X1PdCGpYYcjlhPS6V3leBvoVXWwULZDb9yqK9R/rrFMII+Ll0kIK
DpvqhvXC5mmYzrG16hFfy0y5pILYN3I5kmrdDsk9iOtyYkbg8UR0mk8MY2VnaWXv
OLgLFI+FX8ErKHgAJZb31Qd8FJo7mxq9RPv0MiO/rbVPZq0kNCy9+d2bYUhhG2Dy
6LULMsHRiVTu/xZ6rgMVXb/g6lKH5t5MpVl/U/Po+jmy1fTdwjPp6RaOUhi5++HE
riKbw58Bd5hdCpkNfuAtjCp9GTPLrfZ3NCVia8K8EnUtwZMNTueIvEnINc6SgTy3
lM8PxSzbE9jAXixPl5FheVUrWjYBf3tTltIl9QumSQ+Xuj7UYGEBHNPCT7NY/HlP
XL7fbSsmIHtBpcJn9aWbz5nbps9FoIa1MPaeADhmYYDITzOrRZvsTe6KBnK5wp/e
4/axpQutUcyk5sZKlvuXX14wi+jkyaCHDZA08nT/F76jchojXkRGToASIL7wV8gN
M/pSc1M+OxKBqoYs62nvZPrtVhx/d2PuJG2zEFGcGSSheUcFrUifgXWfSadV/CpW
BinnuF8pB3vZgcybbAazpWEnPIBzz1fvloY2zZYnfHEAeJNm6/rTNNvd1cW+pPOO
IVnINsUdc1yG2PMVJMqS9zjHkjRPBAnh+rI3SliR2kMu+QvdXjbSYxUmBIgmHvGZ
yFFD2MhAXZZx+9xe6IoNWO/nYyZcR+ljK3zWD2zg8u9Ab4sZk1bmpsQ9dKWuwVGx
gaiCLTLHNEGEW7CtsqJ/20j/RwqpjNwpZkr6jRMofdSuWQy2fJYxFJ6RTpiQ9Tp2
rjfrLk01Xpf9+2YN56TgnxmM3aizte6d4XxuoJl9f/zkjzdWs7A8yZUckv8S5fOn
63kFTopcuCTx5XEv5RhykgPtcTdm39zoH8pukhOVN4AkB3y4ZL4jvpptNxWi5CbQ
YyeA+CX+sbcbRNuxEo1LZyNMU3scBVK6BoBFAH5jv/GyrfIHYcRj2y44AgJtbW9h
08orsCLawzucSVrJ3y7gsbg/WaSK8IOk7MjxtgnAFJPTCeJMHUOzwZJy1VcDLXhU
vpU05FXPVMXMJT2YlZIcR8RgtFqxWuLDr1l3pyQbTz0Dr9hJ13EfarxIPrFWWd8L
phnFNXAuWk/PpoZK5Oei0zEzZcTF4iWlES4Y84ZNtvU8SAoM6uuo9cP2l4A/Aiau
JgG2Gje3aHM37ANhvHFzsv/WCK02jppOoZ3J0Kxdl9gLyFKJ0uOmyUO+5dJe2qSX
wISkRhj6o2Pnw5dWEKIzCGeuDenDJGUxN1LvVOu4yOw3OgXaOZmOOSj0+fe7xtpG
tMQDfMmnQql2+nA8uj8u6qvF2yfh2v4AHMdPHdTOaflmJszvNrlwFhUmdk62JpNr
RWyVRh97jRe96RiWi3j0cmoEv+0Dg21JIzH8PFOEUNcOy7ALN4IzemXPHeUZpZFc
pwRyu0jOLX/G3zfqOUtwOYcJZ4sRX3Ikywv/bvlf4gkONJP6cKPjEqiWlylga7Ob
6cMXF47TSFzTj+qapwdJFs/TmlNE4onpzYdTI/yk5rRAXdfifnlCA+qyaA/XmxE8
Zn2Y8pMAAVza49NdfHXr7omUz+205MDESag6yjurK/1Vk76iELzMFxZFQhAneFtA
Y0fq5TEzbLavtUuI3CquVAJ1eJVCXVDrQMZii2GUQPjcTFiWJjKyvep/0U0NYTfV
ZAxu2cKhpPSHUlMw+FgDm8Is0deeh/XWWSQm1zh0pLLgs4NlJb4ylq9IKZJ1Eq2N
JGMlrRELGUUohfuXTJmxcVetWPBQRuTNCdPNm6xZetF3oJ60zB6ybHtqA+C+mKjs
F9XgAmBZx9mZHnAVEJXkKzZ/W+WdFzUfWOqq7SeSNjr/RxCOMYFS9j0krgBPcAtn
gMb/x+yFHla+jCarRnJWggCmyeoXCqj+cWYGf02QrSfC1O8cKVBN2T4JacKAo16p
6xw2bd1a99TexANQl5JN92PxV1cpsqpoCnpdD47qB9fjROxpZOdPwH2r/4wlgNoX
IuGL0woKcvpe2ElJRlBdYJsT5p88dttCfMahRSxW7pH1gf+NO5rMoWJtXr4O8OcQ
pa6V9TBUJ4a8YvYpR+BUlyJTTf/zJJhF4D78lTpRSqElGDwvgtIX89wlRmDLb3bl
yhwN90JfsPRncRyg3OfiG9pNHb4U79FZaZ0CGl6jvCQjqg6terSG3Wz2gcXYfQdt
+8jzyP6Kc9QglYG675Hz5JLon/jSxW7BG3ne/djuWj/gKT/kRY5hQ+K+OW8DXqVQ
PHGE4Hbpy5L/gBLFp5uO/NPpKOKGlu/dApoDdavIGk+qCZNd9A8fSKnLaiZg7r72
3DNFdZfe359AYYomE4m4WsCRaC6nyN5agH0e9XHyGYfmQMG8PKrpkCQREdE1K2FZ
A4YNFPHoCO6QitpmFjtgmwsUTX6bCpacV1ACizuerwEGZwpr70ETZyVJIqOXMCVd
JhBiPOUIzKW4eudRTi0hTJMds1LAJeNl8xrEKtK2n80eUclPJe3zJTy0Sjw6ev+R
CuMLufiUaENdD0nuwbfSI5VeJH+OYb2MP6NKORO1Ns427ww18NM6fduHzWndeSoY
K6QpgQ5L3tKCn9Qsjw9G83/UoJulqNh3oUYyLfaJATlwaiDi0AoQI+o9TST5TJPw
00H+QW8C/EPvkMe5r2AHtWnEQnWKcaceSbQd9w4RBV3Gy8Xk/55enogK2S2TLfWE
jiPhQriST2gNhtbtQ70cO/EDb4FHG/ObE6XRI2o/0lhBBbKXksXJZvVYDID8kzNU
tHf7OzzbrlEB8lHlbtag44/SMk+1llGqy9ob4tL1IZmpNNByZiVD3u4qWk002DZ5
f3l9oYKvKzBC1vIQkXf6onHL9hD4pwV6Juf+YPNMrn/kxE1EyDBpI8Hd5fGz75HA
zAFMxcTxePCemm9bRYoM1Mi62SN9YJhZ6bpEih7hwBKJEJnbj9LRLy885MvYKDvF
4N3mjPW6eCx/zn6XGtb3x0A1EWL8DF3FHfarrs3gCPVCETa+4xN1EYln4kja+OjJ
T1ud11rju0ImZvApewu8z1k4Zl0V8qrp6ebmDhNZjO543u1yHeC+T0aIerifWW9T
8tx9m0A7ARQ+fwF1cTVy7surs61CsD8SJHlZsJBsVJIknTdOLEgLgYNJLyTAcEM/
zKTMPRsvmZ2Qw6df6q7q0OgKV9gibIHgpOlsNm3EV03SWS4MWCr7RjBmeLP8o8ED
sF2xp1Ly7HkgKM+VI54zHE5bguAof1mXwCuQ9cEh7KElQfLMp5V88VhYsaoG7K+P
OpsfPlm2N4zeWv2eM+le+/YzldrTieaTNeTrCANRi1UPdL9wUVG+FGuHYPbJe7Kc
E3SoJvPb6ax0YXOm5eZghXhNRnFs+sJSjd2xsDHZgKhs2414hR1xJR2y2wygrI2/
D5HJEEi+ziMXv9vdaMzGnQCKiri9uXAYOOKLjmw05IwWLjVETLJbYDghzMdypYjM
sc1bmArcY9FV9fX6w5cFDT4MMhf/4+hQFatQQ/O9TgxbNsa04y4projD5+Qtdj4R
Yf7p9YrQPLqRQhIUeURqOaXIuBh9QiFr2QeOhdbdpqwzrnnDvz7cDG6UXjkcu7Ip
4HaIy2puBx1FiKzEmxHBhw4F+8KsD2HD93nzqxv4eef/wEP9ZJfgF1HtH7qR36Xz
FLGMgDlc7spVIxnhivJlWV8jkDKAp5jwzpKqBgw6vdYGvYOmZ/e/Br7kgWkuY6Eo
+IUawqj3SH5wZf6lScY60/5d0I7XG8q+EhA1z6AxlKS5fgvZJQSLL0GrubD/s+3L
bbm6BGu1Lv4vP4SdCYrSeQx7pjhFIh3L88v5re60de+fevSGUUFjnZlAJ5LqWe3X
031HFuCHe+6vuCNAURkEGI7JzvCMJiueNsRxe1GKGWrYwZbhksciHSxyrzWVn/Rs
ATRmhkCBTsd2jcuAivfreHGajsO4jGfhqGxORHZH8lhGLqEAfmcwcU8Siuc1bFN3
dzCL+YrkA8kLDEYe5RyYuecXL+P4GVanSA4/up2JDkcWIZw6c6QdQYZP7LQbauEs
/+Z4jzGoMmmJPU2Pym1T8RdaaZl8eiEhk5s+/uPMtjsVLjmm0+VcT/q53SAIzqMt
bIwmdbRo3+SW3+CIwCOovjoFyB5QT3Cwsnf4ok7TzZ1Hpwmgwj9HjI50fG7WdKV7
sy+41KCBA17h5Wf6KFCMlhvNvr2ZTXf3T0KZf7Oqk09lmLOD5yTlamXlfXWcgX6P
LQWawafGcwHAt/3wuKhfwTzj/t5r1c+KuuiKa1/TLrKr6Rgz6aLF6Prso9pM6FQC
1Me+5FI4VxscBrZfVpXY+P6ehgfCEduRDjEeY8Q0vWAnXLFbAHuzte1KKJjhPpRg
u5XSjpnRIveZnjByyGc72WUEt7zes///i3B2yE7cuCJ2K+R+qzozZZ0DmiVIPhCP
cIXSQMf7T8rkS6CxEgIQueOEr5jRjuUEYxokGSOeWbL1tMLcnDD1/a7947c6hnpd
nPndxWTatJyPJbP4jK/ZYZhLrjaCaNVumD12l8Gfu3GyQZ5OhO+gfE09uWedkO45
juu8HgsoMK6FS8xdaLzPh4O0gtiaaNQWe2EMqkj3upvcvdoGAz80ASEnHozZfXtd
+pYsx+SjIv7JX9nlSieZ/KL4WAwwAgWuRHs98qwnOmr04y15FPys1JZxj0q9EAz3
I+RRN/NxkOlKbdJBQpVj5bynhHgc4Mtr2j/0YbQUHVxUCpOAeLp/5xJQApA57UKZ
za6tHJWyhV3DrI7lcrWNCs5yqiXdO6/rxHqyCtVi1fFcaPyU7Rph0yGEvvI6e4j9
nD2IeCgiWU0aepzUCi+Y+mCA9AQ2HGjZMs/FCu950uGtR8XwjVUXEe7XCURjccKv
L8g2uwv0tFGGvD092csznFwGAK5QsxigWr648GO6pQo+lFhkhNBLiAhz1AC3rk2V
oyoiQHjPD008pUbg9JqnnZBpaTwucH9p0fkXJTI1Cc8YHXw8C9NJP4ChvAscAsMT
kyHtrH6gPUxDJnG1k7T8cb3/cl6HThogbSrX84tWcJG3/vixjikZLVbP40FRoyna
yrrKX2QbEhrEmau/4/RaKpsFnO/RyZ13A6DHpd2+nkJ9H7Y8PkIE0zgbW6wCwn7f
11l3nlrUsnSjvMwFvFa+VrzxuylgvlopAd2wZ1wOmwT5G/MB+M/E6FiXELO5SGH6
mleTXQHUKr+JchT5xBGRhUtYV5ozo8kV83YKt/K2NNsTWGtWDxLQq4tho9ZZlcpF
Sw75Dj5yANJxiPq0jGfefnLuXNXA1eHcqhhVky10rwMq7/+YNI6Y5HoQOaQpKSMR
9oKG61Ffx+I0kT7P3SA1GHdIwz31/U9BbBvkdFMRazjAHDcHzUoQ/SsxXvzgLaTD
8jUD50qo0pKZmMPVJV36CSbAfeNVZ2awyOeOMgy34uRX3W8ZXx+ij04i1zEzdD08
cNg942K1NNonkKrce40i72D4QRCm87fEGsGCqQ82Uli/EMLep4+Ix5FhPtV4QTzX
lij94qY789AjP9+C3Qwxjo/cpp0Xnss6zHBFqFbvI1yvvd1LYImFY8stsMN9pQmm
l00uBTmqq8UqVWvfCj3bDLQnVvjGUf5s0IkdijuMsj8INxoXB9hA5m/gJglfTdwy
5rh4t3rpVQRgxgrhQ4ucaIVADdhEUQmzsITW+KYDbyk9l2ymFKK+U7uucFYa//OH
gNGEl3x3nM7L2SxmGcuIpFj/Q8cIMFrKUbBaGJxRpMpEFlWEz5sKcdRa5TPXi/z/
EaEe8TdLqtrR2XhjqaIaQhhoxiv5m0w8zjApPbzBQ6ZHgXbMRIc0tgySO+CTMK5K
nFCWo7J1lKat2o59evU9vxjuYRULpmHfKnSwp61Zk5BUkV4sFsM+rSvXAvkIBXXH
dxg+aMGX6DICPC37nYThnLAtKUp98y9I77gwZ+X7S4riXjrZJSBfDFuqYVttQt7I
mridVzt9QidJ6p+1pD/nLVB9M96UxeVHZjD0Qlh2Zehf++uEF1lCpcQ03rtuTDvm
OZbgCGP37GO9hb9PYVfAl/+dlkLlSvhNM4MqCt8GSXjdChAxLErt+lzBNs1e4EbG
GYUFn4EkxwLdCYjY3CqxunjdycX64s204qjW97xpdo2MjkcO9TIEwe3wPUq7yCFb
lEq2RSiWfVLA5rJXnJGB4Br8gBuyylrEDFgNVgygh4U1xepz5TTQip4ojp8bYu5f
PJFlGSrlmDzXAPzBd5Jc8PUpjhriLVdFnGRirukplpp71Yq7oaOOHOj8OgFiboOI
7jIkj8ttpmbr+4Wl8aUQ18IxtQLGaVyzXQjf/kE4UijT96UbEbrbh+v8Gd3bHL3f
ek+y65NPMLWUSuP+nl7GCKspfP+BUf9XDb/0GG3Yz3zuX5RPDgP19Rs3AHsdVKB2
7M3nHxQ2BnTVQFsusArEJamOndpVfx9zv9586vPxPsSPRARb4h++nDYe0R04eUqC
JXYUKu/LNc0Uk2MvwUeSwfspFbwF4BWPk2CFIg5AKppYl4a956DWv2Uw7bx2uJss
JqNET+Wem6wkMcVSNTEb6EKFzhXlQw/rPo1fIrFbJNhjxMcAY5xWIj7SZuWchzcI
aYwVh56e1u0QUoMMULdqGEAb6FzvmuuhqnTPOcC6ss1t9CX+Ps8WuHJOdUpP3Hmn
n6dFbtdHr4mSoJg/pvaM81GzITW4nw+IycOIjN22+rVzaFTC8RetXtuOOiAWVEni
XOTVs9SEI4gXIkoXeMxjV//A+u8P+sNdfkOf12LuM1hYiM2VvZF4Btrd2qE94gii
Yw7kRHiGkkUGiGih0xTEqi0EmkMxaRTSCUGRxUoZjLahKaqan4E2M0eL/RPseXrZ
gbio6RVs5lHLKe1vFlNao6r7IbGtzKdJfdZRnJf3lDyLt1Mp0b9YYMoY1fvki/wV
mhb0CqRs3OidWSe5DRv1KCV7LBJehhwR9aSHvOa3wpgcehh0nzFwbjl3ImUHzmO7
4V9yFzpeDrcOibezZ3TFM7Q8y8yragW5UVpobnqr9dhvLAgO2859w4Fz4wWsI6g5
jrYnuwJeppaRJAF0T1qXx3ZIJXoMFF2PmWDvXoVyT02NBfxXEVmEu8+KvPBR913h
fA08WVKKterYghfaTA+l5Im3cjgdDhLNhTmLSu8sOFxvg/1L2tW+WLI6Xek6SxWG
3pjUczv8rsyWHL2AO25243u3BUke0mNb0JDuE56vdLl36vP5XQPHHCa6edvEOy5/
6X15Uh3KFpxeUVeHQwE3FVCr7k24/rZamRn04pHs/Chcz4v917HHPPuDLjFmYDKZ
f6bbN1ouMhUH30yXyJr0VFU0Ic8DShfKctCGhUya7TFBb97ge+sczKprxxK8HTVE
yQrehx3VS6o2lBV1AavURJmboPyXgoGdEqc+eB/qC8Xgfgb7ZLbzZM4vR1v/O3M/
vum4bbG/8bphgqQhY+u/83GJF4lrEynD1bZDlucKRMjAYB404aWTzOIamnrpewks
xPkE55Iv76V3Jq8Q+2rxs0enZGFF2eGK90Pj/DLwG+W5LpdIBoL4nzied5PxAUp6
qMYhUHbycUlFVKiZr8XNlDzTDHsaMZn3zZ9qdL8pFf1uHHNUN/lEh+W1MnLxNAPC
ZujP2QbKjZ3VX46AGPt7T7iq7Kv6F1rZsMNroVlaF7U0BGjw2r1z7ZMEQpXJ/9L7
FU2GDtgZyzI/I//lxedN8JBRfJCzE9ijigYGP8b4wi6ga5X/yBdfu5MZNylkwgEK
mB/eml5HR95BBo5U7lT7sZxXAV8m7G6hLwb19fOiQ+0/8IWWdhqzgYxQ7umsbb30
MkiML2oh9a5fYVoQOrJpnl895XJTvpg0cHKRIyROjr6DOGOcEYNdLHP7b4BC+Rle
KlsVgyLJPRqhG/Fk9WZhC8fZ/sCpjxlu3tUbo2pbgez175s5YCn/WAeARDRZOJTc
kggg4IMg9eVgNkOPvDyOjECohVHQFlJWZ6AUjlYUqZ8LJK1Uxj1dQlkqyOax3M0E
9fHkMvQTdvaMzOWrs+xyq4Gire5wsPa3zjuZkeE4uhxjCMoYzrCyz7hOlNjRy7/d
15uX9Rlcrga0O4/8Xlv8RiW7FbxJAXPiEPkS5OAQmwopV2pZvVGU832dRYzNcQh5
b/ygnb0coMUVX8gLV0uIqS8q7rx1dliN2ylFkaQkrJSS+cHckfeWLozMWVs+lGzr
tqueUn3AnmLpQp5vMI6DPUfdyRaCWKonR/B0ADk5HfZYFPBb7+l92gUMTEOU3yck
AOtTSZLnZZq+OB2Mjj9tyNOrDp41+zv+ldKGYGilMXADWDD8VSp6VwTf68djJjV7
dZRxfzltaZT4c4MtNUHlttntPLuhTZlzuExsQ+Vo1zzD4ZS97VBK8iiIqYMWlV0h
ndYkVnwz+A423xqbWC8hWNeKFGLFxjdPm19A3bcytHey0BXlmbTar5bYKM2Ipe1k
6RESRixzs9Bms7Qb1boiXylXOom9qufBe7Gv8/AeP1n9cWx5Q0J23GF7h9aH0Od7
5JJuZzQLzLo2hHEZlGJZIRd/Jrnv+4SDVDIypZRM6c4fFKOcasZcNwKo/SF9YwAr
oE9Eyv8p+7JaoNAaKC6v+AofcH9ofmSYvWzsLCKJFnej+AJyYfUuqU2VJ5X+U8TX
vKGuUnCO2mm/0BI+jxwJhtDd1vFK1q5VvGn1Sm74pLAEj7HBPsic3XhkIBjymdBI
BDWAY5Q0FqsyVE5TdGm5OQPp6ZQzHh8OYdf/2vlPBur1U/iWqdD+YiaRcXB+uzXu
AEO3OCvp8CP/bWCcuTtbFhPuV1y9ygXdVwnmXMozmse2Dzi6k6eB45BZDqnXRLa+
rMub747/ezga5uL+Sx00DjVGSiBhgMbrcG7+PmsGEZ0gfaUG0XdVwJBH5pF269NN
i5UrXGBOs0CAGLHNVTbTUlFQx3D1oBPFmxsPabnyAYPeJta4G6FFjarRaEAfED9E
suSrXD7PBUXGg7qn95+ogw7jwYVSZj3HVNl71FbcPdjWdkX6YT0rdlq/7SnOR5c2
m/99WC5t9mbQXcZpJPnpdtzCyiqR9Bh4oncoBcD+a6XiuVAZcQDddKGKHYYo91wP
Npohf+SwiFNRkAXxGb7eV94QJ4tVsxzCCfJmf+v5jCfWKDliy/aICh+jzhh9llcq
CzD5rZCc2EM6nl1iEZn16EbohbeGJliWEMJkY2oABPs5+gGQ+X8my83XZji0kS+Z
PdIa6kP/YRXM8elIYeyhdUnJFxIkfQ34aBNBDF+FSTwezzmLQoByGw6pLjUGuUgi
norIA+bUi4HP0aW88G7YHMTtg/6cJvOk8VR4dIm6pvOksJX76/nqT860UsFdEbd8
kcVR5DBhuJnZH7Ll55kMvO7dTjo8z4PD9bT5VHkzBDmEFu1JRiYUqUDuW6UFen12
aQecyWwetjRCvY5Levt9Mb7D5FGk8Pj2MaJHCniY+6fDMFAiTM12MA1xBRiOyjCA
Y+wSaZH+q58Af3yj3YPV5C6Gp+ITrYk7fT9UuoBWen160B45QolIXhoPhqTQjqEt
M8CVscWDVX8n/vCjMCBytO9V7bJpC+tWu+mnPmmz62ytp0I6vC+yENHKzXBY4oaa
IhK0wPvkrDMGaNTGhuHRtg+H0m0kHA4WOfUmTdRX7CTtTXWTr64IuvQpeWzppNUy
cSlhnZ2dImO8Zu/HCSZpOTkKE0ulXcnZhLZ67WVB0ZXwB1jDIKyO+xFMPe+f2PpQ
DqNr8hyd0GdoKIpePSWnxwBtLy8O2Z+9wuKBgPz5MEgRJvrwxoJOxciE3yjPXtut
kZUCG7HsRDJwdxd1VdIbA8PrS39EHDFijWHI/N/u+I+aACAiYbL0sVIkMAs+Rbu+
WUi3xGCwYINCBtyGulJaIsVZhay8X3/IhIoYMEd0mSOiamgGYRYrIcx/ijL5CHR5
reJAMaWFUmpa6NbEAK/2b0cBkGkQFBt1McQqK3UwSk9QvCGlLAaWr9fR9UcUSBgZ
enQ4iTAZsY9DFnlE/NJVRP7QJMR04uV2KSiZ4lurkRXc1Is9/bs2zPJqckgBxYh7
SysP1Cts5kA7F/meSuZdK8JxgHd/w+uzSn+Gcpf8oUXhOcAOWLFzzL1ah4CiRvHI
7rc37s0pvEPcYJV/jKe5d8w7OkvLWZpjlRJ03MREvE4KwhI8ulVvUWrECu4caUyI
DVUO8mqib7jqSvmptvoC1MnZ12peapFpvIZuROPvwyx/a7K9VGTTTQkVWwUnzvjM
YLUO3iie2md9pR+xLmBOcEPrC5z1XYBs4+/DifIppOjxSh+RCjU+/Dto/Ij9E4Ry
3mSlnFImZd+ikDtAR8KFhISkyXEKRELkKmVWmivM40uH36U05GEUOYqAm7EbDb2D
bt3o39kD3fvh5JHLCx5g6RjHaxCaiHxHGKvJvozO503HqDm6F3aGa3jAo0IX26s6
twiwpVdy1oyApT5A/YNCARpNHE/j+Rjqb9Hz5ZdlSU9B74hmINu7iA7H+oS4H478
B6cMcYBdl82KBmU0Hi/vQkS1UvWkJO/a4MrbkUvBuxzMPfEDevMBtheTOA5Dwz62
HahiQREPvkltPG6lgdh+wVyeD9sq5nvNWivR90w8/29Ni2DWtupMluzIpEJgjFgd
DkECyH+BibLO/DKQ3CFemvbYWYWhYDNa0in/HmU+Sgr5IaNH8cZdlAHMdaGa6px7
n1NAptgaYVXHuSgenTHmejUJY2+9C9IDteDmYg32KtZofNQmSKmmqleCJUtokOtm
OKBVt02ZjW4/oaWSD0V6R96oFBDEy+I4iBTM1x82tYhz+qQiAKGnubHSj8kECYyv
fQlmvVlNl/WZ1X244IEzrw+zCngH2jY0tyP3bBPotOcBRssGluXuRxIsr9yxVBxK
Fi/S84yJqM+WdEx8i8iFIczJXktLyKnsaawmwbR136DVVoX0dyUXGMx02WO/6Yzs
LvczEsTdUpjDHTf4EV36SzPgyaghIx82Gh9HKDJjQsqZjvPEZp5Tw6XFNkJH0vFL
b2qAuD8dGdLfrZm3porbzX22T/ukysQEOI72to20aFXeY1Wc/xE9pgn12Ss12m6j
az+Fen9kEMRAkdNP/d6rcIr3R3eeRdU6MqmE6ZnzDa8V8YE6QtFoiTykMDgRNyW4
ssbqDLL1/eNgHfMF6zOhzioJaL2qSbJbXqISBaWaof/BI3pBL15plxvla6YWQ2wj
s8UZmkkR1rpfAsA1fC+SJihHKtHXWjHPt66R18quPUN4Vt0Df2cb3199Swwu+XjP
UoJbKw2yr1k3w44UHg2al5mR+Y+cRcFt9F/6L78PDzGItzmn/JjmHmObxkOHzjZu
CQ9nEQwEZ0LHrWO2ezBLvGPJ6Hpy+vqEy9PAB9C6tIisIutSzSGkr95zDGOEuYJQ
0QIOlYTjh01+8M7TtBmkX+jFmRG6R9Eq5txmPxLbon1JPqP5rKlXztegsLDNGDNY
M8H/wqOBN87EQzUSCY9K4RxwMVYNT4auSVutQfBogrN0VtxOtALAHsv7LHfdcRLH
v2XQt6EIKhYjJmAWYKNjKztDxCq7CBsfn0Qw8aURr8FEtpNK94t/LDPaJx7t1yyh
wykyQg7DFE6Oa831tj/nVFzo+wtnRkeCakt6Z7+RbRnBF49Ua1mBVIUa0fDYspCR
EjNo2HKOo9jacdM9BYv4PPLb6ZAWiC2T4xQcoyhULS6FsNRqJ+K09utwYpltSz1x
Ub6ypmSAG41i4pBfIW2bVAKo3QQonn3yoYpAWh9Tg5pZkNldsr9VnuryUfAY3i3d
0xPdY+xKDC7qB5dw7JwL7+o0Obr/+vINRuh1/eWQBQ7qNdvZQyGUIF5SAqqAVf9G
w43YluYSuXgpdJXjBdoR65OlMHv/cTVXJJGDnkBHB/ib40dfxaWjxzvNM9zzNw/t
F6mfp8/U8VKVJOQECaxm3y/yyBJHaiMrh6XQdC3DZGWhs+/WcWT7icMhb/nxUMd9
vzfKCcvIOPbivtkYP4Nsu3z8uf7xiDxel4sotlSNPO0mlZxFVrj4P9LLoCMgb4MR
1mHPVZE/qSdtwZ7LfKpT5JBn5vfP5RzyiiQzyHbqdeMpfBZYTghmD4rcHcPbMr41
+YwzQxeXQZCP0xzURSccggG2qG4KLEvl+lEEmq0TqmR7FSao1MZDqt8wRW6dgod6
eXOspHTJJw1+aQBU9PKRRv0seQq+HqLY+7kE08WvdJphtwSvTSGKdbvkQ9asSmkq
MuU7K+qR9vdpqrT/tBHF2FKc0I90l75G2hPsjKu72QOV9FL/fjHBPcz7dAhoiy0t
7P0TDRT3r1t0Hc36DLYYmdRCiRLiTl43Y4iR6R7j/aaWl7bhZm9/SPsTIY7my/9s
N/s1ZfgGkb/WadBbEqL75Kfgw3w/Y8k7zkv5rAjLMiR4uM8HelrA2cjUMNWCaAvb
CqAlHnI4v3U1kzN8xqUROtvjqYydptrRcSvnLKXRstSZZhIuqgpmvtsKklAiMj0A
bJYG/LNuQSC+UJvzyp/i9kCTBVoZzKLqMaaOhjhrX8ch+T6QlE8ljnEhykmLE8xd
deJlomcqdKZSJbTQhxc31ikoW7ZJyJJyiain+WuT3vbNpoU0kfbIdkrUtLVbOqhz
gUHkVpoeqoUiTD039upX6cw9NMrq55nsszhjwnYu3NGXupczYIkZoKdS/jA6pgtL
6aqYi97jAFWPOt98BptyrJ0DD3HnXD9VeOcX0K3G0X1gE/oYNWRSkO1EN8ELBezY
6aMHGT1QEs2csddy7uDEp3rTKupSjkGvb73GlOUWGa4JOdfU7H3GwhhE2XCAxgV3
hWdV8zh+eTX9VWvMkVzlgnI2pvn8nUKdPyx5yj9Y3IGZgvxadKUnr3W0y3nS+Z/M
JB6WFOu/7s1DFFG0SYwOo8RhhMbRB2M9uR/x+ZDjLnSoRZoeSPvNqK76mG0lP69b
RfrW/dR77MnpKBCvdl+UCRMbvTnUjsmYzyNwuYIMUASGabJNQnWtzvYKQs3hjhGg
jdKZ63Y9JXg0s7Dk2JgtuHSC1LU6aPPK7OHxra3yVaX5lUkyT5mT4QeqgoihPBTD
K9KC7rTj/f2mr6VtFqbt+rd6ZkZlzUdZx1Ebwww9Y8JnpW+oJu1jSpCzHhR16M9K
osLetz2MSTUY7oCoh0/JhyC0RnEUKtUwPW+aTNGm/ZpWgXtRgUI6vh5tTom4Smfq
1pdQZDnwotrWcR8dCZiA0i6IrSiuIYxejiyVGGY1U67Fbfm+nTwnGst7EbeQSG7H
ABqL4YjdPvkBEpAHnok8cvkfzAKjVv7ohBvDt5q6/KqMWjvT1ha5EqABfHJu4EvX
hRAbsW46hlLoHPo8IFUa56jwZzs+Xtcwf9ywfXZ77S26rtkr5Tqpu8FOIiZVLW81
yPGZFD+3VS/JJi24ktNv1eOnvdAt/IqMuAPcZRp3FBj8l2UoeZsfLMZQ3mLCR9P/
rf6lzWScIOKldA+r37j5GgAAdiXTXm6egFm24DqykGwBf3v5eHqYHBIeZR8l44gy
U9jhJYY4atrysrO2/l9ovkBi1auomCnlok3oGpfsQFZg7pSriDg5gSfB4d2xJMNH
fOZ46WI2QhoPBr2dxsH9ArfEBugUyhqNtj42gm/gcfEQXo8Rgh72u2PCHXGCkbV9
OyJPc3Z9GAUvxmYb1Tdw117OmpzLlnqCsr+KwZFd7ZK7Ws0iTRYCinJ3naQM0k/b
bRntfSmKdKFH1zHqrR0vgmDCzr0CEO09GXDcltholHpNLxQJ9aq12s+l3siWsCiO
ybjxSeCRVcrv8vQswQPAhwcQrlRpN+SRlgPyCZdqWJdZ4vO9rTUiJAZPBR+w3vUj
jdHDue1tA0u3G5Quf/HhfZPeLXfDtuHRN4hKA6dj4qGzxj8h1LVeFf+/9IgXZIyT
XcVeYdDfkyhk8fnTMEpFSFmS9kG3gHz4IBIOVRzILzZVmUkThmO/DidzDvJSa4qj
di9/OLrNgi1xXdSjexG5ebZT9tejQ6SGV40O0CLBNMIHgEZp9q2dn9DqCXY4w3/T
HuvQHaMoJ7iq0EMmkBeX+CLp61ti3FdbfojxQjoUvYRwZLbIe1gwEh9NF94bDPSv
eubPnq3phcQaetK7SGOLNwv4eVEiOlIuxoeLBUiCOfU+yIhQK73ogNFe+iHKiX/c
l1gy3KIWuxX3bdOxh0A3kLJqok5GoUic48ZlV1zKyL/44mzZXgi5URV5lLquG4mF
xK1J9H9kQdhGwcTrKOB9PICWZpS++/EKrZHsjAj36hLeP0aeDC76DFf/ZOpDOa5j
9pl+QhsSz73virLoyc2M1jtgHCsfkkbtM8g5licxnpdIplvsaoeYmyUALdUK3wtW
fdpVx7zZ0xXLJvN1jO8wRWtKJJyfDvK7grEPo5UOAq1KsJFavrp+aEwsAsI+1MCs
T3vW/+3Of71d7JenMKqgDcPn+duEHjMSreHbMB1Kqe1AouX1pKQbiYwQ3qA3+4+G
c8N5eeAjotRDiZfkJTXY0RlNyX8hi6np0fDkj2XhK0KnP0lE/GbfkBhXsAS2lzny
EJ5oZkT4DuuXKjSRiP0YLdmgdAsP7PAR+tAVsFijN3kRejzvG+gfEeDz568rPUnM
7FT+oqGwUbjV3xwUwWJKagJuLkQoOFUVruIdmVNOVRd5vZiR6c3hFM9M+54LbS02
AhqVJCic0RNyZhPolgLNd+4KijbG7hxwCEufNEUrFNmGUU6nsk40JYPqTuxDaUql
OjpZAHtXRFE/ZjtIRpkpFs3+CE2u2s26XPS33J4p3ih1+CHZ8OK5/zl4uL77HppL
NvrtDUgYO39Dbw4prcOOVYVbPBATXs8i4qK8D9Ve/klqobQUc8fxN4GbMZcbG+ZL
e47U532IQIZh/9Bo0IGA8mq3Y1+NR7Tnw3W4fIcPX3+7/uyLXRLSQzXspD0NaJxr
7dsjwKu+lZeFRQ947l6sPoI4YjzrR1UN3x9Imaej5/obTnkf63GVRaFwZXldQJX6
YBNR1WJfces1JUrIkITHsZfzxFvxKiXX3EQlNTCil1cTy1VJ9Tw4MjQpyl/NsRrU
9QrR4P2YDj3nbX5YgPZ4KctK3F3Qu5OUmrWwZdNvPfKC+PNC0QHsTZJLWEGp/ZVt
r0L5iJExnQhKHftRLGoPuw50Ii1GFH33vOAmyc/rOXcHLrCmZ5ycWhbdvrDBtHvm
VwA+6vCktmpULux17Vbe4VspAC8YWFYcd486QjmfP7XUEdOeUhXYDIghfxMqXd1H
LMlF0wM5zdI/ShMsTm1kVRFMcRAGuRCr2YhJKka9iBzp1jvgwYeduBXIDFCGIa1B
5P9HOw+2UugPaDAXQFRgaU6dh60WpBC9zurPs+aj5Y1kUqThgI8Lo3d7DusbcjcV
HZV5H+63LQ4ysTiCl9BSDe7GSWQlbVYbt/iVxsInN1EwEbkZOriJvCQSqxJ07Wyd
qNa97m01G8PSWNtrMBJzMTRJuTTEAOdZmVHFGfFW+uuDcJJLvUMl3XLeNJez+kzO
f6ZPxXNtgmyLSGlSyPS0yIUXB3sXc3pWkvDkEfU87FVBhRzFLKfWWzF7WUxkaYZy
M0FvNhZIzbv2PT5Ita/yN9i9RXwIoK+C95RUHIKRY4CCh4Nu2lcGszDJ5EI8BCrQ
fQjo4vMqUmKDWmtYTPxQzsw3n2qZ6dQd71WNpnTzmV2MJp4YR0PYIGilvDajx9Wp
5qcb9lu6n4WZrH4O1aKW7dxVY1KOM/nKIXdvCYVgvkgx7cUq+NbLd4/akSwc4Zo8
B02bhlPLvELCRKdA3vaElnZLCyZawG90JTflc7XRr53ga9vLi/YkdQBDmqyl0Z1t
/bzQS7EsBuLlEw9mUQHPFXXto8sAOpKShCpUTnT19uCExfyaGKnBuNcr1OikfhcT
pkwai1mJGWietup0MmHpRECCEsqD991IJe0OuqlwvBVfDYPpXz2cdXWv4EQIO9ZR
x1T4M8CBTVll/YSm1UBsTAUpHmCTkj7H8ziJm7YeZNgkWEoEeB7JuU6Py1yshd3L
lTgrpg+wVZd8M2GES4y2KYLg594ttDDPTj4GYlK8EJbFwwwg+X2rLK4bAvtN2uqW
+jhZXVlrJnXd+73frIsiC4iW4pb5c6xa0i9oYTmNTM7GxTnAVXnwmJB3Wlh82yeC
NTg5WjRp4tmKxVKlBYw1uPjEkkqMjsJRwbOVUqvjt+GQVM7YM6nsCv236xQxfnY/
rD87ip984Z2heAvgF0+Q1UkvslNjQ9vKidULQf4SFww5z4Hf1yN3sXInnDvfTgt8
npx86ij4MjPLR39vR2zY+agsnkTLxbCnWkvKeMd4KKXcf2AmNNo1FK+nSpZugpV3
JQaHyOJoujENgzACmg1MRFDXW7brdJpydwSzFVV4JMcpecnoUpH8Ycb1Ovi+BhpW
pfBGyAeb05zRWdnTy7KH+7jSo++c872W9HUwoS9+XjolyNYJ8He8s6A/Xa6VWS17
4kwslk1zjZLrEDilh+7n00WSEy1Fdjfefuav5xBkQQiaj55US5FpmHOLh7Q7kLcH
INDUKrKadp1sg2p0aHwRUqL/5fV6U/oFyKlwpwhz2g5hvOrpcESw1rlsDkzLf3zk
2OQu234xT8wTnkqYsEfh9eg+0v4utKKU2tmDEIc7PMgVLoEYlR24kS6EtMGA2Qqf
PHibkAaYVYyVrbh4a0Gh1QtuVi4GWLXumJFKiBjBvJknkmav3Y74jh3fxtT9AO09
qzrPvOTJTiFBbV/OWLMcgndsu0LnltFIiNnbml93m3sdKbNYBGDSP4Td0uRBj2S5
WZmOiOylOOxIY3c7VcIQVXWXY4yYnZdubhQgJb9enaNcokZZT2fzV2rSY+PqGzIU
K8STN1hc+291G8s+BkSKJ33cg78QPln6I8Z8jPvlvkgAZKaFOx6USYtDnr1AWENd
gBP49TeBF7GAUQAJVR/hVewVdY+kz/aDLFuF79+KeFrSnaxLEljoCPMuMxNeDrNd
Tda1tSZ4vZR7KfwLl6aUtVH7q5Qc1N9BoA1wSXusfn48lKbH23epPkM40cfepxlS
dMqvNv1Oqprwke7F/FIW/PPonACBQlKPBncO82h28NhqANI1RFMfJclUOxz2mPED
sC2p9GmhmouQlEiKvUtFV3l6JSXZNLb8RUPQTOwb2UxN0IsG6spRb652ufjUToAX
FFH/rWMS1Q9XzcKjZuPlRPQbmDRHlM2SKM9irdAwo1Q+Es2h20PFB4zzcsGGL+co
HDGSMgwmU/LPnMxjLPC1ZyyNrfDDkOPEOtn8SeZAp/E9A95HraRrsbSZ+22N5Tdn
SUyVssiAYHCyJfc0ty5h19sIFXBkx1/JF64cDkjNk7P9RY8g1g66UdG9zBegFWrj
lG1rdSVHy7IBv5mxzAlu2JUsaztpsd7ldecbEXU+1s5U6hchuiJ2/JeMdnUAsvOB
RWgNwYsxoW0S+RBoWf5HgA4t6V/1Pt+8iBbtj3jD6F46MFJzmctdyR66PFSG9F6c
ApG6R1q1E2GbGn5j2CH/j63SQ8h6Z5ITfAqtOpdjxf885RQQ4pVReTM/Ir7XQLLw
9CS5XekeAmcd7R/zsQztCz4fsuWR8sQYyEciJ9b6nJO3n/TA1NiEz+Tv7k8+nGgL
xmz8z+orJ0W3gsTlccsGUlfG0Vv2b59Z5wWaTPQliimUlFCuPpvabW7uvwFeG+d3
3/4SnQfK7kV0mCozEAeDbzh9JFI5mTrqja2LFnAeXpOu/NkXWdR5k9by6qaNR+KB
fgXbtYDH9hWKp6nCMpClVKR1W9lCVIDaGccnX7sm5ybEXMg9XCeY8W8FuiFyYFYj
eJaYUs6k88TmwTg1k3JxsSP+ambAQ4GlaTy9Bg9PSFh0gkz0nbIqiJpGIN5phPmP
nf/LFLX5GB1AJKI8Cx+x+UJU8tDM1WoR96olLP0Q/9L1EJZoB0JVTidtONcH4baU
m3/TtttBwbL3BiDunD0NM3Bg5UtyAceYPaOfbAf+HBFnrel8UNnIoO/GyxNFuwXc
PrZdNCX1rUy2no6OPZ5grdOLb/+vkLdocQ9t4QReQIi9eONTuSxESzchc1d4Rqo4
G0AaKctOqSZPdpyjg0tbs5O419E72K8KqrGaWYBGXqekigJq0tyiNscwL/GvLTGu
J3ELTITFFW5Jjp6liR+5Xe0A+zonzq1BaAZY6CoSct017jl118aVUrmh6ihmoiXN
sahZbJRS353BgJeymBd1AGaU1FWiAJM1rtbYuFBNT4+oenDcYEynSEnwI1Qlq0Hw
ODIsX6mAyigmruPDO8LE6xugO0CzhilZjGjs9j5FWcFX7JmrIm9rwSmlpo1wvGzq
ucZksW57qxGQ1HSzhJsOljc1LTPNyuYU3sLFsC6Qtlf25y65HQ7OgJQCycfh+Ane
ZX+pBKbssGmJOaBKvJOCMfm0ur5LtthRAohpZ7ncbXNA39jYzjd6HbFke7cXoRu/
2cxaLUtgWPV6qB7kpSrTQIcOddKCk8wLIwnk0CqjQQSzcWUWuTAKs86w4znv7U2F
y+Njr7aNo4GrYrZaUccIjQ9ss9zW62LflTEO7ye0c3lqjL6qXYMIM1D5UjQBGBtq
jGWntL+kcCNL3QdnjQHKhVuNscQtzj1mjVaMOQJ9ti9qRoJlJlZRyjf1AI5jG6CE
ahvnuwftxnIgVhPXbwyk3SULqOQjd7AzVjfDBx9UctQ+XHQnHBVcJfkHnXBc/1en
6LaIdqZIMfKvpDcdDcx7lEzF9DzaZbuCj43Ai8q2foVH2LT4Ul/cq5CLpsquvZ78
M2GQ8I4udvTvPAzsm+qko2q6ai35RwD23ungwE/axn1KB0AAIwkfiZNK1Lf7MICn
8yTPokJXT0/5RvMu3GSr/G+/Cz+CKJHm7t11EvozTkkrMgyV1aX54kKEsuOB6TZr
Kl/+Csg//A0Xasg9YRm/PaU5g4LrDXWucpnI9vqDIbsajpDz0KcKvGS6x25gg4Y/
uXOCTdX/LGdabAfDNclp2WaqQ+ZFJGjWNrni+7QniF0bpRweVKfCLMr4bvHc/6hm
vv4r6sd4Rg6LkUXodT2s55iwMv1IdcO89woeQ0kBnYGstkk5ecjaO9AZxyQz9X7X
fCUw5UEaojDaTl6ptjHX9P2qHGOTRyFmSdgEp2P+4vQiMXbdRX8y5EjLNHiDVpxv
lB1+tEQk6E4v++jcmAMTdJ6TKLXpo0IfXVEAM7pi9vjLftELoLRV+mkl8cmGp/31
xm2qdPWQWzLCC8l4f5Ph3pFkX4cVPPSIyW3Yg9Aqd6wdN2ptvvic50x5hBDjhNGW
ToEyQg6CRjfkYfm3AW2qhHmfNY04BJlLL1sqbFIebw2czfo7LxVDdWtefWE6ZYcX
7XDOiri4rtHZk8pbwYsYGv6yUUlGBCfDxH1Q8qPJ4F/51Y9xbkQjBaGvJLcyAzlH
+JZddF11alqRH8Ak64Q01b+lSWx96tkJaJ9thvCDKCfsO3GarSSHv/KEINpMnmXd
us0G6PcGsGpSNTglMvWuc/qaPnKATlQfjKwzbxH5sEUl7oq12Ije2wglTRkIw721
V/yChAeEnWTxWG7zXfj6y/H1ZEdfbbRIIAg91AOAEtQxIohIB1WjKqTdYGs4tPJQ
z5K92WhwtYykiSEZZnWfcTxSqRu+kyvpgpAtaaYYeswNAuFpRVcpcJExLMREHyfA
PJcV4UNxYGKi9qjZ5OiDEHd38DK9244T3Z23XXBf3SSZao/MleO9TqeTx9IEQ7c0
W0c3tdv7OBNvIYlyRHGe4HVmBZ5KS45Wem9j0t3ibZKYvw1zl9sB648RTBfx8Sqb
5H7YeVNFTIEddrJ/SQ7QF/A4w/RGx4AjJ6S6cUT/8i4LuB5tXXJ/Tr1MFFyPLQ09
59E1CPvPkbBCzpkvI1e302oZunQt3Ytn30SlokS0TzrJYM402/S9KnVEoAfzcCYm
AKSLE/cl9bEH47tx98UFf1Q5lM28bivu/sQ/WS7j8FH7BPRD+WrzmCnlIYM9MXzE
XS8wp7cHnRQtK0M0GAR3OBik0NMS5oXWpD2f9loOgkMRL19NxaBfOF2cSFDqBiOa
CSQmf3Q92B65tEQ3dKVsE4x03NhImgMZpQaYSRzqIpC6pkOlU+6gqArdm4vCG+pi
JfFWGmfioG7Zlg529Ws2uwJwYd8onXZ1MOE3/PPLrQS5QRxlvKDcN6JFGPj6/jHu
1EweJPKYNjwqwGmmCqnWREW/esRM3oiWc6hVYzIWXBdGh9B6QZjNPgf2w2lBQfHe
v/cxf132HFDlEByHbaLoFCYF0qepzQ/1fWKdc8e0S4L14vkP1f27idtqLwOh1IWK
1MXbls/L4U/rAaaTnY0FPBrnUQOa3OHP5vFM3BsHV6z42xW8nUZqCrvxdT9O8MyU
zTW5DGaEWPS35PEp9vtzdXo1VaHTwt4Omyb1xMqfBvwLuYAYBR/j7xFdboXM7EIZ
7GHDYwB+DYx/PHV0a+cTdUTaLJ4aJGYXP7/RPkKBuWNE4kZ4Uk90iZQT0yta97st
CshYqxOtB4gG/pD2s16gmnRzWDaQf5D1au7AsOo1BUr4FgCt/V2d+QtR1LzKuKgZ
Cv/UazUyg+bVSMiMX+bnZQd6lkbF2fY8m1prt5lOMLHCaMFc9N9OpmxOnyriuHtF
90nGrCsD/u0RasaQNHboOAh48W+xqQqEbWiw7yf+O+0gZyO/YZvyyWFyXUBj4WCf
VDZouKnx75EcuFxQM8gqVwVcJ3lPOGvDX3ADprHBcsm9PW/5ZwztAmtFMM8wKMRp
JNR+ayoKxNLRaHXwZJoX0EyRERLPCj4952OLlbrG2AurGbmmOdYQZEQdM0TfyjQL
6kpIr1Vad/mbuDLvI4/xvU3kNGhS3UjY5IH9+NW/boM6r3C+Mjzar+GLpRkYvczW
WtUES2s1uIeXwIxKljRQZhgwcKoWQ6F6pdNQpFRRXJLkX8tM7PBUXklECJOcreyK
vDV11JGvaKDYiD22xZyGyi08d3M6N3DLFmwEHV8XLJ3QKcdQ1Qpk+rhPdtf9ZzHK
AYn4cFNadp1lQHqvq1ej4dBLsoHwPXLDmnOAmIqU/m94zh9r3GZ/CnRw5Zp+FZGl
sG+XfK/wwH66a/HoZGrssF+KjNNSJCTiqRFoPt3I9ebqUEYB1o66CMkhDCcupUFf
mWX5DpcqUkv58EqFWsqmF8xGUPhdXqX8NCsESaGiUktZ7NUcXe1LCvBFnusRi/s1
01AZnzsPA2CnxSr/s1u9arCCnsh9DepQcZ/J1RilPoIL++lPQMYLhc8xB8jsd1tY
6v5SUzE8k/XAj40aH334JJQJ1qItyNtMMlCdWz5GcTCNz+ZWOWtuoUwLuIRmQ9g9
W+iKGgraKgWe03GuMx/aPiQbRT7t+waFnKqgcX6d7+2A/QJDAaCcDmuWSy/wtg8/
WFU6zYPCqec/0jwFHEVeZHWUEx8WXVCGbFkIyoJ2fc+geXUXhGEzPORXWL4eoAuS
bAmXHPO2Fl6ZnLTzHiFU2bgutSMzO/G2Rq8SfCDsUjqrbDODq3LeWTVWFT+C5dul
UjPYNj3fU5wDylGRlkVk4LSw/6pG1wRAS3ikzL3npgRKRPledLGPlNElIh5tdNTS
Dw9X/anxiIQwj/1LMBod9M71eAyy9bJ4R0EF14p59U6IJy7ehxSKBSwX4kZXaVb1
uAucJCpeItfA7ZBmWvOkBbEHuvdy8XIHg4USb1+uFS8RRl9qy82NHYjh8DAwlR23
tPzNStNJClum5tHsg5PVsHQkAUFwgMoAXvDuaDTzb1uLo4JshDYAwqRxZYSKYccq
pnVyqnzi2RZK+jufXwOQ5mletBYyqeiy2T0eiAXDM3BHlYoEuZURvkDntU1M815f
9EwJbJ4uMdxdFwWXAlI5HIn6r/QbaEckMmGHfYlTZxUMUuPICOgd2WDbF77cHOg4
XOVTpfouvXkiGCMrKX6KXM4G1CtozyARCGpZaDe9U3OlB8GdMgfJPMBOByL7WoTU
0+9Esr/lpAx/r/l80wlgUS41bU64HSALhqE4lc/rafIV5AVkgp8zJsQmVXzp9N1z
mkRlGaIQYtWdKDToYJZrWAHNj8S1cAjTjCB62aWRwIru+/mZvaxbnIT4/Lv69n+w
1WjCjqwStrhruc2bSLXy9zZFIiH2RZ/7HauYTDCCcDIvXpkJI/hFLqnN3+6mCOyB
rt8Gxb1DRchJB9ERHF7WRrbUrzcXgvnBqLRfW8Yppjg9FmmOui4cGAc8PjKUaKOk
SIGivYh0E4TTfLz1t+6z2IjOiQayavVyM1UwfO3GK9+UMdZ/svJfyVvt31zgURzU
qDYMtKKrrCKOFDsBokh/OiX4fkqaVS73/b50gIW4Kibd8QZqajNGzo0W7kEKR+8C
Efc9ZCoQ3Qb00HCpB5xHvHDNzNpziLsxHwptdkOPQXyOEWPlqtF7Q7Fkaa4DQWOM
H0dqQ1jE2RsuwRABIYDYVBuh7L0pGpjYON1cBYvKGG+AFZrYH8iIlAQm/d1RYXDZ
5U+TJTQJ5NY5DVx29OTTbXDAqTK7sQDns0PrHqZxYzlqDInQB/3Rp+gCR0+bFzjg
R2ElnAr7wAmgDFrdjGpJu18KHQxSVotnkG7CNYERD3EEhOTplRKK8Tg7cqxLYnJR
Z5T6Gl8LqmCsjQwk1IxfEwsNk4lqkYoxxblEKlbnOT31qNNvnfmPlqzZGeid6yG7
OpaJ1HKro/wQzx1BF7eGpUiR6OUrNnFZg5cahB2JdesoU3DU3iQJYGTY8uozZaHO
3l4A+1bfxsO4wE/p8SRO06Cm/JYCbpSU0cR39AxigLL10s5+FSb3d/pk2DFMHJ9a
jIu1gjwkYpR9nBX4u/cPs5GYtWM+RPkybY9mlioRKBs3iOrd6gW4t5gHf2NyaDYQ
H5jqTur/xSQDicIUi85aU7HO5yBqyoTvJ71FX++Cr7+yJpdZWyd8pXq/vs9I3K+x
nuyhgCYXK57/S0hMZm/Mp66I2uO/dbkVXTkA9SD+YHWo94XPAixQEHd9o7IBytem
bSH9IDSMoNVVGy/tJoTbr77o03rGPSFd+7R4/0eQuFu1R0mmhsli9ssqgnI+Vnze
CyvK/+uFXzS1i1EjCQbWjarHsS4C3keNsCrpz6OTvL53HutgVxMRZX7tTuNE1qu7
1fIX23+VsYJjdGdZ4+GjuVlK0VV4dGBhCkhmnI6kG2hOe8uOysZsKj/YuuLOVA/H
rrj8huocdouRUyjyorGLA82ShWG1mlz8AVILrDZH3V4l2pwonC/EC7ZDaUgHfnOv
/x+JZueNSWN8dpRZeGqF0N1gZ4qF8qo60mp2cq0iuKYemeFubJ1kOyUOfN1AwRsG
V5OxGm3HZyW/aDEz3jl4lDr+nwm+zvqkuXPENjOKUTis/I7x6j1tg6gPLFaRXyxE
4iQpqQY4+pa79hovBzW7iY2DGLUS8UQR7LZlG//fP9VUL8koXM0gJ6fsNoTStslh
oCUCqRwQ6SFgqdnf9zIt77ZSB6HVD+0uzQLKe4u9Po7D3oRdXxmogM/bDpCDn6x2
QRek//MuQDEPCaQAoLnvQO6uB/0Hb2/Y5qbDBLZ+66JY5ekARXnObcfty3rDMC59
cpONf2LdA1xXPpWoolQuJ0hba9cYrJq/5fe8124sTDcnYdPhES2R5/WBf0yB9p0f
dngw8owczx2XV9KZKFYXCqW+kfnjnbA/2YBupeGIqFRhgGD0k82cAIL3MnXErw7S
VqY6e/H7adpvODmoF+k4O8hpKczQxGIF9ksoUnUfIUTvdDzz0242A57exT1Rgnvb
ej7o532eZrfoXqyootiEv2iwKeF1Jwk/L1xc8QQjaG6ITqiLjnz33Dn4Btou1Bh7
gfZl5BQefaFZSzwy+0gZKhzZIGuY6ou6/nApbOquaSD/SVR7rA2ESNmzmz2fu5FE
3sm2MR4Mp5N9FXpIzsbxovqoujYifmFBBhvQr4y+2NTYidI1VJHQsfpJWn9m1dow
mro3zDRIHLDNaL4GAFWpewDApccMx07lLAjFlMr0f+fTwtARtLyRwVWek5ywYkPH
8rY6XnRXRAnIkrfDbskdhnz7m3D5VZ4I+zP0YH8O1GoAXnztAGrC7yVUYPHezSII
hXCMYe9GSEgSMegdEMttiq7SCR2DR2vUO2nunUpooGkpbRR89sTua3NMFaxdNt5T
icM5DVIYB4KkSTCjCbSj1gzDE7o/zXFCGH+t47ca+2jkVWhoHCF9aEI1RQcfK8bY
8iEgYHF0xTbdSyZixGB7KJyEaww1cC/AIU9NJpw1RhEbKE/7bKmXZ0tenRbCD5Xa
eLIRvqzsUjJAg6elezjpEAcUlgbUyQqQC7huuJpX3FNxfGmmaMatnL9sjotpwP11
2CN4cZ/7PPkdMVufwVGj7x0mScnwVDX7zQTKhng86FdrOTgmCLEjXZBqV482e9zp
L3HXpJGM37vkKOT5ecnkS+5DtgUo+BnFPy9OKAUU+6FV13ZQKnYRdE3T7ucNc5VV
8nI5NYlBFt2ybibSBp+CioXBeYFnaRUx/GQiKPXTLY89EfalWuZumf3mLsKfT84M
nGozWGYNqqyDpSX+5pQa0U5A3xQ3ZWMWmAwhB9S8/Ly9UsU56Yt0gBKWIwSid8Ww
yno2zNyj3Q4tKXt/PVOFhMeIW0PnrRyzRSryA8+kas7UV0TAc8U0BJ6TNVOurBfA
/rY++HgTWgRhajPl13Gq9M6SCu2wAyvxGT7nUCFeu6RZSfT0lgfw9IMcMowRZsND
38R2Sud3eh+kKCX4f2JDDKK34SDjTKL85SOzVWwSyk/aYAV9Vc7K/xBf8WjTkzTd
JciOx1FKyMrALK1+pPAzubmFLj3n4BaijB+oDbEwemVa9PEYCAasyjQcpa5Im7OK
vaV+KYW7lk+4EaMMOtrtYxDK72BN7LweZCKv1ZUp2WnDrJQIo+LFW9G0DI79zOsV
FGscDMwP4DCR5IhvwZinCsnS0dsyBunxEegfx0EzCew86SXLNYf8wCS7CHSH6lT/
99sQQZbBeUcg4lPwt8DvveVzcgullbdfN74NhnU8kMmKl/YkzCmpkYA9yR1THj53
tBfp9VLbhmVEClnP4q4NHIutuWnC7jiEgpGufuA7Vl/Uce8DZoaoSnj3UYdEQZt+
G1Tl0XgnD9g8r6zUrC8NBsjN0YyWEwUtYLhyNHvTiQhqDlKiKG4eBBSWaLQ2sFUM
vk0thcWE0lEHrsN/bP4qb+/vLqUHwAidD1KdlnwPhmUpqctpU79BS8kCyGPZTluU
bDXvMmvH7Px5S4Hamf/mNmzlFGpOrRs61XCrfWDDntnHDPakDEL9x2D0GUmRLpgt
KlF0Kkqrx/n1ZL/4mpBgqo9ibTYCynLBPWK2pu1sW9+xLKRzeSxI6pE7dKEJxOYq
zYe1YAbMIoNzvJHkFyd7ubQ+EfTBHrkhpy3FZtdp6/dlVXZTgnnPh2GoydNwjxZN
nj/8Pz4dM2Ci1pdNLpKsfldL1J2WvFqwh2iynNu6xx34BnEPeBgh4KMqlI4BKOiF
3yHkteqTLm26q0y7/3YSbxl771HQXF0CwG6ZYgw14JKb1JiFKFRC0IaVKBHg3fno
IqyWJEaFvJ+RirxoxFJPLtHj2ixmRz03mkNrS+d8Jn7/09APejd2+1RtWOiXKdNb
Cduo+7Wsdsq3XFLhJiDN184FLqwb6JA887ExD2OQeHETxHcPGa5SW6QPq1Ie6UdP
Cy3BhpJKLSnPo4tbJpkEArkb+PUBDbRIfBCyZ7FVDAMiekkv8evk7NPgpcxn39fS
IaOs/1cHjAUDFJZUYpcvwjCytBwpbS9avTirfueMNU3VrJnZnTEGrpVaz1uKAYwr
6iQpx1dtC6LSkznaMLMVqdIbJANXQm4uQYxUF0lhugYmCbN2uGr0cc9k5rQ4NZsA
mLkSnZCLziylnds3fNiGK9bQyhIYAVVNxi3ww7009ax1fdpSDfhPnvtS9tDNLlJc
Lc6bmtbMo7lb3Oaa/SEDnU8/+ozu1H6SM/pByG7rcw4xNwj876MaRFBT80NIaN78
Btr7YDIPstGUE7FTHfV6XkAyLBEY6rRxKwTifgR4eFRcXBDmGyHITgswjdHSsgyn
pTKj3bUQ4/ujEOHrlhi3Q0UuIfQPWSGvfm+6sJv+eXAYP5tIh4CKYVoYfr+g3MeA
vYh8rkD/2cWym5phSeuXeJwP5xzECiuiYYAGmk5gPIvgwv/2n2TRaaLNCwj7gJtM
iKjGCKRRItGJmZWD5Uuk9TQjumZy5AYwl5jJPntBu+7NFbW9eHO7WMWdeBS+Ev/U
p/JwocTtmrHMz+BcRXRNFehIfGgmZdw6IMBIh0vOCrdT1eGQMuvUu0O4FVjLz9i+
Qlkea4QpjAzuIQJaQdKFE0CrJy14DTs4Obzbu80qnWD7dhP9sbLsxqqLOjOp/DLt
5SWa1mLGf/BnThcEfqF5c7gFQ0lMoOdOCoa+h4V+2gjC6QO6j+6qLGWncIVa9mhZ
holiODjDe/+upfDBQ6KeCmtEQetP39zMn16IIa/T3oIYEyJ3y6A8e9iFCF8tXvbD
EXUqGUPX7Abscs7bMsQCC57ZxXeXdiuiSRRUusNF38BXGfCC7WLrX2PfUgcL2Vx3
HyPWhkMvLOIrTnAmA06H/B87ou76xJJh6dOL/z4W6MsUtZURSuzmOuFegbpTc4QD
mOsRvcumxlHIktjyJIaBL2DMcsgjmcTtACDp+j7HZf6rahMoFW3+hPLklYVacIDq
3tfnIK5X6Te0oPTeET4XYKCVQLtG16o84KMyeYiM2wau0mJ9QLMXPV4QYzdQFonm
pYvN8W6SsW4Yq5PB8SPnfWTRQilk181SZMiBgCwJay3wgeEy25zZLuHwqZw6ytzl
v3PyeYNHCeejx3jKc5V9AKSG7i7BK8gSMUGn8Lotfa+jXaZo19K456QZSFY+I+TE
pNln/NtTgC9+uMUFstwjUcrS4wR78DB5PyHgAY3euwLTwoBkl5mqidLbTf4qLwXa
88dFoOYleJonwb8VdNnYaQzibfPhUmJeXyaGNMuuF3dMGR7qA+C38Q52lrhOWqz7
RAw2o2YsaAPWK79P5aAhvAtmtzZUME3J3bLXEjKpUmfm9Dmmp1UIWCPfk5R2Qgnp
8u1b1yEckMz94mH+mbtYguhXd3FfMto4N5MCZMYQC4TLj+dAZkQwV5PkyY4PxW0r
Uv9bJVYQDQu3aAtJ+rmK8DScHcqjw6C/yAlMjwDm5epLDjuqVXida6k950ERRNsI
BITYUlTPJ1gw1b6ILTxs5EQpz/AFjYfD2XfzbusvL3AXDTRwG80CYM/1/Xzg7z7s
AMqZIM+FVLzE7dBCyt4RcRcVZPQ9qZBHk4nUKSej/gsonZavvCzbEIo6CSqiHXuy
51Oh73haknPraLpJ+r2KCsYPg6pyaBv53708HQq7LtLJvPo3vVkouZFWYNFm8y0L
NEmZugTwdkNELfQIRBJK40Z6Eo1ymO4NltJCz3bCL7q3HWvB2X3TvTw1+ESzVipL
sIgrfoj2sXzfQcyr3OzEje1bpYhrIDUfWQBSqdvqKqj/l3l5a6dLplmhK2Snd6Da
C+k0nnhDmVhSAj8mmkhP67vZ9BwOUhL9Rz9aJPHvj/zNwCYfwKo8vwNxzMsYLwt9
CEjvbNcJ8KPavReBK8nm5FIj4v7zXSXo5A8HQ20D1vfW2TiXdLD0Gk4zjo9+cVP/
EhR4kkJIU8y2GKdpzVdys+a60ERFSGKChPhdBQk3WqDJqzcGLtzlsZtEyrSB4Koc
f2AipOjQPeY9X4NtGs5TXsJ09ZxBwKBeveQMrIvw6UsZPWBuJKNVFSkGGiNuJRvn
TdCqtb1Ds39/gkNUl99+OR16lnV06GZ+/CM+dR5O041vudnj0SE9gZMiLAhnfvia
UjEhv/7BUb//67Pb+c4JcfgDmJNijJ6R17tTnEJrA+RoSLZtz3VeSMQnuNoNEg9C
1GFhl8431CFbuo1uaI2qKiC4pmIW6Bx/rQouXb7B5LfWndSgKbsFHPXeUG+pSm2z
Amk0koLhCqu0NYkHSyY18sWkAsHCWaVjpqaolsFw/9tlUDhgT9zyYxJlzwSmGAYc
tA/Y1FU7/PfFfIP1ZcHj2eiC8CaHYWl38fj26o0YXprJMwfvdBHR/QZEYrwuhFcE
WgR1lWBnuaa5cUMWv0eSuXyl/A5FNWTgqfdTAqHn1Y0oj5hnx8ILX0z54h6/hx0R
wlLWI920hJpWJ6Rul+2THWGZmY5i2DELmReyMyR6OsWS438it5WYbuwu6jjdk1VE
esvPqRzItYWnsxolReh1cdUgN3A3RwZ9nEe0/qr+H7L1cQCTDBIvSJ0gRBdAeWED
UDaJcv/P8KVK2+tDjSdwLTHqG9qy+FrltI1Ueyy9SKTUfEUywi4p9znAkQUAQ7sk
Zya7yeSNVQFw8+caa/suui2kBfzPDlBjeAkRG2C+Occg2lzuTk+uCklw7rCRu16o
ElxT4E9dLN5IKzEeJgWfyTK/5ei3UafpjuT0+X0rAyixEur702uEuKfTDap2BAib
ZQfmWQmBaghY0yslLndnjsc0lC8WZxxxYgO/WDsweOl6N4Atqos5dtDF1eOUvWeY
0xyJvos4Gi5DBOGAnbl7KkNMHYTcIrMA37k/7dMRYjiGGAj8n/tRK1MLkvGBp0Bg
3wu4wx/DDO/BM+YBv/ZQruXrlmYniMtU4rnJBP+LMXBTk7tkBtRzZRT6NbSsMCwD
49ZLClGGK8k8fnJM5XIHhGAdLC71wwf4Rmw0dImd2Rwhl/Ihyc5HLMWVopeVZnDM
ir0F7AZZt1VPDlHGD9u8TtRrRGsgXSch6m7P43RxYW0jB4r1ssDc8fTddbVXloQG
rH3dHWpwZyl+TeKjA1RfSCRFv2tA64HVkgVY+gP8+AY2Tn2Yvm6ZqHkDnVYylZho
Yp9Htv6gsza6H4mvKtCd7AatZSFEWZzDFlhiJxn64kW6T6YapG/FPB3cBpELHJWz
iMSlplEfpc5lFzoJQ+7r54Dhr5W0CPAHscDfMyR2XL26+okj1Gz1PBRQ34Ia/Mv5
fSCaNE5bvaeViNZwRavj6N1wp5wutKNn6MnyszRSVouuTbkHOHZMghKzLEAYTvAy
rCaRy4iSmadPixLtQGtZC0uiMqqp6iuJP3HKQinqgKlmRagXUJ7cM9ZrmCVqLKUU
whCmEJhmIzT4cnEd0QsNefnIlt51ROUNqvlcsejJWSYvJ31GagsE4ywCq76hi9il
I7lJ6eciPwYhUjnGK4cMCqpcFv++3+UEXEw4+//1wcJFbRZ8eFPsXW1rAYnW9/Pu
WG491n9pHcMYj9koC3KgFvgCsfiD/RHt9EXGeGoa0qrOspSuhcM5ZeNelaf95YOV
f5AGv9jWS+Z3785QZc43D5EO/tZouazC/cbRB/56SKtIjLOBjxOZaU8cIuonNxfE
8AnMGnL28hE4HpcJzdf2g76cnt3MzO5Yn3AGcLZBjOSkH5Io09TBtK/8eBalDNUF
eFlCeabyh3HbtUAp6FxoEaZ6GaJ2K9r1oWMWFO7dITPxxgule1JtJzATx4ftS5N/
tpDn5K5Q7zg96T3eoo0yBZWcz3UX8p0nN8EdjYMH5arelDoF7P+Nq0mpuwMulvrS
e051Fpb3Lz2czmcPT9b1KucYptqmHmXwwEEgUF0xZSE7QDISiB/qcCMiRzCzkhFr
bBPT9eQh8/P9tkee7FLqaUKRdadLVWwWRIZGMFsjxVV+hIktPjvxlLKRlP1dIwHG
phYXaPHUPXPc0gneSI6QZ16QS/kL0I3W/DUOgqzwHY/kjELOyOiTsLxr+50++I7r
j4qKTl/xV/j0bymdLyB8dGcq/slrMD+Gay9/Vpe8MzJlvXvnU5zVpwtUuMB5W5/U
f2lHNytw4QkUEcIteLvavGU9h4tVFnR/JubpCoaePqdV7jExrqEaGux5cT4apTd1
DvXldCXw13+Riz5E8VTr5RuiXv2Db88lMiwZFQkay9aoOy8sJc38NagTgOnSpfQF
SU12HTJ4a1s9tBKNUD9n4aeKPMlpp/wfG9nBpE6J24khBPITiT+UCxLz6e27Uvf0
4r1jrt49VC4ouNe6QmSMsO+mkzj37d6OgrqF+QIKFayKKuuGBqKvT5grJq8Kp6mJ
y3WPbuYtUHrNGm0c3nEW5jk+l2NbuxQ04agFBS5s1VBYCpXGh9wR0N7wAkUxWEyn
Mm6GleMACyZBPz7OVI1JR5XJCJvU4HyEACTsxbt+oyEFDc73URUO3elonyNlpoEU
mK6uNf9FpZoCqEOrxpmvwMKysXGd27eaRN/IZ3VKGdEhpXi6gpUUrBnZQxF0qKor
7UmlOH7x07fDqfAMYfRd92JYqNcxtzZv/KqJ9YiJOcPUAiFHr1ehsupXIwqU78e9
zMe6vhiKtzxmjOL/ri3XunPOFi5rJdaSwf+mcrEnF6BfIHqOykr7qhrknfZTYvz5
XJ4/X83ueAJcunrQ4nXsHSSnuXT0atH/kUtW22SObHm+t5mLlxPqjIDuxi8/hSNF
0OC3olL5CSqmdeIxvYdD+YV8ZjuH/6RXrY3FF8J0QtXWxugCNjMUINnY8L9J6klD
7DguxoGK4twEy0is5EJicreOKJ3uaDlq6JcnDmyyEoCU2KmAJXDauqR3rpBxyxtM
GZjCuvmNXMdmx9R856a/qglbpKF6o9yIvXIUN7v96SRFsk/P/iuXGnMrdKZx63o1
LYKkhVaQxtjfUCctkqrGn0rn81hDEJVNoO7wu4ZwFRW2dilf2bp5B9x09DEjW0wf
5USzFZPCclIN8fePnY3YOak5XgfNsiujLFXaRrztsqgCL5rYdpp6TDmnKijb4Rs/
UL2he8Xz+IdJMEzeWTry6g0NU7FVw9i7khvmGWKf6mWx/wMbiy2fA4APbQ1Evkrf
K3ZwEajBDN2/Zr4nRXHaJQCl+Z/W/21tgGAq20aHViyc2MbvjYIcSbUNeAleHSH5
4WLMR26EtVK/NRdMZw8PbSdXc/7PqfnmB/MS6q01LWtXINeun2+xaSMSobgfu5fz
lZft8paWWfVjI54nGg6u8/oZZDl6R81exsa+O7SdrHeBex+wzr2g7cBM64Dj0CMR
3t281ZNVo+vTAyjYJludtahzWfxiWg/RQdiEtnBcThrxJOAOhdYbPZxTNysRgf/D
Wz+j0O47j/mJSghrQ19TbvyiUaEk5d2THbN+N1wnjvdd+MFhOiCzkqIwvazAtnIH
uzcd6fwuvEDwxUyklQ6Stmq/P2G2Zko5yB2R4YP8g2UpvscofyfCCSrA1+kyRZf8
YG/MQ9d+YPIBk1RGQNs/B2eF+ofaTarY59YpWVPui39cBVy+96MYJ284SElWpMA+
zHOYSRYLmW1tzMGrda9oMARlIrNoEZzLzu1VWulx64kEZnJq9hkLmLfcUJwRTPKn
lnS7pifdj71us3071oCt1s8eE9/T/tbTvv7a/CZ+x5/XZlo3zMcYgcwUwiWPT4eu
SMk+md2Udx7owk4D43yRubAePW5WS+PRe/pIuRf1zOLsMh1juRm1Tb6PgVT80zbu
WDpWR+mJxxm6/l5c9SBfw2owv3MrhssVk4qh1m4J6aSHrLApYCTBjqhMwv5463dH
BeuB1g5H3qRZwREcd4P1H/FY97AtexJQWNdrqpmcR35LhpNB4xTShQJexyLveB1r
07+ZCcU+Gd1H5BSrUlGtuTHwdxdpxmBbjTMDrl+ylt7ACC1ghDlq5TwQvOj4U4Je
E+MYjDKBMP7pyaLqrHuN1Kys3+LLqAJGHUb5X82lEDYVauM04q1dwID+hWq3YpYr
ILC7Ydlm8fsAMT00ZfGZMVaUYeOkxWpT6rQyDbZ3PtguBRK0LWDEgNzt5/Nc57YR
bECm/6xP5pSMTymxLS++A7MTWRYfHDvYCh04Iupjqsqmyjzej83lDnr6ZfVL9YGc
NDzDZLW6Jav7AKTzEMYig8onck9Yuhx7aHdwCWy+Ha81gPOcHA65+ncM8wj5WCT3
iP7QVcOIA9s70gRe9HTFH+9vaIzP7gsQ/+N1I21MCEsAnAUoQjx+l1IZXU9h7IOH
dnH0iFa2wZ+QQ2udUYjknA0bVCPS0N0xzf3iRqH8gHdxK3Sg6iF+DefA98T1UO8k
fhuDigHbUyHBOsVhYCCiSTpAf7jAbu6cWGzyU0IMH0p5ZPF+QQzD9/ipWs8PkSgI
xLHIdRXLhvb87Xks06ZWV55NHZU5WZC7QDwF5Y8njnNphvRHQ7uzYuwM/wsTOB7X
NCA5nnW+UhCedYK+TjqXuBB0W+vZKrsw/9PNxf7zLZbQSD9CRLQ88IvxZGK91ef5
x/8p+N4GukTXBBzR1+rm56zAQbnInNwV6ONINQK3kXYPgDMznXbpXNpDlSNQG5zk
3IMLvjv9jyHG5Qh7JkPAYRxXOEInZ6VypElcmG1gehlAqfaQoCnRmmEKLxWhCavU
4IKY5gf5z5laU4g2cz4MhmtyMQJoVc277AaORZM30P6RtbXbl+ws3rehDpjfUCpK
QiOjXvzo3K1k1wOIPkQ37KiWOJ5K7d/uvRWhOuQ5nc0VjIS30RUkVhPlnSOc/UpZ
a3DsA1SVYNuBmqoyPwsuLExlvx9UbRFlQG6ijSEyJPF0lM9LpLGLRM1rvDX9q5jD
xp8QdaCvHPQRArE2XtvbLqXUnOa3JKZUHB0ULKHWf/ah3uZ2OPdjRDaHVIJozYfZ
8utCdjHZUrZrbcmJCLjh5Knp4q/iaMRG4/PDju+ttXfCJiso4or0Vd2e+qx0DKBH
y3ky+jWaoklH2cmHSxFqnkDKBCaDOigGPmQJLmVpF+bYIuZscSxpWiPmk7gKzD5o
afwYSD/60xH2C1l0B2X4CVQhTIEWiVsQ1dRHVbZQQbc2ELYuZItZFZnvvPp6rRcz
xuspd9SE3PQh5RDLdOTEj92+zJ6iCrWTpTgxg0/hsViOf/PI0wKi5qnZSboGvNPm
Rwx7gQHHydidhwzIR8qblzX73o4322s/qdc2n/dOsxnketJt16epkbB3tgZMIop4
F/xr6XdgXLjJzCp3mHep0RkUry/5yvLwuXWZepq/m+uh8x9SA+HXYeYAByTG4rT4
rmP8agmFwd6uFmc57j4HFexZ8bpjqMlMlO2NBKv9Bl3bj6Y/s140yZAETssyxNkC
LLHaGcGwPTPBeL4QOaxbqtCauKmoiTH76cOozTLkOaSOwwXnJomNYqKLj/R4Qakm
/+x0nexUMX9bi64UAUcXE3Vz/qzWLrr+V20Pe//4ryrzujVvEc1WU7md+ctUhzOu
BdkA0jkquqVF07qnwmoDVaGSHWUIDEUyTL/M9TqCVePMy+ClkROm47VwqProwkpa
oifPcmHvptlcxDPMnclUvPmN+fePvWsk5GnMYbm8wdVESnhtcn1eIe+4XIGd40yJ
RmLPUQf1M6CAOGZSM087gwqIu7FTLdisLwW1QjFBrbbYhgomxqT9a0WT6DeETrTF
PySO73H8B6+8bvrh+0hPanxCQuYFC8iq4Y+TxLKr1Xmlo9jPbYHlJ5C8rgiKtPTh
KSX2ZPIoWWXmJEeP2tIfF4sog9+G7EOgqeBUTDEXKFKufrRnM0J4vY6UgqU/Rcel
OBkxVePF1UA1DFRshAWdeJM/b8FHFnAOwoiVSQDF/ZO0kIhuuV5tJrBHmysERMz7
L1GjVRB9+X0wptTLKrSY4p+cpL+Hvr7RF09i7vni/hFbjRAsNB9o2Pz8M3/rfHg8
GDTPjxKmXeGzHeB/fMx7F11ZHeaGO3sawLcupN7nENXpE0vKeHzptc9o/APkm/81
/IfQ4atqg8Wzj5kPqKqxn9C0TWVYHVxKjABlIyNYYxjGblqq/ynZdkHWdNtN4bxK
l668cmpKxSmwEpDlidTciQksyyMp3f+ynry5wJFCnuhJLAuNqDuCl/ADicXE0SvQ
th6qGFaK+4kPBS9PleeeKXWmEEv/iKtsMyjF1/fYKrWLYLXYSNPQyWSCjUEuUbHJ
yU4eFJRij4PCOANXauQMy6Vf/k8FUKScvoqUGKv+DcdIEm2z3Ld6uw1IwBoIcWVj
O3E03vApUK1qycCcaDJa3clGbZGkAJ9Fosy71nv1ox79V+ej3gAl4u77ewg96okh
5H/NKJ5asZPk+ZaXvrAUeMyBAJuGL0IlgCeTgb39kHOm4tEjCS0/xZMrFzPYzCjc
mPcHC2yWx//Y3JH+FiIHL8HXDVRyWEEBtmtdJYtPLdJK7Ntjfjgjbp0sKI49zIkX
R1t6P8ZJ8GQeyA6ZNcJbWpIkEospZmzYfydzHSYWzLC/vXgZEcdfXZHZpjLCWK7R
USjs5ZIM9+bGHpqw8nTDzm2ABKYrDgLTR4IDdCgDulsoqahDswg/TrkEt3wd4qH2
GCpu25bn7wBhdERTqR9b4qblCIoTSWVdGIzxYto6ynxM2VjPKDWgo6U4LEBQEW7B
VlSWYkfUAJPiP9DhedjGB7MzdkvrTEdNcYiB33/zEXYCxsOFqLMjLebln7r5C9eU
stabZfOwS1X9VVcpCLjAXG3c5tz9XAu40iMr8JaHnJfUJ4vNgdewGRdnkQ+xYp8s
PXx+WXQ7JWxuvtZC9ipFHawGmVX9g7fQ4jpfA60EEw9LctqVrJisYNHOAU960zD+
CIwg8/Cdx7Qufhdq4UGtPI+TVnqh15gjCfz+vLQFeV6uu8hBr0YJeiU+Bow6vmQH
aMqXo6eSBgiE/RlbIfgowsHQKpA12HYWT28ShOwlIH/xvrYuYYpNt5+4oeJYr1Yx
m2iBttIMw0r3l5LD5691hmLqmSS55qllnkcsGk3vr/CmJ/kbf31/6JewthuRKfeQ
hQj+ZWiNxVcfLJw+DsrdSmhh/dnnJQGtvm7Hi5S+b5zc07hnhWpnpiMybdD4MUnj
9m5dtQjUeCqKo4oOVUkYbUXTzr6YZztKXs+2Vnpx114QO5Y3JpMVM6jHNVxBrcDv
14/qLYyMJGXs2XsTxJpMXp9oenAC7MUBn5lQLMSDXLQsVIYftCBGxdZKQvIyPGjr
8l7RBExwoRm1n81avMEFNDnbfTKGejKCtR0aS5ejB1XUAgQirXZtewG0wYook0uS
Y+N/anDOr0L6d8mh2fuo/QvaRpTBE2jzqhdQc92eHY6uU4mknMuHnTRFG3lS34Ro
t/ssGxNW0eB/S2Ym/t7IYmU1VZ6lz5AcxlWZZrU1Y5N6FVDQi6xv41BQBlEW4zT7
wTlcS+7xKd/3mTA/lOK5By2zRnfSAa7GtQSeAFSstUrnXeAPnl/wDEacXMGQg2vN
vCKXKiI6wDkQ/5yo7vXXXI3hpDpxJkoB0N3Hhcd8e4qwKKm/h0+5GTgmfgakqwBq
DaMqTf+l3tBQlHBjgYJhBEnlHAdgu5tkHdLnc/xApHTCY0Wb3KziRyzNiSYiu2vg
yK/U6hboh4oxbQrgeYmxFP5kjcFljRUY34sAHWYddOQgw36axRlpLz2yKxOaXBL7
QgFUdaDW/ajBQ2V7r9fOrxMGy3f1JBAhsivBfBBb2QHqTFAx2bFmd2E54OoxE1LE
znmvQt6Lt3J00364GDqvMClpCaGnzracXM1pXkHkWVI6SBfuhFeQjA2jAiIzeUDw
uRrdxMksY4vO4+lS9Ysn2o2UoykK3op7DweZX08WUyG0cBUTCVypxEwTzA2PG9b2
FmKBxZe2MF7sbDvoqeaydODUg4SMx8JMUC19SDAEZgsiOuig2Fc9sHP8WFogv+at
E2cqhhAyXWMr4n14Q5N87e+OEj2QOPrKm3znqOFKoVWo0aO+2/aM015Taa9lsPta
5aIGoEFzLsbGD8AeQ4APQbXFnsDFhF9lvVfTcjH9KBuOJNJ/G8u9dy5qIEEt8QR8
eiLmNh1cWbIXfxaPp6Adros54sH+cZGEvBuakNYk9Gia9bUHYx22EKeBNtfq2lY8
Xg7SMKzJyp8kdLzu4KoEFyZ0gffjbbpGYsAsSzwnHXuRETKnBdQnPy8OKOStjlFI
hJNyuo6BS94wgPR6hDhQmrWUtqANPxaxw6pEcZccx+ZzBk489aKQ14AM4jRfSImm
1jI/2RXcP2ZYrcag+1MDxzDx3E6nkBofwgixtgLGUneLQ0kbwwgRCVScfsHQthUc
kE8uIb2t1TdoMgDPNoo5aj3aNX/4bTXKvu/4jx+d36ak59qGDdznpU4Be1hqqtxh
B3Fkbn2FTvs9/iGAHN2NTdZupVylBlXwoCxxoP6AMAS5ZTfmRUUdiq5AaFVciT02
Gm9RjfrMBnqVUERtwCR/SJt/VVJtVENrOZYBUfySnXlp3sDDAd6ls9yuL7Tk5+Fj
hqiiCOd4QXtsfJlVf8OJCKiMuvDVHIy9+VZkjp4MbAhnEE+mKWkyxqRPDmYdg4IF
q+Yl5iYutstCmyjBvSxSZd89L0lyqMxAG5ZHxBsuEgZ2puJZfRiDTIvQb3mlTpng
+9Gj76vUIDC1FULd1MNk4iv+ZfzLJ5EDpVFXlJw+HdHgHTsFit90Zso545GuQI5v
ipaD1+Xz7VzNDHMPEa6ecsiAhxno3YHOWlG7MEdhlb+50AgwMgkdDI48yk+2N3j1
60PcEboeY/xOqSvzdwuhFWY7mLMj8wymaiJE5TwY0tC4RMxA9z+fZ5weSibjC4e5
yKdWabFbxE/tPcbdxN92HjwiMw//EQgDLxQ9IxsK/VNP4bbpB45x87R3RjCLAz73
1yww9lOB+OmHTiMkBEvQoVjI4MQA+ZtlcuHlzT4zoF3Lpte5tvWyURHm7LSlc/uj
y5IQaokzp+oEKUuqX38eDwxBvsKJmNzvJzZ+ZjPKA8Ss1kDGt9Vubj0q7Rvs4nED
VAuUjn66+flcGlkyvf86DHrfiW7bkoEKNpF31muI3a4HfYYPqgWFm+1MIsxf7Ox2
f5Bg1og1fXoYEjnR80X6Wxr7GouizTzR0OlSoPeHZ/6J6tm+deHwGkmby7AxdqEL
gDcHmVNgKyHPP331Vj65b5PCCCoqsLFLwJsrPkEZChoobP5JF99/J41SuLJfGLgY
GL7dKl07lgjUlpC/PTyBphkZQAjnPuHL8z7bYUlJI0kVXtu/gR8w/jSYBjqrU1hQ
s9Lz+FVBUOT5a+gq0p+sViIiTmxWKRhzANtn0C7SCjpWIikPMqoKwhzXS2v0YXBM
8oKKFhYjctgfT9HpM4UxkypOJZeUkmTOAojwIZW5OA5CKHtcK+4wOdMYbOzbcvsi
Z6+QZXumNsVTJMm6NhBJ8h0SP+Az6SmgpU6TIr4o9+fXpmJTXO0SV8H+b05tt83d
IDPH2tzf608t4zld6uQ+33pQjbaLVX/TxrODY2TLW4TF1D3kE0ouZXb4asSttbDq
rGW7e/J7W06kmMxM7wwD1xSg7aDrDBscxRb2lGyy95Eykx/tJUrKBFBvOpky2Zsv
zBFqymnHaD11YoC4SbjdwMDG79YLQ/EK4n4lx0pR2A5HYOp3cGrsyotcPQndFQ30
i69TrLj0v9c+nxZjek00+Hy9PrAWzw7zm1PGIueoKVYId1zZCrH9Q6A2EjBxqTZn
kgcEMh5wlcApdOFVKLOZr3HXFJ8Q1/5vsWew7qZrweW/S6+MtXKkk8H+M/KBQMVl
7ykw7aj59i70aakddYZlMrUP7AFn3M55K3YwkQ17BA8Rp15Q+PROU4l1gbDk2HXn
qiy1ZRwr0iOSyoGNd367guMmowiEmJJRT9oRDE0gFMmc1rwoCfMKarr3ukLl8WGC
3FKEXNWxkGGppG8qOQ1MuBXVo4sol517JDYX6J/pv3yTdYIewBFvoRZqHTepAgsw
NQjwu7E/yN8LpQzPGd5+mtGDIRWGrZkDd05LXqE0JKLWmy5zn1fJg05wBzlN0Nxd
bPAK6lSGqhcDLEWc9R4RyxhC5EnK9rnmDOLrCY5SKYLojCTk/DHoFw1qr5ykRag0
jsk2eAkic45h2aHMN5ylOLT6WCv9jm7/dT7K8GMnv3KJJhatCo7BVKcZyfXfnbAR
/Tt7hsu8UDnGY8xNh5J3hErjPGm8x1a5UBj0Hl2AyR/dbItoatFPiJqWmB/zUH9b
TWox+8o6FOZ66PC807pb3TRO6LpxBpLLglFHTcrY+eY4s7NgDwPZLwmL6j6O9LfJ
WuyYU8u0mZgIvQr2Gh8a9oBU7kwS5sabUrBoumhYKf1DBrqEluIuT/Cs9UwHWaAi
VO76k9GFPWnezc6SiI8Sgx50wREBeuC8NbWda6p0lzWOHkHHd9XvD+b+hvjF20rB
qLgdWQJcRb6q2tWqxeeyKqBkYrKnXLFbXmCm4WPH9vDw3XC3vLZyombBfUZcPWAV
eSnIy2byo+u5xwesaZotc3wA8w0Lr9nuCXVYxLnuzSIbH30Q7TJL+xyweZamhH0z
bBX0lb4GWOYeAC6WsnQAqL2+jv6xUmJJtqj5rjzJ4Kvnuj9umobCqGzShk3b/+pt
aVGiJ9LMF+vdcqWJTtteis9yMABroiqrDUxsoHHrqCRusPllVOfQiLOdjn6H3tqN
y5kXUdSJ1JAXSyOxPFMvO6V35JhXtDyje2yPWLlwOVmChifm7YxR4JvoMGVkD3bO
Mz5Ojl39TkUfbDf+lWMrtEkFqshjgKvSi9xgi0j/m4I0O8j/eqvDNrfL30bJLNJ9
6SoVewlunlUabwtvrxFGmr3IUkCH1uKZvK4GzSivRkbDxlN8AYfrgqNmwurbAbZX
7srt5BMY6zaOhFkmw/iDunpOTW3XsGMGWzNw2BBYADLis0N1b3QidOhKo2vokXIu
tjJFd7HTbpQTVEm4h6O/3DmqjZi14GEIWkXA2SsJPFD/U7dDwyMjwHvh+u68xQ9y
sDJTFvIWrDHbVnxIK481T0wpr9HnYbPE7DbTAXhkq8cLjkeRDXEZw6u0V/QaSjmH
cdm0nwEbdo3iliD91Iv7te2YhZw3XliLKPGveQbNNPhutxmnGBdVp1OxkLZRzNGm
XuQDk7i51avZ1hBfusUyG19LFaxLRy3kgzPXfTViUUvcDnz29Op4BYXyG21G1qmi
8qXRlKLxG46XpvKXqRzitvy1zeReoqB1ulWN1A7fWg8Gyq9z7qHPIPA076D7MWxb
f3njeYA9/sNd+JCoOulWNgQiIE0eOTiUauR4OXMd1vTWOoGx0FTMDa8fzeXOoele
GxaORlYrjnYzIzOv/EyEFS6kwm7dKmoFcKP1zzNL1kj2YclGRPa92w7t9YETmfJv
7elLHeHg9/+tGRMXNyNN3OV9L7CHYEFuQjmqOQghjnzgd2zNKE41tVygUfjk8QPu
9ZSp+c0Tu4g1yBgeKlZS9S02FH5gSo/G2rJAzM320UT05jkSJha/wsmgdJJPrLyv
esuMRXNa7HA/3EHwuGXHGlP/64jz2f5qDmx3lzaQ5zO4iLQX8NcFYR2DLALt+a0Y
goG83uBP+BwoEp7R1om6K+NEc59wHfh1TxHXWDET/51e2wlIcItDXVzsiVMzMDnX
uPzIxm988kyFHVBANe7x4FJsgR58zZTCDmVyXdq/QBM7RmR4W56iL5O2PPi3T/zY
qg+Hr6VonCn7yUvK3TQbAik7NB/TdbjYiOUo6XwzQOX02HhAj8guYt8c3wvYA3+1
B9oRwpJZ/3z2nZPZsjaQI9P3u05Pbtp1xuNImhEHKC5tvNp+DsKPDv5x8vdYey6T
Bl/m0R04nM9KfiXPznho78vv5JDKwHsmxDWhV9mWXaLBVdDBEypw0uFuM1MXzjHY
OeAXZvJi8XWtPx6RpEf9LbxoKpaSc4kVVYFTGQm22SQt3iZTgqa0CD2yuYSxg4sj
22EfLAzJ6oLREhB4i7d3fvLze1yIzWL1MUdoNZnPpVuFAnQkZ1tnNdBwu5leEVC7
PENpDVV+lorMyuMKWvGn5LCJUQX8Fpg8ClfJk7ZrRhiwZV1NkPkm7bpDQiEgUEta
QtbSzbt2NESdg2P+oJweXbfp3o7x4EhhBQUMLCpZ7200kT+jQtoLgBR/L0NH+LVQ
8L+28AnzSoeNqV2SRb+yJK2RSttQThKC1SjOfsgJc+TWSBNSUtIu7yYBohXzhEv5
h+egZbMHonaZIFz6WO2QmUnKzzsu1qNi2eFDs2/NZcma3XMu8ZrF3iD9hymvb/UN
tsfkENdpd2Y4nCXRJUEIMNysCE8YlNstyZHCK9eFT2eWyHVDIO9UCa5it2gdliKl
PBK2Pc6aCvyZXH43WQSvwQrLqKpQtSkIKlnhAkHgZ1gJf5lKfRf59EHyqSonH78q
02roZfLYK0t9EmfKJZd74DX/TtBppf/OohkntoQcwtd2qFb4qh+7zWTeeL/ZDJxN
kJLRkfJZuPM4ubkXWezL4YsKnp6sBWj9njaoMSqTJULvmcuv/xrElPuHa2t1C28M
XrSPrO5RhIZDV92mw3ZJep/CrKRTVLrG1OH/ebLlh+1x9/aru2aSDGxe/n/SAnSU
sLW4mnyfHvhDaIWXAS38spowELe4MGWZ0FdGjvJoNvIzICu2hJbxaL2J/snbhQ3z
6HA1pCaU5xSnbJ9NAcsBTTJFB18MTHbe93+10u8LwAorzFJrVWtEuC0EwB13qwvF
FScald0nGlTrs5p8TJuIHgozkmbuQ0Z6NJyHkK8MYy7kGWFN9ehQHhb6XOUV0Pun
ZeEIoTmnDYEQTm535sDMO1gLLPXFMx8nFh7hS4VoVP2X26yWuJXRvTphbpwmfc8K
LAbg9kzHI1zNej9RV2uiLx62MffVxlVYcAvBO71c6YIlOZbroxcjTsA928sM9hvI
euYPMImuN9iQnigyxXEnx0wRKDQ/5i41DQx9tbmZ7cJZzC2ALmBEr6xhiNnNh0cn
tKs77FSdxdJQgQvCKpwFj4PNmj6geC/foRZ2nTWjM8tLoFinvF7zVwFjiyBdlY00
Yl9DXY3NANIGWdzBJs6DabYtER8iIaAzI14dNcZMw3ObMMvO9MZuF+Qt2GfkrvDW
ERwDDDigT9C8uVP4ufMWp9L+MKY88LsnOo97hIN9FcgyuXolpQy+8T/u6uqgP/Kg
nU6khoKn0WM8e1IVvqsHjtpYyAwCeapqvc/jf59hLa5d+T6Fr6PgmTfC/UjyGXUC
CjtnXuQy0PRFWddeJwrDi2yolfu2NJXS9MElNw9f1Mi2GtjTJm7ytSl54GbUMTjD
9e0fDI848HmPipS5OIScJOCd4XEOllDnnsO79rio8pytfXJ70g151zvO5sushCxL
keKp+DFqeienICcKe0GcvgvRg9nvqEDuj74fdJVukIAYUdCClItrEPlPdbUimBL7
XH7kMeOJZrHkMtM2khDsfQqNfYn8a1eWr1aOzZxBesnx58d5Xb1ex6ZIdVzR1rmz
bV4iUVPEZgKo/ZX82rSu4kKTTZLPmAK3eVhJ0iWRzTZ/HmQFMXa8Mdm8rHfEVFma
T5tHrTH6EIZJKRdlb2MLMl0Q30cd+fb1aEY27RLV+Xzz+NtJcZzlA8G9z8IoVqSf
EfEOq3I/t580q7Q2PaL/ypA6prh35ucGXjas+1ey3SvCM8CZ3VVwE6FwJmBbv2V2
KRFTUZ4TQhJrv3ibU7gmv4bcSB9F0MMqRLAHcmIwXcbxkAX11799k6hOa7AFEogI
BfsxFlzRKtO4DDv8qgkdtGsrff49m7tc3rM4J7exi1N/n+YTE0WtrKrEPDBsTd7L
ScZHBD4HgwVpnxmL1yJHVI116c47lEh03nmckJNYyABHdwA6NngqhDAHTLPj8ZGG
Ho61wL/rruPIh3iec4NDGLL7JEtAFc1HTZDdvq1DLUMF8bFHKKNS/ecJrxNqkaqC
iWdRLyjfJFkxFCfp1LJJfFNc0/CJmTlQxjHbrJSc/Re/hV+GDk8J/Of5rshAmC7X
rQzlDZyVQL7Nb5E1TBgZTOQAWss2FbwjxDglRXif/9NCcMRJBnur4OldkWUWb8Tx
gGg/Q9rKjUqQUa57ftOmCUwcQq9i/D2gRtk3tSyz6Nq3Menrqk4LgPU4ar0oQ6M/
UF5ccftuci1gDQd3brmiFMjvCJGxa04cJ+BAZT+FwDJsSkaAYD3eCZEb69zkfvH7
+3yy20DdlemMzobhM3sOjJMu/sjhSiOVJOlAGfh+pS3G/w3+CJL7VHmPVSPcOvvj
TUROTedD4+UVLD9ec+ag2nM4Bgs4HkOeRFQxSJ8tJsEaY7XoFpG3G0hKjUyzdYHa
cdeW/jdMu4cMbrbDV82VrZ6aYhLnyAtU0gE9BPqY2T+O0s7etr484cErHPDEcqlX
59v+JOvFDnM70Nbg2r+PjO4zIL7RD9yNDTNNIjZCfvxRasJVB7AlXMqYttVENCgv
WLiSRhwxM40llHiRblNPLZVe931J9Czn5yyI7ldpFmxt+iDAq5sHpnivRZniijwg
cVeC1kzzVxYDdVyetA6DX6ExGH/xyK/hlO3GeBm/rCw1ZRCtSusTN4VcwhhgK9Fh
JEEJ5bjERqDwiTNrw9DtXTf/WaQ6Sh/Og/9kBdtvj0NVFuzZE0yYmyollj4WDVve
Zl413OPPWbH54/uobRZKIDBXJGiZlUVQXQj0yrzRMS0GB2arpnUsMz+2SsJnDY4u
eP3HbB9+fKyOG9FCOat/vqviOTRXDGRLNkeuXSacPPF5XRUgO/uW9US0cIM7RlvT
omSGkFIpzifeZLG3jLvClB8za4e4VTjRyqzTyvZ5SPKQJCPw+zzTP0Vb/vpjR43s
2ewb/3xJJ9Ft0um7yGX1P8bcHOrC8x/91fpp+LGwlwEbkahcjdswSgNsC6cWJdqh
3DKCr9+LqcaDWVAijTDl42jAMutAQquKqAJZmhJO651Vm9jYjK4xr/shCwsA5gGX
o3aA159vRMPcLaHkxQ/bu3Mx7pW1tuoP3+/4ybU2zmIflsRKOqYCCUX2HpKzL3jM
Jsdo0lxuEBz8vEQ86sSnY3VggNivqR/08+eOqa2Xc5aHPNGKvsqXy8DtU8LLSTY1
r4rAzrH9+eR7pVVd5GvIpnRJzBdrItoqsjj4tCx9RWIVxo5Q05I1+VTa+MAtvcIO
Grhto4EA1TjaVgyj5l+QXMHWkvCgdOpL+CeE5lHf54kNuidRllvZUHYlnFZm1AC5
V3N4T4anGNFLbi2Es2qp3CKNAn+lR0NmGWsFWpjUxqLHs6N5Z1DSrxjUUEOrc1uR
6DpNy/h/z1yPhUlbffrWRlwG9eyMlTlBxqwc1pIhGzMjWAkutNf+Uu4+bDIIIgoa
Gwddrw9h+ZkKi1P8KJ4Vxiq06VfrtC6OdshljTNIQ4r3mOTcm0jWKVSjqnpm3jiV
dXiuU+poIqPHGytXF+3Rm8D93nsUNPEh00MUBfp700FwQzljx17js3F3fCFFmEbp
WTRa1zTSsn8ZPQaXhH0iRmzt6sU9ZpwS2MvCdxErAeWoO153X8qVp2dFErSTq79O
mda5x6u5u9xAd0Pu7rt7l/KLzYbIelj885PzGXoSWX3keqemCFMF4KV3e2A2DuKm
Xxsr/37k+0Dq6Ej4nNKfBxRWelgogCo2YK3r9G8aWMnsOM0Bi29tJExgFjRpw2sW
OBhRNEcRy+A4QFpFYIxb58sArxJWmVG+63HilHod+dHOkXpVOrQRGyDYeroL8Aal
mBFEgwIv1xw6/sfiRvW/P5aLOE++OQjPzLAyLxW0AQDIWBuM3zva0xK6r21Rt/sZ
NpOTQIi7AGne6853fm0BZ/o6JftdV0Gz56uQnVCLdaxIFcWc/g+xcgVFmeMbw/Xc
98psqVl8aGIdSK8HQTOXjjrJIXVOsIcj2r/n5AnJgY1gBQ7QmUflqM6ZdvQTxeu0
xjGRl430OJV8HrmOJbi40jlhuQlTWevqNu9cGbGq8GS2nm9wOoHmVZN5lAC4dIT8
eLLz9F2xgqXu4q3ey+nMud/OIoNXBlrvqu8TmUBByRgbCmnN0VAs4Gg/dd0y0aW6
c67jnLhVXW6SUo2dk/eQyFzyVM84sQtpm24yaqI4RNT1KjFsO3onlStD4RmzZd0C
qXINa7KGajzdTCMdIrqm4W4EkOqi6wBiVzpVcGMvlYGcW4REfdxCELL4Fz4GyArk
TFYuq4uVHjd79UzlEhg7bzGSn1dUZgZURjHwwKQtVRHyXi9noGD1m7+jHFZpmE9V
cI7cUqNHEueu2tGOGq2L+NjrpIM8VLBRBYOArCaWqRiYfCu2JcYFs+CmUPKoeV3Y
C67wdVOarQdE2dO/moK2xLNXJVxIgfEuCfuhYSXN6KViIGDLnuop+iWIe3TCW/Op
d0i6xyCD2c4n+uP+fLC9DXinTDAJefihqEgntiweUI6XCIeBf9M00sWefXw6uAcN
I6SSvPf4aSSqhf2De7t4M29QLw3KaB/cNO/RaS0o+4PYEw7DH8wK9aM79RKHdoad
dsN363ekt8tgF2nSkwYorb7oRJNyTLNKrXnofREvtlrsAxd3dO02l7iLGbkAJDEs
cBhkyevP2KdokMjXv3sPdceYXNKbzCBbS6bGOD6Gzo92s9GrJd7A7TmSVHBMiWwH
wCL3PmdWU4M27vFuCmvDX5WFoME28EQhIr6k1OY0uL5PrcLEXdzLxl/zyLJQaOIM
7cprK5nWcaV4C/e/7qXyAJNXi44/ikwu7LdjDnR2dwZ5RrnDMrOx6Pa1a0FrUEbP
FTOseBzvhve7awyz+DKzq4JAkJHwaDGRqsbdQQ7UL0t/DV/0eLqyoCJT/eZNsOiR
wvp+1erVsVLKwZHuigyJKRIJH0RiV1tZVNfOQKSGSMsDcUwnhMpcAJXjH20hEm9H
rkZyv2Nx3T9ZTPVAhIQEaDjJFM2Dv5KVvVgJXrbrOTex78zkNUDoeLRYgtLli9GY
G3WIOhAbA6kc4WptRpnaz4n4g7fnuRpDWEwmXl9uUAlCYr+w3wHj5wFD7dBJZJHZ
mXxIuRO3yScYolJ3wam2WyDGtqo/y2k9RFLNaoGqhN8uWMeYQlzuFVXR5VK1+Ap7
4Rndiq8/Bp+/3UfybWomXVnUfEn+bWPlsEcksgkOjX7Idjp58erz5yXathVtvsqq
fLWtMzzScbu94VkxBxCOAdScFfWOnZGY7OVCcy81Ixux4A9070yfluRdj6oIOe/x
xluePiDyBw4oziIdsLcS9bmQRoSsuiBQOg4ySx5GaDhmY3fsQQNSYeXOc4pYbOFa
W2nUs6q9EC/r2je+RTnOFMFeuPIwSYUqAOeOoaSYK9KZi+iPbjlCLPr4WPAtFYk2
pas9YG9Oas79U3obsLXGPBfSLYKLipYejkqYg04/xWQ3eGvNZDduyvyGoHJHYATm
T58hLxu3fUwAT7qzOk+warypfLOixW6HMYkRbVL+d1J5HwyiKB+FPlWw4zZEXzbv
RuQAmkTOklEHRuYht6XtryqqqB3UbhI3kYv6rNlcMXFAT5ceEDH3skxXvgZOacxc
3pM1f1XQQQqIVXfThA4pio758HWX+6Kv32sWCoiBjWsVyVsRly/pFB5EKJSN3II2
FAktCCHDRxA2iNEQyjspVJcsmsLUNdqSZnkD2IDih+WftPO7b58N9XlPq5YxWI+q
GjGArujdEGrFTtnWq9LKj7G5guJ7blPbuTuUuIoBlWFQF87ZDuOZe4dqsu1WC+3K
BjyjDD5AVp7eCeqYGHZWB8xwLazNbJlYpinai23qMqosusLt1wvF6zlmzMAjDtYE
TANzzxOjGLdh3BffQJnkznB4RvGnp6SO3+huwW6jz1E4xf6yffI/Axc+sA5ZdvXE
Ra5k26AXu1vy+CvwBrvbqn0x50MCz108p1s3Te/cGo7+Zgduvs6+oVFdZLAFy5nF
CC5OR020+ZbVMDGw/EV/U0M3utsAn1FxH+LHgdzteP22Yq580eY5Z0Qfnl/3E54t
0z4sTdU5PifTQ6IRi4GDmUDWerWjzw+hhppV725X033YuOs1bV8ld44tbME1k5jB
EgPjzz9nNactUkb5yjHr/qV5fzZYMTuU2hdDUcjTdl1X33eG9rmJJDTBgkHHDil5
yDMQr8XnLPzgy350kDXSxoH8462ju+0Hz5lRqsyBHTFLkDf0Bf9gCveR4O2rnMaV
rdXkZKf/ZycVHc29YYfFVZ6wSeyeAt1zEJxN9avaesN4CLALEkhGyI0Zm5mUGI17
vgL6MesjHft6I2ESJIUHiDDlNAqi2yeNNgrM3Pq63ciECShra4wOiEvA8XPQrdFs
lx0e5BXxRg14D7TIpzGYoxkk/vFgZ1ZVZ2/2Ca+CikQS6ccnMx9ASyZMVBf58PdH
9TpdiHNTp4P6bPi7HkxrrUSSBTf4VQpK68kYVwmRzRurlmqevwTEEQemR2c0AXBF
akjIWzCHiFDbT6nKTgwqkp4Y82INwbRUp/uShLbcp+vlKaF9Jpf8XEsvFWQXosQW
qT8uMvtJkUP+cIi1UPFvZ7XWKsvwIkfTnwA6V6e9g12QSlu+pyiyRHiqDv0gX+ky
aIVBRJx7lFySVY9xATVMvvziFBQu06itHNgcuK/HpppbVJaGWndRzE3/Qgvm1rIc
DgGEVZ2m3+n4NAaM101sISCxIOuWSiZa5VHXEk6eQg/Zsd3TFH03kj/ehh39Ds+i
4Ic827uPRDynetfZNhmRmaKGLwN6FmkQOb1klZRuJjsZzr65FZgDLb9m7JpRhfHR
uZ9WN2OUCutnCx1DqtO/kfDb/DIZcYiAVffLB8SShDyibZbgrQxE3x9g6dXryCbL
qt7TbYfuHenp5CbH3uMn9vjwFW3y/dkZKAX+au3lCg/JtJtslbWsUaqjMDOfTxtY
IsgJnGpTCJyU7yvFOSdzYK4zNqKa7vOy3tyjgc0sYbRtaOw/Qju+y7LgvnqoUntf
1MOUU1GJTqW7eI8d4EAA0IX/fA69HghIEpIzslDct5oa27lKNqswogg14BAq1nSm
NLjnyUV0Y94OivmoRbKNKgnDfubsdSGEr4SrdZYhmRmeQSgBlh/P1VM07FHMM/Ki
AZLZ763m8Gwu8DF1v0RHT7FmKHyc9/gi2YxvaS63IaRwKmYV92kpEydLEyWv5ddw
yFTXN2TYyjjLkBHdB6saAz4HvhQdReq9p1R1NYgI8YSwTn7IE6ddsSs9dpTd7dqb
4ofeiz1pnKiOjLGWdkzZ07DuOS/sk5fkCUTBuH/Jct1DsXar7IyV0FgDxVk1OYk6
wPuz2BiiPbKnq7IjNa0EqEmZUD1zTM1yNVD3m7k35DMKC9FTi76opStkbTF1KAx6
tLI08Zt3Ojs7I5phPx8jfxGwdRjI3uXw7OGdqscPX5RUVErMWsaMcZWSwE7u6YeD
87+di6P4vN89JyQa4ibjozuqAYnrVcR5LwIVrMVaoHI72K+ChGlOFDtqGxFMn+YN
3+gAcw/B8EmCLLrjIzzrrpYiNUy1eQ8Sgp1aDWxqZoM4Kloc/qtZGalhRlkWS1Lc
j/cgjpx0fy0pgsNmbpyhVSSutQhCPGluV1SLH3Ya9HnQOqbJGvPE89bG3dlyoprd
8Gm1CBu2U5t3BuJEIGqE7Yy/doW4k+Pf0sj0J2zOj8WRVLPt+rVQu4ZoV9VxyF5A
zhGjBV3lL9fxEpyEiDHxNyeFFfdhFHwaaazlYMjzHIkKu7fYYzZksTn1Hziajh7q
c46nBV78nOBU9JVd1I9XXXvl4sBo+hi8QYPbOu+QgtVDU8ll0iBnbE7Q7YELtPg8
ljIlHoGDWWEEFEBPph7iRDjggtLugbgoXLoiBxdtP6NuE8XmnQZuVLWx0zof2nqW
aEpfsLi12RKKcSMb9s1O/Rtt5r9oFAYgZcgoW8j2vQMciDbuSGoYuW53WOv1a8F0
kaxUKkoaSLZtr5Ohs2Pn/0RokIbfT7dKnooiOHqlMSQqRRnZirODDeh0zkE3aiQx
oOK6lrVZISolIPPGnl+BZ5TLwHrpBcpq/t96g5DvWop6pVwFIg3jCDuKvdPBeNQg
XkUlt+/OfIK2eEP8JyBrbABQAVKOYy80PqF1RYISLzHufcjstCIzqOyF9MTqtWFr
REfm/VWzyPiyX+fY9S9drWGjouSrPB33eFVEKhTcPmEjc/6mzbzxVuGb/CpalYi5
R6QsCukprz55o1A4vYgZuBXv8beXuMHPBQY3PMJqToez6CJfd9nudQO8tCzGXe/p
u6peDC5leW90NNz7F3QcvYxrix6sMZBz9ltZ+cgH1mq9CavfZ69m1oND6k32XSoD
2HYkNg5RLu9JaT18n7qg6psJB6RQkkOs3sGztbE0lX6iVXuX/TEr/4CgzDJg7OSH
+d7OskUqNBftbNAbbtE10kWxRRQzPcO+kLZSQD9w/DUb/JQN79/XVfoaZE2l5FHV
WPZSl2mQMBjBIj9isg1i45MmvYX7FBoPfVXn2ACo4qQUDwxAiZXlgaPypmBWffKZ
0QHssOKBAQ5UYZ4mHWjoJlDlpkfIQQih9iPCvCaG5Xoh+aX4whVDjyiDdvR42YiV
FFxGNpGrKUfZCvl0LoTHoxGgn5oYuJdOl2JmuxsRyrLKGf4tVoHCdm9Nlqo+XMIf
25sqRAsi0wSLtM6ZNOSu0cGPW0wwNS/FFViUjpFLi/eSWJD0c2WEszbQpS5XH5+5
fgeauiNTUQQ5HviMMzbcb/ueB8ZF5N6ypwCy9ZUG41bCA7XJrL9UqH+5OYw/qpnU
Hox0Nb5zsHmFwXtZE2A4ZatDRJTQWz20y1U5+MZEmfbnirtjELmzIz07gS7HyTtC
ELG1aqC+IELsDV/TplUPGc5+9kBrvycRHOmRn4vPZzBHZCuEY7I8j2KxTI+MYiRz
343P0TguIg11DXJQAfaHlgXYY/zSyFmPuOJB7jymUfkNfsh62hBsVKe45jrlHgpS
v/RmPxf2lQ/ftmTuzFHJaa1udxUDLonWcARr05VaJSp6CW82hWPWhWT7A3JTZKbC
W93WBWrngAHucpf+sFjP2Vz8h3UancwsGkAT6tNhqEeLp7jpGIvqaKszKvWoPbSB
ntl8QNUC7xAIGcdOH+P2nKXJb+Lkv3y3iUAUraDVul94WnYvFynZ332q7D9XJUFn
GCQPps6i+w/aGBWf7nAk6ggjmCoyhxUTE+eksspAtaHywYNsYzFQ1miAJwa5HLnb
D1D2Tkna1DOOAYmahvDdgekKhRCk1xnSFjBv0wTZ0UNXaglQG21hcKaauEedYeY1
1XHmO+G6bd80un8ZaLE3FqMf40wJrH5GWrtBuHecIczWiNSL+OhdDRKX4WcFeWfm
TVOsKnU4cXUlaRMFvfYxZlTs/5/spXbNrcaunzt75/egtALJOZOo1H/14PCNDffx
14miI1C53FhrO8MkBNwBNgR++xHZtJgZXkPMN0tlciwAn53NBhzbbN5xuVLUir9f
i6tIqmqmuu6cDO4CYU8cZPCqSUPqGKbaB3amxg9T8Rt38EYXGMuBwguPmCXxPbtf
zqOKuCnSx9YX5Pgh5imZwLPiL0//gnIjmiTAL6dCultmdBvpB55Ri+vbFvHX16mS
u9nOClXPEHdSFXWWfV0AQcrGMwaUVDtZG9Zmv5SjbXqH/wFD1nXIKvfUVI/NTm70
KlCQvmn1CSkAmtrlldKnz67drSlBGU6x85tNyzt57dHLKDEgaU7E3IkuF1EzklkS
VPEtPXh7dzxe8yQZBcyoQEmzW+Qyu3bHye7/g1I6djr4QsYk9GoLCVcMkqgdCa1C
VvuUn23faBVRkfhmSAw5m1M93kMsHp6eTW6qL2nmYMe+3O1R8pJyahyKtMldpAUJ
Ow6JtedMlWDg1LE5MCQ/rOvalUlqzRAiWJsnMzxcArkGPZufT6PJf5/QNG8JKWj3
jahFTxkoBLfRVE/Wx47nmAHCQfO1OfNikp//oQywHS89uB00t18GuMgXNObdOsju
nw5XQ2Zhr6kZmwFU9Tlo9ednMR2AhoJy8PdZpKqxkOArd1LO1SGViKew65KtcnUk
HkKd4PoI1a4TJrjJ4SBXl3IXipDgVGqIL6TPOjWz9f4Szjx93GXyAlxFdzIli9ON
e3gqS8MbpzSGnCnOkOJNJWfP3G9hsq9dtvqbyKKRKHs=
`pragma protect end_protected
