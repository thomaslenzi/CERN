// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cG9W0z65n1GglqNTBI6sVlly7l/XlhFHERunhK75hIC1/ncRzqkmhQXbouyaWPWA
4AAYzhX/7rpdaiDiRYDEmSj30NgnPJFBeM07MtiXgw0AR4KqmzW1SIHM84tTbSAd
b3BSMyvPoI3dVX+sAcI/KKkz/Vx6Zs7bRTT941zJbPE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18784)
9TNDzSqi7GEXAOxHTgj7DnByIA8k5cxYFVg6lsSp4DJoEV4r+/S7S1RfVACtUWT/
cRrngcaLJ5vC4g5CM2gBg7YUXSIcfABx4S92Va0/Dx5PP3uNwDrM47ER319c0kt3
py4WJ+Xylm/z5yMa76Zt4fbOFoE7PDHrN5CQVJtYMWSXxKV0O2eyJx0PycsweD9l
Fy2GLcpSaDsSdX32W/8TWB4rfhRFQ9KG2L6GGj8SAtm/FJySqq2hjP23GXUzIIzT
tNnQwUaDVenkTM8RTLqqMYLmdHHE3cEo8jiiv6SiZVeMEDFTLxuWoN9EDz8xiGpg
VwhPFlHKgA02PsDABVGaZpVx+Zu2mCTKy3wxYY3XoHje+4nGh5lhzPJCnlUiuEYO
6w/MFhYj+AkGX5cPOmEM4soTHIQDu2WpmHs4IXI0L/yjsrvOd8w2Hcobea3jPYj5
RQ2MMMjiWL0WV6qwZfFR/SaJXi9ynFdQfinPwH3eZ7uL/A8xPEjpMcu02C1nRe+r
o1gNvZl/XTaUVlYDbibjogrIHk5RBnZpXvDmVrGQZ7IJYQ+TF+m2OhSsBcGrBWjq
aYNJkXpGWp7m0qt7d+I06EGLduDq0Eo8bkivmoqjxXN+VeR1XXmXGSCdINra4LnP
gk8iZSc+wCIkgsrhrL3jb7c1ZDD1LP0jQm9mNmIXFMCbR/tJBe997ojzNQKLwCKO
5spB7cMEuM40LpcBXi8NeVYQQrecccLJWZt+CcDomvxZ+IlY8uFD6ZlRtzO4Ut+2
X8P/1MCQESHBWdLmGzEa7Gpy5sYTCe28uHx0YPecx6XqgFJwtlnwdvgIN8ChoEo/
x1nu6W8ejR3haiB9xhAOMqQV/BckJ1w7SzYaV1YQX21dm28qzZzOZxkXToxWpnJF
HnRVT98OJxHuFHqJfQ3/FoDR/bKtVa0KxmyY2hUGJx2uD58tUZxfPT/bK9YxhzPW
eFqV5M5rSH+fi6b20k3XKmqsZDEB+lWyhcZF1NvdqEP2b13Y0e4Qfp+qpdd8qPU+
rAz37zDUK+rnI/Dh0P8FHfu+SmD0eEk9qHebhc5T+kJd40PZk3WfvZrZB/SWYfVG
QAwMi7ByQEy3JPmVVKdWCfsItA19Y1XHXxhASnabwSjsQrvB/TOslyf66gNAHY4/
FezIh6+YhZdqZFOV+LUqAulRzScMm6Db7K47to6zXU1YnUN049wG9i2p4/Xc/vX0
Zy1QAgN4Iu+y08INkxKB+l2Pvt4YDomkq+g9WzmWJ6ypeTqrbCWWcEU07gOi78Te
RJ2NEg02lnGCzvh6HaZ9K09d4f32bZf9IsVQTUY9xgiZqjTIz0PPmtW1MHMiT14U
AB1JLcX3en0AZ7cWLhbVZRrlrMmUjECY4T/QSXw83y/Q1vZEdNzDxNaDvXdMJw6V
c1alO/Cgl5uYvxdw1ar5Z9izLBEsLo2MG39c81Lpjq9D0TnfzCEDiTY38lY0HJrA
SkxuAs+48Rdr2F/4gbd8R3FSc/pS+AgWottuATP42n1iS21thWjip4c7scbS8wG/
A9w5vyzQsXLeyX+kxGbwriIhiqNrLy9MLlNWZ2oDx7ODnfNzohIgQCepgIqOElYu
DRnVjiSppdRRP97TjWB3dHhcBqtxCbJ18zWvBirnfOCd7cHotIKsKF/H4UOHKy+l
FvcooARQ7vH+FgcUGRfoT6hsZGRX/PMNt3znr141ISdclQyFvTz1socSET2mbkXT
nW6aPUiGJKOADS+wy17TDdcI1BXPVk+U9TYWh5ZoIP3iNL3APIEIzNDZvJOS6Uvg
w4vzycGKUqSuBpKIO7wpI7nbFoJhYsNC69TcBG8cufpKu/kfhS0Pjk3eZ/SByPY1
mlxw1fuWBZ1k+WnenTD/DILY4kN8Eoy+DxJMLFRueNic3DBigwRE/e8RgClZ4v11
kMKdxQzFpFZ+e0oW0NrW7QgTl0vgO04uubu7M7/h3GVNR4uOz3pmViZXc3u2cfYI
RpgUXGkbXYue0gC+KfLjN9gW3zikkdkSp8Oq/Ief606soDVhJ1GF6WPEIF5QjokZ
siU6yZZGvVCuC7Dd4zg7VhSZI2RgVhHiYKKddadAYQbQQx9btPOvRyA4xFVLICoL
LFTn2NXQasvz7VFkktB2y7H/dxrj4skHonJr7JaTBagRQFQ7XE5pC3IgJxQM50oR
3739NYjWnJG2dJMGFgkiXQXz7ZNXuy+wXMGG6dd0ACLKwxO7Rvciee+3zZJ4zTgx
i3wAx2pXq8ReqgYCFHasuSWnK8M5Yn8MS6S8/nsp4uBDlDdPa50xOFNm8kRTE1E4
MD4FTLLoQPYz+DKIB/Hwrwnvqi4wjvY0bN/h8WlDuPVu/3OFbHIMQIEKfw/LM4lR
nvGBXGYyKOl7jFuvcpu0P7MAi05q4vrGaRnnAg8posZlmNMkc9ix60hEYcsZrdtX
Xd6ByuQnktK97VttklyW2+R/CtvIJvTe+75UaKiR5qRawsCyb6MjIk9GpgqH3XMR
VjOwSNPSYGTzNfQAynbYJARunhkdYDxb42hRYUcXS7HnVs7XTonBucGsyS0PSeFs
ALilODQjLUxiz26GFDfvL8fPH8fC8kRE3hj9zO3AuhruJ4FVf/XQt8G0It69WyHW
GNaWy9h8nBnSoQQVF4/K1B5yqf4D7gwgHH1/PyOxCW+dtqojvvIK0KQ5et/Tl5Lh
hEA+9gsf40K6TRfFVZZ33c8PNJr1+gX+Q6GDlvDfRdVxnM/ryv7mr4ldbF8dIaVF
1Oix3RxrAfRtZ9VqIDWzRpLNmDE3vH729kFMWkQAPQ0utV7+e+01ifmUcZsyGIpA
WuTwRcMyyD7XMSp7mPI4sfdgtMTRKVgxez2PtYuyDeSKMHUXyrEscBLh93D5UpqC
RBFm+nhekazCA+WOYGPN9sM7GN3ezVh7COIQBT0HK5df3eB28Bk/5MOGreoHKqZr
u6yqDng3wREONITNCu2lrulZklozTHDRMol3Zo5NfiFXdrTqmTkl899ErnmY2REB
M8JR36aQw/qOlhxMqj+eCw8t7T4CaqJ5uLsX5Dvn1GOVq6r4vztDSreeT/BRx1YN
LjAvgcTLT9D7uL4xnA4PaF+NUFvUtC0lT+XjJ6diJ8KP03BQelc4ssO1Eu9rDmnF
xPBLcyLSDMgUJ56ZUVaOlO+26aPA8h0Rwx1wfcLhyu0VISgZwgit3zPloylphPAJ
rGKXHl4vwwgzGeXB2FJd8OQ+NL0JiP0VcXgCUyiTCvzOr6iKLZfXFlpanQt/2e/r
EHlyut9SlZzjeMbsbeLIWPH5YMqw1KsBG0sLKmVh34jIu7QF3AH0eWFvo7ZkcB6L
HXezP6gsjHCXwnYLkplZRAXn8xwY7GpR4Myu0ES/Nbg15pRCyTri35KRaTgB2m99
RNQceuzDp35pBH0l/gKAzAIVg5TxkILj1UyOaxkI6awisYlailwxEYlQs+jz9PcY
m2+/G4g7bllAPRW/ZsUpEGM6cLuBnUcYgBaScWmAyASuG+ZdFMkY0WbfVSsSxf+f
Tp+Thf6CjsvO0CwFTm7DE0bcpjG4eFeRO7i6y/EFQmHF0P1AVZ+jAKc/9UyFnwLH
QmCU54WQdrhxWkU9dhfRJRCpAU/hy+P9GdFMqUVbEkA0HNXrP6goKTcLvxOSAQ/p
CS3+j6+hMXJmFZ4QhD/35irge60oaFpKp2lywallEsh3UJBnlb5Xve9cW002AwaP
ebmm8cNStquZUYkZ+ETxLtF2wDzWA7Xq7Plv8nq7gNGquETtYKKTNxVFbr4eJ7lc
XM3fxdlTxh3JT6Zy16tXDxx2wAVKvx1WN7yhAgIG30lYQbkCK45dYKldKSvKeePa
fz+3p8QrLacZpTLRLpUfo9M3LOBpeUFmsCa97jUj8TTZ4/PYZvTl3TGgOw0OGjk8
irTVg894PKLPF4R0+5LsOlaoxKAFrCRqyP2frxF9EZjMKuBt/S42iA7xoHZyMFtf
1QGkKtwpQLCZrC+YadH7lFrdPgEKnLyzmuBdxPD2oeY4H7s3yfb3FH9ZQT29oTKX
XCcGcy4h0W+CfCJYla3ANSPcvYnGIEZYSnvG3ASfrwebKjDzLnJHWJnGn+u7HIIn
UjSwyrnCnbWOawfBG/A980nn5zcrj5tpagRfAfPBwfpaKXesRerr7nLX4NsUjBia
gjz98q5fFRtOxMVuRoJ7TgGdNPx+/yiLFc0HOZnMGjJcFweDGfMckwMmft03jtvs
nao7RawhrZ4WNr/VohmMF0EP9bUx8NL1uz1+DIGxQg82EMBtZykW1u0e420/sl8a
gsM7hHYcCuDsCDBDOMHKlteCXAIfnKO87+YFQDCgQwzbgPaEPXGANn4FB3jitfkw
MGJim8PV8qEhLJcIDoNW0laXxOZXxtQHTs7uLAYgdhd7c+8yTZl9taxn2xS/Uu07
/LfSraavi6p/Ad7GwdUZE3z0246eIWFiTX7HfTIMX8E+Egkoo9FB266BCTigl1hV
B2VnKjhB5qB2naDaO/AiuZ8SXWVKfn58ur39vDLQ3MD7YB2BanRPCpwfQhBjYOkH
+ucc6nYDLtROsskXs3+aCs9oiB10F6Kp8OeU93+aquszvIu4pIttY8J1/9t9K6IS
QSe5bJ4HpxhtOuwu3Scx0JcxfSLQGuWuGvPFUEUgJapmhNNouwqBcYUPkWjUEMut
Irt5DE+lIZpOQd9VRotiaZLdtEP5TZOpkbC9dkvgAUe8pxa/uXgxqGVkfZMj4Bsj
mDPUuixCf/neSNSKjeBVi/MUIFgjZc+apbvTVI8GYYUgxDADiIjHPZxX+wHgDB0+
bEpaUuNEaWCLkJd0WrLWAHBdX8hVVMdmRhVFWMi6eAMlsi8uCpefsPX1opkJXYui
ZvWTvPlzDno5yXLj/iy/RObk26miaeSE5KoxHOn2p9XcB9PX0RrnYHtt8JtDzJ7+
mXqZQ+kkVTe+h4DCxOG2OEblMr7d4Mk/5kV2HbPu2RntHoor39vubR1DymqfICK8
Qr3BD6ZkmDed38SpLmb7yVedxboYnEOkav01b1cYtggYGqvRtDJEdQ6I0GmiCJY5
FL6iWGDYj6gKIpvLRROgXlZKURBma/XV01p1d6HgqvCAHwbcywrtGaIOqOqrgv6e
reIHYBcNJVfou03tIZJUIe4kSaDVFw0gHI8PAYzTn5FOsNy93t4BYG31jruLzb9V
tBxYB4DFZieECBPVozDyMZelTEkVwqnxTo8gotjqC1jkqmR35Wh+3E0IhpMaDUyg
nx7KheRxRsyPdD4qwjwOJcmjfaFfws2R40CqslVm1Idu5lznx4kra40ggQTd+KxI
qTgLN3qNsHGlZ8zQIEsKE9vs/EFLW8UnhxEifYXh5sbZiBl8SnruHVOfWzTOhHpK
tgurfGRX8hDWZ3EwBBBorczfNDn2wSlHAeTbdYnyOcL1GLoaCr+c8w7FsycXICkr
nmQWHwhyLj7FK0znLTRyKKhMx46SS6h+pbiOomjEtVwab8Hr3Ji87EascnLisNsx
oMAH+b/J63e37eWNoQ43HTfMZNIq5yN+KQfczlIsGl/tt2X1MOSv9H1VJtsMWG3x
Qzw1L/eG/0bloSePELwv6og3fkAMUq0/Tz22Nu6t7O4SIlqCsrg8+WXVd62tcknG
JlWANFdlxIknypUrU+9VB+GgrdVuuxzIOtyc7F7CgJBi2iv1NYbWexTR3sZkC1Rt
R3A5k4eX2ujkpyah87MV+IPzylllHicZzLy7p4BsjHVxWPXVn4Oenss2AqA3tmZD
BitgY4JAqy/8pH0yIhUiGN6XW8H+R+Rr8i6bS73YSXQ8s+oUMvDpgnEnhc+fJzC9
R0j9vJnRIrd575qHvbdVg7nNLvIJ0XuwD7hrPwBU2yntwP/mHREPnDJXIhTbKliU
vGCJknTql1v/dFFHb/+iztgRs/Q/tET/oE8581l1l794FGqBVZJEJSN4KB4ROZK6
nPj0fvS1T/6RkXJhqqa5Nyny1FkTgcZ2YSjirvN2KNHti6Q+HqkISlFDO2q3YBQp
3/d+uEUxcn7o9mP04A/XZw3GzFqlS1hLkIwmIT76peGcPUJyJn4c84oUAWalaA6a
NBza5FviHR0RX0p6n/p5jXVUXGdYx67qqqHqijhLahfa1qxDYcOreEjzB/oP6mxv
/ajSZMdusmars5F62+6Q0Oc5NRU4aTQY6tH2MPF/LPr3zklOZOP7btm0LbIn03Vx
tBdxiejBshu7KIxFQkL0wsZVnXoujOtMlYUhDAMkNfoAkby+X9k5MnBUWpxE0LfW
YSIrAwhAnvN/E7SObrsX+ju2j+xWQrU0x/mzcJ2fssAwJB8PN3Fb2AHIuyuzEbLi
UoDNS5B3wNcGoawFO4RSpSKVcCvoCm5lhGcFNdqPXAqWluTm8xsgzL/uhu7V+Fhd
5Xf8BPMNpv3A8a6U0RPKG97f7l2XMAMCHgIwX7sr2+QkUr2wGONXUCeIfv0/QkRT
j5umSfMU6TwAbzInGa33CpkGNHtEilxEmkqLSWZLyUjLqMcJSNyb3POC4I77cV3d
DZRw3zdKd88s+CE4uXo0fUj9/dpF+ktAgKkNhs1M/gvPoT1bk3ey4lALRrzKMoPm
580tPlkKcfpcm9Hlx3KT2Ikt+4emzZYuxEYoRWCMCmCx0z30zk3xeG+bKdQWsHZK
kCkzSn2EPaBP7khwUM+t5paNMAxZ0L248Mp/SW3z3tRHXDuUEvv7Y/hlCz6HbcKy
afKjpDpuVPoVbMDYjGjwlvl/UMS+HL4w3Qt043IPwI8bbYLH8QdOY6pxRclZsbn/
qm+rgODj3jqmc2cSMdauNYhHG60CYZPoGj3XbVLnQXpy9u1thX2MrDsT4qWj8U/d
YHtVU2MAJj97cWjLzHFzxlMbYuHbnaqo1wfUWY5Tsp+Y12FYJk553dCQto5U+V0x
NEsBjQ0hZnuQhSFolzTAmQKWEC7V/RKZNxWKTf5ifNIU0jfw+3DrnOQjTSc5PzHZ
PA+R4woOlpgClcvcW5B/lFz1TAc/joIQjMNQwN2DpKE+7MFNKEqPNC1EXPOp0yoS
nqvZaXx9VEmTYkUex2pMmqsnDTkWea4e6ObJxYv6AGNKqGOcPKofjKeZ/+THUzLd
Wp5+OsSkcqoNDF9s5l4oKuGNfbWhaISQ23sHMYnHZTkXbJTaiCMqBLNcL9y1SNjh
iGywhwGIT1O8tP7YhGuPh6bQm6vQ2TqpRm1cq7HlEbTDlIfZlv5NVd8DY3xl8SZ1
4NSPXlL2j2i3gzis+aPWQaTEONTZA/J0uF3uIw1+cGkK2552H+iQRpuOLRvz5RZ+
DKdpE7txVgvGahjOaRIBEKzXtf4P4iJif6t8vr1NqWrQCMtjNpxQZS1mj2xKkVQu
FbnOyYtQU9QzjSmM0MgzgkkKyN6xchIcqXLvp4JDEPfdqmdLH/4bwVDU5nzem3W+
cdmmp4zk7zZdhsk3x0ldbe25AQAdQjizEF/OtoqX0yK9R+HevIKU36TtFnlw0KVG
XKctfM9JAPubPr8bG790BN3Aqm/y+PO0mptdco3BVMAPz8/6eq2kKuKbFHrtbRHQ
q5WtXvDVhalsotK88pzh5CpeBpqgybFBjjwrnLetq0vGBgUGDeEOBptGAQtI5dF5
WVi5udgb2o+PPvAO8GG9BZhhhqo45km5N1rVl+AHVuKeMnkC1/DzNfWsVKhhvKmY
jx5/BBlY0EVEd4K7NrjSAPKb48s29yh9+6tg43ndDpe9a82db6mbf1IRFRUzEwZr
bm8h6S67AMbsWqMUyVt0w0OOwV6g3Hk3QX/Xfq8mrUaar0jvY5o57IvNjTrqd/+Q
lr1y23sV/YCxLU1pPZzFGhiF/c+RKrNUb1rH3xyqDEG3fNXntuVhiKdA90WOTmLE
so7vlIjdgBDxNf8YpFXWZeU0G/rlB7/xKQt+rC2ptdrAb5JRdyHJTHaoJnEpm2EW
OKM0C+p/bfNEIpKlqO+pZmETrCvwgV4Jw2Q7ojh/OkY9BZMW2FHwxgJvA2Fxk5ue
xZ8UWl8oUa/ksdMOW3qGxeWmmEswd1UVA95HANHCMYdwCaQs/b231CqTKfAcDg7P
wwPFsKx0/iZRLr4JbT20SOqWnKxQg6C5Q/zY97Fz6jV7f30hykk1CuHhmNS7y3EW
o5TYKKRuDnezKog7EIUBlHS9dC5+dvA5p8aLMvMZImqk3jRV0qW1okqUkxwd5nsU
gGOO9BtMU0srF5J/cBV73VP8o1HYreOa+yqdeFWVUAW0F42IQ0acGhuMYIfMe1Yd
x266f68gXErm5KFOFzOaLCaYqNbTYhJ2NVsFZeRoEF0Lxm9tSmpSHFZsfvJpJ/L/
jtbC93kXziKza6aDOxLiDw+jksgtpA8NHjIwl7EtIz//G9viEJ3YR0gaIgUVx8V/
dbdHtljDXZV0oimLN7RQP/DwY79g6eNtwI6Zqk0EalxYwneUoQs3F5/hCAdOMHl/
1BsCjnxLBa6iCPvY7hHfZr9bOW6RFS6iyqDlvrLx0h+8R+DxpdgXlm9InKCLHIWj
58SOrWLiYkS8BQ7I0IRRKW+e6JeuUPWVlHzJWmT+QfxFDlL0G4YRFqVpvps1EYf0
w8B7UbTkv50/lVIJH6bxEOo6+BQLPsN7gPdCNQK9ylY4K1xjJNiMzWFKbm5x7dg2
XiwpPCpSi3Azp0t3f0cP5NoEi+40yx/+m1Mis9qlw3rKV8Ac4pPxr8/Oyidlk9Pd
g1WaRju2fxgN/uV3aOSiLwsauVKRDbuydgGnWOEeQHC+cfw7DM85nsje9ikWYVp/
+N8MBFYMvrbvf48nfaXVCSUCndou7ZLjSiXnZTMU1p3qU2RThCf9luaYDVViSw2+
INlJz30ldNJzA7ynad3W/nt1EVEjeg2ihHpoycxsjHyteON3zeD8KSlfJpbbl5Gm
4BgvDsIIq6XF49Hwj/rUxDyoWL5OWwUYbm5vV+3EVQm/wK+gjkeryPpT9fUBOlyU
RzuOYMr7YI9C0Io8ASSv46lB59s3qhTqvhchXtjAOJjeWT2p0XZXOLnY+EbozquT
k1HxAL2AXxkX3tGQFY5HLed/nxNSvDDLEo6j6K2KpJUQMBwf2ilfMGdpteLUng7f
MUE3QUKqSEisPA6KuPENV+0vx7FZX4S0O8JiIrC8oE9vb1itiiIcVKPjFJ0qSPKD
3yQyIRHxS3BxUZxoMGSeOI9BQeCKsYOksDv8CzFENghdxZhcuWq7cyuH6O8eV1AC
pUKMiMmaCcG8/n4jy/9ZY1NQaFSDF0dIPKFV/cf+7KoI+CJHoLHKBnfBEFKQWdC+
NALsR6nVbu8JAp42dyNTs95g6JNOHCoKWxT3pwrNqtbdKNss+5qlblZl4PCEU77G
IjqzPxzGDLbTQ3q7AbvUQiIctsQD5Kayys62ejbZJVMrucKpreh/8BZbB1drF1Ow
ZTLlTFMqrfuv4sPSZBn1rcZKEot+TwSuqa3BslCUmtW9wEvZEntO91cDhMEXkE6n
V5/xIOQqQRNc2MoCosHdL+matM++qPKgwe+GQSzmywTwAjkLSS1Q31LoBF2kiLY7
J7KrenByVxm+zm+HPc0kmuvzL6l5ipOzYH/5JbYqdklASE8FI4AJNaA8lHfGxJ8m
pcR/3tRTVgk/ed/BOrjLDD7g+XA2stLG20/i3zdIDDlMR5kwSCAQGd5yQ5UYGzG4
eiyvl0nzPC77vgGXI5YKSb02DWfCL7em1q3F6AlJb7qWMnSfIJC8Ga366KCPKAk+
/RPGImDnqfhpM327owGL0MHQPEo+pdsnn58jpVHCgdKDsmbrlOZ4LJFxLNK5n9ve
dPKK67Z0hOtXTjpvMQ1eVXEbxQ6TeUm10CjRO0v6p0Qi4ynxJxPm0b40/iyn04W1
AJtXLjDA1KE2UNoYZFbdDCtpzxsrPOQFdEBfNRxsYvpcHOX19KDqqwrgGMDoFLiw
UlFRVO7CL26o2+3ODYZgSwgFolFvae9PcoMblE/X81EgdkZM5GqpULDGC0xUV4V5
QC+vYaTF4uk0qxf/rCRkVpaPygJVjE9a8WCh6zE+tjozbsoLFFqnU4NR0u2A4sDg
dxTSvf0an+x9ZELUzT/Ygk3nce1wUpSk9AI973UQiPnVpC58KchZ7+ORL6USkAf8
ni2UfTno4xBLvSAhgqJEgk9Z+cfJxlADJ5u9Ln7enBf20B8R4zIiB8z230/xSyWO
e+1GWIrsn1cITw/0gueC3nSZKZ3KWJWJlpD02KZZQNbQQNBYz6Ed28nGw1NGwQ09
mJEp6fwhJwcdSNx5fYSUPaCC/P5nr59aRNBaGWxn4M9DnLfIghT2IqXvgNzRxDBj
KQo6s0ON4fLX+26r4ZBhgEzjYEPXajJiA0JFpn2kNFmQsvAWpVDlkAdBeR719bEW
ttsYrTFKd6iWS2/0wSdGXYXImavoWBp+d9F9Q+I4nPM7gJ52yO3F+bYDrkSkIhqr
U8neWyBX2clly82WNx9ikqsa9lLPjUX7fClwuiN+ICJEq/CeHzH9CrbThGEZ7/0V
gIJ8+maZtoxqxc0PFWVB1vc/Sclf8h8HOOnUSYmV0Y/7XWk4mLZP33NaCF3PTw1n
OKw89rpDFMu8X9Y2FIP0h1HGyAWQ/gEit9SGtgn2mA2PJpypoOfsHVNV76FX9KYW
crNYMv5ds/A64+42t/V10Tt2AtGJ1LUtLBnCqSxarNYj4o7/DjoSNDCnzO8a8X7/
n7GI29h5KH3hFworzpb5Ab19zAgj0Kw6z5y5VgIbCnzKqU7Dv5Q69UqJZjyQDFq0
cQTnJmIb9Q+DAzfdqYpQt2ZLPidmnd/noE2k0crTzf/Vit2llBNoWuvjQJxNPRUV
a3UiFqJuPQELSfREUh2BJPAO9yBOrUOvWV5dx+4OKqKS6DJPCe8dFootX5GDlgxO
3RvdSewD5zetxIgMw6NUvXmjqAaHedzDB4AGIohMyw+K75PbTznxx9Y+yaFGWgu6
Z2QAh0FEzBNtG55zCaMWPm0womDT5UY+EAJcW6czVlpps1jMV5mxfJULHXUJGOLF
OQt0+2T9F3oqRAp6XmXQMyrkSR/+hUYbQtNCiX6fXwjapJJOhZZusU/5dVes8fPr
cvbXuuxz9JkvcfVwPf+k0d/PLj4S70m+g5edZCrWvANBpZXqbgTz46Vd0s0u5Cn6
hJuvkclqbW0MjltwZXeYQklEeCGyxC/dpT8TyfGItpbNrquFDTMBnMQ26gaZ5zVu
I0HE1fHL2xseeXQrHV4Hse1K8AjDHOY45iIIvPUPA7LvJAJoRSKQpniG1bcD9huL
JhdYerfOvTTNDHEHOaJzL03DOG+I/oxZe0nV9pdy8Op8MwPXKNLJAmG5MlHWe5tq
jyvg+wcoWC0salYXpl/KniIk6hV6VzZKD7kgk/9hR8Bw8L0xhBowPWesVgQH8nG/
QLZx1NDgVImivTJfOp5c3wRnDspboauJQRz7mfwnVAe83H9E5X74tLJWXsaYaibA
snj27gF6TXbG+E89F5FJA8UksuRM8etDXz65f8SP03CyVAHPFyGeasZeHfmwH1Z8
RsSCImgsaw42zZeicMrt4KPAECzJNpN59xYDODDE9/0EfT6nnkgWfzmxDOfE35IR
O6VT/Itn9dH+WzuhtJ/A0dFU51noJTMvh22WTLo4GigO6swWk/PswVNcLOJhYTiX
TeISiD+OvXAexMOXUGBqo0SjlPVH/G5wx1QAY/gmMKb9Z6IDcCG/egIiT5yiYtAC
+XoETBSsVUV4vkJnJ4pznyruOy4T6HA8L1jggSHtVXJwRB+o84m7VFKBzC2BZ/7q
HkIvRImdzAxwyeScVhfsD225GRD0BR66eqCeRW5N8HinjygW6NnZi/AwalCUFE99
5rJaiywpJLRn8xpnHe+8WL9recQ8xt3ZlpGjC7BIQBpNB1HAYRipKV2N93dgmCjg
9iyROsYTa6UaZRkJxT5E7OgbjlZEtcz11IjPU9Y9j306whAXM523fyafOoieEmvi
o6hzCbYU9QQI5t5raHBERqfW7g8L8b8nJAtRXcUlqrk3H7r1GrXeGKxdaI93X4eD
jx7GJcTC6O4jYalhmI070ZPPtxfMvX2xf3nflMSKcPJqJcPI4Eqz53eF4XhOll2l
qabWWJJgG9ytYzUXOgnBi5yAyXhvI3WEOiTQ2/0d7yJn1Ht8hU40tRxKHszsbirA
tr0cMppLkhFV6+n5Y7d4I5v0Yc1/5tzDBmEa8SYlzUQK+Yoc2EAa8YELOCyOiuEv
PVkfgtWh28roR1kZHawpgmMbcTdF1MCu5DGOPjim1zgilV+t1T1kEevwOtMdb4NL
9aht4PTdczJejKnnR3kRtf1vhLTeDzsUKtRRIg76SUhmu+26+gmTNKUb0hJWVCOL
3ZwHeLdKOqbqyackZsvxaK8XBrQ/7PXEEUTQwuVpZiUSKSunEyiwio1YFkiEG34n
bHePta9UIFjEqdiYm0pIxgaawPCfQBTnenTOwN0DZGUQLr5erxi1hV+6rqSm1mT5
6uvYs1Wp8XDhUnIo8wMbbpwYGwSHcc2lYpF6Hf8MoYczxzTu47P43zxt8w7dQe5B
YqacXUP5awkBzz7S5QrHr9fk3/JVws7Nhk4+hBm/iVNgLQ51hntv/PIl185YwK6b
SP8BXujRsm6MCnh9knQVSf26n2Q01Q9nCMzz8vSQkvm4gRxo3idzuSx8hGLMH/Ww
VXdKAisirHU6NcRr62Fd7edJsQUVjuNj3pShtIKWO8CLStGeAQsDs8YrNb6koG7G
YVxyX0hES41AmqycoU6G1EkuQzbPHIOch/e2DqtkvVDQclU5hIKX7mbEGmw6w2TP
4sJta2nJxk7eBDE2PjYKV6aF7FXn785ABOMkgd1mtA7m7UKJbrvagBtuYQ2oZey1
xzWMyrNlQhg3Ee8VkMEKBGEAak9Hg+aZsDkevQo8dcR+RxB2y4p7iisil5JBzD8f
hD096MikPXA23efP7ZGoqm8lOQj2E7/GXXW3rXcNAdPRizHnMtfmtLF1QLpsAuSn
Bi8YqqbeoxH3RIJvxF4rfcI7Hqpqj5EmoEs0rovf36/LQizSqv8qBkvv6SgSKYkd
r0rfyzSMiSQtwMsLQiHQAdRlSWcp/0MBcrKRbWB0Dk+LZleqmQoPmBMAkmBBEVSr
IFjTUUzarvdhFt82sxqKEWmG7V4lldUeVRb94kWIGM7br7iTaK64QXfjYQlOnmRl
/ky1HOOavInQ6i7jMoJasib04pphFOWMl0qIYcxkZ3ut6LHPfov37xzhrkrUFovj
s+ONKcthX6my5mOLB/X07X69/gUjkdTx0nzf/Gnrly8j4PJQmS8PwLVzX/2PQDh9
yW+biECxt6neoF9DfBWtyPsnDEPG6srWkljavRV5dAvALvKr9js9xiMky/C+ELv+
BF1+nUKkRU2g08rMkBCZT30d6xmNP63Z8DNdUdo5ibmyT9j3n3mDwcFqlq4jegXl
q5K8fT/zQXGeghEQqbN5ksB2nPqA5cFB9rumMO2Z7dE4QxfFP/Bd9vnW9+CVqrqQ
K8n98LPr7iShYCqD2i+UykzPtK2erICYanqidPTJFeo18yVUR0czrwGiZquPZB9p
Qr5WKLvpDuhmELpp9sbAGbT1ZGBWXoIFVVfLnq3JSiP2Z4fwhQuGLkseEQBFfZNZ
rTXXZ+7PAd/MH7qjsDl+woqt1ptFVsjY2zqU5DT9q4IAQStyZoDuPjflZB1HKcVD
wo9m1a9IRSTfxG13sxLDKduxcf9HoOyFMy+IG0sRsM81xMfE7U5QWNoVJsyym/rq
YLGxRxKLz7XRXW4pCRLICptn1A8axBv3h9UB+r+9qPBJCQuq33tneX8hTjy5b+6p
xKZXnNb45LyH31GL1ewNCGW6s4bBu7hUCgK8Ryi5ZkJMLzzN27G1oJZVCu3AZ+eB
z2yHSHKGV+ALr1QhOR1BXqjjiMgbLVHioBSu9anZ4j+d8PplxcfP0EKqzVkF9vIR
ZsEnIOWgIjijlcF1EP646vw4D1tesKsy0pXZLdInYOS9YDDjnxvQ3ulfqqLhhb36
D+CJgvdF6L/pw+t+ra86hJqKyfuqBCjn4gX0T21Tg3duG79FG3vP7QO33K0S5gwJ
rraJ8PDvyCVTev4Rs1yEdtFlPE6XhSivajkzaLJ/fPV6goqK0mowD7iXswUT7YtD
k8QSoUBYt+I+L1Ji/yNxFDxf9LQRmD9Jzxhg1Rc5ywbb8SBInnAl/8+XOsF3mf9n
/VLPfDTegA8Z1Z4htCml8do+RjrtOooFsENk2vwFYpBA7/GScrk/9aq6n8LTgORd
zkqrDQyWyklqrsPucRkWR1WepshqE1hHt+RVkzWxeW8q+mIyMV3Xu+5k49zIOXkZ
Ohz/zWWYRXA7LgO0WktLDkEVg+lM/JItrBozPXzbyHIPh/BHSKlX/r9PgslaX66/
IS4gy4jpm2GVru6I0OaBaffXq3tGwBp0X6PhtXYGvW82TY8+jtljiicIhRNes1g5
vgq+fgm37zHFtOT6rnUv8bINdX0LJ01KbVEtMKHspP7NjQI7zn++EIymtlWTaeKU
7L+foE7XLnd3mR0IYWgzHTP1m9smoAxlAFMT8f4pBAGPCBuaJGi4gyRTpyCm9BwU
wlaXXd0Fh9BVA59BwpYXk3drfMi3NSbZ56mqeb0FLrvN9H7Ji+1VaOpSIqPwMvpw
7ZcMl7ujFPiGu8FeFTjVoAIhgpvAmeaM+s7wWa/SsvIDut3l7WQN4uNqma5XDVUR
wYm/Uh7Vb9ib/ddf+CXtqZRgkx3+g9qpnJfF5D65X73enuHsNvaCjkv6/ctcvXjB
9Y9RuFpUL50Rij/951KRz1BKruhzDaGtWKfSlQcNVWS38notci+1Q7ydiNOjviB0
oHd4aMUS5yQJzlNAOKOiUKjSYDAiR5MI/MZocbYo6i0JFZPCztW9be3Ijgay6cUq
hZrC7r8J7/tpR988FswDa4sNxebCSc3unp3qkdjC9m1Ug30y6RsTyolpETBer9tr
4jxM+LQaTYczWqgKTlyDNMVFw25KDrd5QxC6s3Q8evhg2vzG3YX01ekuIaN9RPkB
Lmoj1h45ouEdkgeu2xu2Our4S2wRsW/Ska5us3cCn8XsBiOVwUBuO5h2illErEJX
lzmQkDALGPlapCX0B9+LeBUg83MsjRbLN0IF6L1oVC3ELnDU79AI+OkAM/GYK4nU
D5xUZctYxMLWieoMfUjHUrtgKHw0yylmgFzWtibyL8ydQFf8P/Vb/Z+0B3lmA3ns
s2852vf4T4eo2PsOk5/SHZ/BYuYkFbkPRe2+wJZar6WHg8dkeHvhJ8I3J4ClyDxS
jHDwTO2IRLFD7UrRsxB7UuJQ3yY+BWJw823HBiPNBEUMzR0MFAzM8URODUI5655b
mpliWuQQlhM91sDnsZVcN3n6WRc1yKNv6N24ElE4h6LYy9RXLyJO6C1qDKEvPco+
MxYLl3INqtDmFPc6kV/0sYf4D51KFOs5g8d6d139noE0OKXxrkOPfCU9Q89bNZVJ
LDUMjc2mXLOCxODLpS8GrW8i3caXFeetLR0F65N6XqWQNCPeaJ1E1kAqQuCGQWFk
ktGVrP6UZs9jlngI/u39BloE85of0Lmisxmn6RqO1skwhgrpPMCgJOgpwMd2yiwm
lCE+cmuJ1wGkNrjZWyyfno2QB5D3HeMeh6NCd0wKCgw0V2x1oBPjG9vpuXUbgi2e
52u7lt4C7ASpQ5pFed+aWJJFxxy3yv0snMV7jlMu6BMWiqEpaHtwy7H2IEKB1zH+
A8cW91IFzWJ6LyvVffD6uJSF3kZr809MjzFMx9UWZA/JwMZHJDIXGPsAN+J8rQOW
wsSCk2Ju4egOkDyeLVBZ6P6rWn+71sYH4IKw129356m1arjyC69/Js1xnRcz/iYY
juUuXjRdyCuWPb92tTjodcF3gxJthfwHMWhhOmduYwX1d7r4Ocb3DRsyPgq+RijO
coTcSbesJ7I8XNtpizzdtxH0etbvom3rGYVvnhZPiZa++Alm9OS8YYZWv7Ju9Dd9
Cc0J/o2C2qp8/U7V1ItgsmvJx3T+Sg9ZY7Ilv28iLqeGz8T4S8Q4HMmmia8gS/1S
YoYU8DuRhKfW5oUuEBbYOfJE/oYJCHvH1J6yh4/IzJvH3li+6GnBCuxiy5Ep6WS/
w0RC3UchZYRakiLlr5lhwBNmMGHOfzbK70lACoO/4y1Ibn6WP3N6SYhwmAEOHpNl
vbeVi4nHYLmQ53/2m5TkqmamxwTpl3kXfFZNtGtnJX8CcaA/ec4B53xQAVyqAqdH
G/e8raXArdvHYVKZ3Pq/c+WXwDGxZ8VNIwQ+xQr+gxzqB43QS6sqqlnglzh7a2PL
ukN6EwaHJh2A3jSzXvr7F9VwFLmUFZRFP9zEWDaE3BQzhaE8dOOs+h8URPuKdLDN
HC403MwfFj6U/olLk2/onS6/9x0qTPqvVPgIZZhNVnW4iHOyqW8/WVSDbMB2ZeHG
FH/ly7R+ey5vt2GSy0kgkD7319XD8O/DGk8MWbLOPw+/TRU5I+o9EMGs52uCNXBL
snQHxc8vsLXjTbbQQ8nbp74gKeSkEs7CTyC/tsFrB7052ZFHZBP6ltIy/l096gYQ
avmVuVIH/ISdLqiIqetbtSdYJKxPmLOY+sxP3HlD2SNh1gG0umMOTgZyHjghV3YP
XDWRdQfgedyyPWSCW52QRb7jidtTc+AOdyV56leK4R8KZ2vSzDFKn3ddsUHevXYO
Rp8BZeB7pxrMLTu38crwTg+xNduBX/vSr3pjer0NxAWg/vSAu0Qg9/9Ibxk0XYHL
K1zVUFqmu6FbLXh5DuShIq+wjIIRfjAFYqlpANiNl2r1PeB1DPAQFp/s5oH68ogh
DzZ3VAFTXxXlgH05eouPGiV5H3YkiOh7eYu7+XX64vTSQNgsvb90vOo9GX4FyivF
WJI0b6AT7R0F7pUmZCYdgBndrohAeNM398I7OvQgnxA4zyZE0+W/DEXZMTx4R1LW
qFZBwF4VwnZrkWIC/lZ17Y/RE3H3dO/vWkJIBdUqN7s2mOtGsisP4JidpT9gwEGb
ihtDNot0rzB4k8r0ngHFJr3FEId7k+MQ3miDJDXFoT8VLiKwzb5Ja515AzWy4ydq
JbFeSwV+LndNMFnB2uuGIrlrfArWS20vLg7ujTzTLI43sIwRk9aE8V43dy10MT/b
LcJ8+buT+/Hpxhgx54D3zAYKYjWZTJa+kbyYRa+0rINOD3EXm6QZq1sRt7AFJ911
V3Zk6TU9iL9FcaUvtBql+cmjAJxqCPQ5hTPCWri+d36E5k39NL/6Ty1fDe931jsL
l6JmYN6qS51viTC/fFpOmYc9O+nmjgCxLbxSev5GuB89Es1EAZnzSnDQXtsp/p4s
0tg4VyBs4Exws8AypiQfnzkhY5MXJGvKtv7zqYGxlYHt2EzLxd7mZ57HdWa9hrxt
tfp37JReCbfGK/K+i+lm9LN3v7FOwooDT7tir8tTX+sCQ8SCdsWt4hCY1tkP0nGQ
zGjWzAE8mfMFxV9uN/fGuN+qniaOLBGuHPAdNgHLUf/88rXh+EE1kzBnGDl/qXxA
Ul1G6YT3DK2r2cLoknnciaoC34+Ebi1w8yxMlW9OW0l7S9/a8HeJyphsSmq2s29E
QooUf3NfmV4FQT5RIGp9H+8bmQi4Mzalsa6IRND2PvCqhCw00qhtzwuY97IF+YQr
JkA7JI8Or5gdBjXJywq9p5sD0Zq58XSXx4Ev9Qoy4z90n9rBWbBXYqqqoGjZJP78
BiSQPmQi7EVziSfaLWac3jHpqFYj6VouOPlM+Sb9011ZumJ37ebVB5/YM23LRwzR
g+xW4Ub7ODScFtfcSBBIY78IbTon6p0HwV4c9v3kAndq18bkSg0ltI5kcHgPcZ6h
Q4LO/KDZ3HxDLUQ1/bBOY6nYmlSOAGBy3C0w8xpO6G1lfYMcrJ27iNU+devs9JXE
saNwW2yJVmjL2krzs2n3U48pJWtq+vWqECywrIh0yD9XE9vDPDGsawoxPnXPrknX
Mcx7x9UsocyJ5PxNRGx3XXMhCrsSs2h3wAJOYS2kcvgPI2XtRO6UO1HwUBvwfzWH
eJlAdHy3tztORDYfh9yJv0jUAvs93ylyucCeQwXwfbe2Fh4H1+ymnD4MV0eaYFg8
3GxYdV6rs51gkd33uGUrFXm3LDOUWhHy2C7lcVeHYZT1kFGE2BLgnPY1bpD3oc9U
kD3Pt27Em/T+zaByAgI2ndafcGL7C6+I27eH/KpUH9BpeAx6jq56IGHWLVbQXABk
qOVNHGMhwSx3dcACuJGbdP1xCUwiOzq7i0wgwBKghM0Wd9edkfvOmR3xCDqOKMOU
yaK8KtxQuqUiaV+rGJFxuxUEIh77vBDPT5ULR5w2XYr1Y84ed22zSAEGO2T+lHyJ
ZdYijV+6yAawGZsbMVFyHAbq9P5YhrBDvYXYEj/xKGKwM12n8rDu2HSoiIHXFWzS
vTp/RtP6kHLz1QiXqQjqu9JCcPS6ECn8/wHnhkQIyHUFTSyUZH8RaoSCgPpZvgKV
l4kjyDlnPB/KmtBsNmU9jBGT1yb1GzVxPSvpPNBZPqMbbh88qA0Hc4cbSUxHTz++
Ibe0Y6Sbq9h+P5ly/BUGOOPBCy2ELequxrbhuuiYXPlbIM/mAMshkKwEz3Cmp0C9
XwL0zakJpSEwnQpUu9DT3QJQjSPdWyhSXnmXjj2Wj9mns9SJ2yVJ280h80PFZfIl
utfFbVm77AX/vIEaIuATEdbxevbI1TEY8vPls3tQpTNoAGgGRma3xdxG4PficsRQ
VojkX2A1HMoyFzZt5LW+E3y5xepKbKvVndnYAW2nTeqBvZL9UvgWT+yWcERzCBeO
F9adL2x4XPDw88LLvhkim1vL0NJXvyby8hI2zZcYhO5Ni8Ym/zCIdcsv4O4SyqXd
b/nW9EHZXJz4uzmMinbtardPv2YfbCMeUY0YpQGw47tPrZb8CpdpIPfrZPsvGqmN
Nix904RpvZgo4kTxMjderBwIDqKd664JyH/qS8XSrf+AkusnRLM7KE0YjGwayFOX
MkpgkvWZ2W52/Jiura7KnkRRK8e92gfiU8baIUJeX740nDxH5mfoAVn8Qx8oEm7R
6B5uJm9+u276KGgVlpdOV+gaW/e7sssjjosauXFRXjOzE1HYfVyRhMWPZL37Dcsj
KRKzaejTwJs770bdxUl+fn+IXUGvjL/JDleJDofTS1MEynB2Y8pGkRbN7vvmWkDX
VMu65+zpqLnzyPgpMjC4+naAKkPKtqGf9FiFNX1uxgDl7kzpbeXDbFizXvBHuWxA
4k1xE22jNkReCSKJBIwYcX8WkIBNvcRyzs81oWas5WdhzwyaKbgOZDnpolRSHOI9
FVMvJDGHcsXyRz46xtvcD1E2NNdhn02hMsnae3QWhi/Vi9LfueQ1dW42jbUATU1j
8iIIF9Hcce56ES8xhsNN5ELI2oV3CkU3HIpYm4JrV4iZk2uQX5ZczGKZ0nToFOAO
oXGQE4WU+lKKH4CFs4RV0JOP2mgNdI/4Q5T4JsY899o7EPFKr64Uu96mu5C4Xb+8
JZkf7SUbVodLxfR/sluYyxbbXybALZre6IeOtTcZcfJM07MFTslVowG8EdI3hZik
DG/r8azpZ1mmiWhcJ5mCAph4n5O4Kgn/O8r5PG28A6ujlpeUDsSsIsQZSbyrcfER
RHrHhSuKqmlHWwPklIMjVi6CH8SEfyLC7RrfXnkaKI5CMo3LezoMQXsja1FcBeCX
zVWg4fhyktSyNWpn1+Oi5926D69/Y+5Y0uK1+b7ZjMndUdjeMkx4BiV1nIYo5jZt
TuMomoKPuAZCnk+/Uw9UTxGkaFk0u4wiCbk1jwWas2POjifptMdZX3f50rBsyOws
HLGAAtGx+geVdx9FVXYwH72PX4is6s+4BhQWgbcESSkOhXLg8C++lA0PdVSYm+i/
Q/Kfsxt1f7KwBR5tnL6uXQCm+2qE4ET1Cy8Qg6wFdLKUgm3BE9hlhwTdHvJW3tZb
02Ygkde1GQqmqXrqFBrxGbCm44V0VgsnUg/4L/eA1bKymK3z9PNohLsuBSs3A7O+
zrDGB0sOIJob5+vfus8kfQzyWPYJYH1ABp4h0BqLtxrZGq2nfPuyH2IyQWoAMR5s
oO5RNRhfbwh8BOhf/hUBFclglbDSO8MYFs+xVvKpq9W5jKzvX79JKnD8V9no+yo6
TXXDP4xC98RgaCQb/YycxgfCR16AvZPGLpTfTFphaLvigkxV6hB016sKJThTYtZv
XtEoFbSGvteHVP8U7CFK8jR9anXq2zSNDZk4LQ/mLQDpggo9OnRXmUalYhYGiUaI
LsXBdzjkDGBC4XjSxPRwI4fbjLF08ECRGJ5dZRJHg1+AB8bK6wXaoPXaAc+2lUca
paWu4zYBP4gFjVsVyPfeXXLEw1TkLtgELob/MXGlCqhyunHOE5zgdVkGAGXLixFK
0UI3bjl9khXBndeEhJpYd5M5zI1RIltA1DG4paE913OutEH2lvn9zwViO6r4w9vk
VwS3qAo33rc3vNCl6mc8rHI9gvfmUkzc7Mkc8gcORtbDvs9mEGGGuDW6uyuSznn/
n0iO0D6LkSZu+lQNTB0xzOvL+FlWmrbkiSRSYo0qMU3fPpnUgUwTwL8flNS1RbWl
tiCDR0ZF/DlRNqUv+9+9urz0ygEGWi+isrer5DtOK8onYKv1FAPRPaQ21A/5yGGh
33bwA0TgQM2YXj0dISozM/aLquKf/0Jqzl/wnBSgJAsSWYFvZ6dAr7LVWWNvh+3C
JbqXvHngHlnlRgA3OqWwshvmq2yJP8z+KiHln9e9NPRdxDCPDap0VLnftXhflV5J
3snJfhaWyCWdLAIzgvlwUnOX2cFKJE7FwIjXwSjg+WMiOvH6HJwIA7NhWLsjuwNu
IbhVU7225uolMzioLUEHWfYLFgR6v7asAJmBgUP8UC2CtX9NM4qByVxVKYjmlHw9
eQepny5vEU9hvftKSwmsiGq8oPSBSU4Tr2R+h33VyasMOLuyQmPS6JB0Xvh50xkY
+HC0qwojQcmdDfDvo9tdbCtE4z5rG0d2LN60L13gvJssZtVNRXl2+5IEjGREBOJG
tegcAispe8/gWBIB97cNXAnAYpXeMNoIviAsjLB4Jd7/eQVMm9tBB672RbmnFp3J
KANQYRDoTR4iKwGY7Lxblb8Of/Hl+yMUMD/S5htfVOovDvtqU08WmFXEOjIvtEIV
Zqkad6wo90lcvKOEmoJMb3Nxun6hLsNhXQ8gPa1hYICMaNUEi3Qrv4uu+qitzial
gyCj+fyIi6c7BGXlQ3nwBnyqjwWJFpxI8vqYb+bUkUCZlAvw69z84juut5EV+yQf
JmF8eWxnK5VuvcvmAtXC8SUOOo2KkKsXUh2VWQ7Wtz6FebyBFQqhwa75OppKeeNg
l1sow0io/eD3PtavbF3oSdIEHzti0KD8pZEbENaouR+OnskWZVbITt+nMGBy8MTt
YdtJaBwE2fyfnPoFhT6wRHy57trB6D6kzzkZNM2U04wFeOvj6XZQId55SJ2x4bMI
qRqaDdmDo6fmmBRZspbFpVxlFq+BOaXzhVkpBk9Q5Vh38T0PsKuQhSB1bCIKyAx+
wRvaGmxd5bAUuldG9yREh47l2X+a5tMRrG1j2yE+hrYrvPmGPAFu2fp0Bp4Z42pN
v+PpS3uzpFeGJmg06zzVzkh63E9ssrwzDeaE+5eg6hv5K7dblcW9So/u1+IH2xIO
UuJ35FsqZ7+2+y5r54cWkeDxf/wRn6/udA3jiMmy0mqgoHlSqeSj1FIbnvyZUGzc
6WkEPUsqGGQ2V9ZTrgwundnrN0eBNM9P/TsqIExX0U/31s8HtuxFliaS9+qNTxgW
x5ibkv1vic/Ug/Cr1/zh+J1HKJjnvyEYhldhXMrqy6mKDpjcaqF6daGbsvSq5k/B
U6Lt1GnQ25PoPhg0ZdBl/DtT59qFxKcVK2XMUwluQaFb9meDFTLieYU2KCNDxIWi
GsmfxioXdxHt1FC5+FGO0uXN65Kc0ZbewafPTf1Ri+E+iqsUw47+9NN3iDC18H3X
SmKYysvbB0S4laccrD4OosiUxGWX7ClpGXnlqUSh4rHWSfHQ6aZ8GIv7H9LWGX2k
b3dbnVRedBoWEk94UfzhKQHNJLfpHSZjpqFjbYFtZo5i15Fx86p1+DwVc9AU7/7V
cp5k9339ltLkRa5Yq7NlPkw7up4S/FHBOtyDRX7ZMIl8kOkL+tm+Gwy/MXVnfzWJ
Q7n2pN0Vp8vV4utN4nVMf1kUp+e7x/iRtKeXka22hOTVjCJ8rjdWFZ6ly/ef4/2f
H5J4bOfH5niZLQcqIK0mqQU69+4nhOLC/298Yhi8bDllwKgluwQe4I2Mtyr/wQgg
UM3145gDfQc0HwljFwy49N5/DC9ntgleWGQfVxNRzkWa36G+msKG5BCC+guqu9o3
8t+EsepiIo27+4hB1Tm+8cuVl0B9snZWOZ4AJXeGsO6FeIP6vKC6illYLx7SEhx8
Mmz8EFOia35nuViPXRwk+3Zz6lmaL8UR+8auWjbWWRbzC7WOkDxjN2utk9llPHJF
CLSu3+9dGAQL+rIhMPSiaxn5vtoUF5iVnLQeYVHkn8yuV440puMv9f73h3Kl1u36
rgx51eh6qn6RLcfju0+f4Hwi8Yx0HUHV6jDbZ3YkEzZI+BcS4zi85eGeYIV0SkWl
ipMrES7uH6biDd2SB9iNM6KS8KkwGgLoClEiuyoVv+ejgM84+kswwN2FYdxkq3LH
4claV1qTA6hpl3FMalzr338ycxrhrqKraDm+XxcZMC6hfvJfe9PaN9qNLTONSpoX
4tFey6Hm1u2SboVntA5GvZZZIs+d8nmXAMAQgvtBMi3eh3HKAxNMJXhZh4Gu6fGA
jt2jlG3yjHYA70bgwYFQkJvIzSICKNQTZ+w2CvA9Th6tnj/WNPIksrghnFMlsOQa
Dntk7nZh//KQKndWKkhhVPOVzw1NPHElnjnkJheiKEdJZCvg8VcJ3OLAmujNLLNY
Bnve+GVzUOjWuW4PbeETeh6l52L00kl9stxAAWH2X6UCr6sSrH/419mSvBmNYwtC
ZqLjHtcLdYuXbcU1M79gqgIWOySYBN3yyOHb2STcsd52SulBftr/BIj2U1diQzrN
CmX53uG2W/+U9KV7xJHleTYKPgfG2bPyej2CwYWiH5NDQiT+CU8NckrZveE07HLg
9n+G5RPvddPJjXcdW02buaKf1QqiS6KLtsE5bv+BORGUfcXUByVzqKeEHI9FXsEG
o7fJvCcSgCOoQvMnZk0bHX0Kf/7uK/u6EFj/j2rSuv5jFtZ40FzkdrlDckthRLty
qzMwqLRaH86YA5MlbyJ0EwmWTeMHuEvuyunN/YrIMEi6llzJ9LpjY9w6pMStGcwq
9Z5zyullsrrU5pLCeJmYD6e0NrORN4+c2KG5wNmNghJnjdGXDUitXnCPHmZIoQpY
ixNCfj2nP+YCUl+IxLdKf5SBm2VFmLtxxNTpKFt1dyOntQ6JbMcF1TmTASa/3LL8
VdQvTbFtBGPWyaM5AWyiMSO/vkLkbePbkULEpqweFnobU67/t1t82PayZvjrjOwo
7pjS+6kLf11y29zG7CgThEWP/b86C09I857+Lv1BOiOUbO7cQzEXoeTjN3Es812s
yw73z5mDMHxczUotnSeC9Pjj4DJvhSFVtVnyKb4V792wryxjx7KLDABmqE1liU1e
7a31og4n7DF+oij96F1Gw/FQDKQIht+5gReSIjI8sSA52KWpFAavCoMpiBco/JZs
1os7c7yb9cWEAPZM2eI30scGFeT3wX4YHgM3Dtjt22uyi1ggnuy8M5o7dEQ2RwVc
TeuXX+XUt4y5UBTrD462VC3+DlitL3O+K0EzmPVQMLrt2QeXZ+gcfZIstDG42vqK
/uYPjMglby4GHaIK+Bvr/MzBHaPqWp1KM1rOkRvDsvNmNBRWbiETJTq1Ipp9B+f5
H6OZhuUoLaGe5I7wkeg9nexfeIU5mnoehKVDiFqDIBt8IDRXb/ZK6YBqY6+S/6RW
0PiS1PJ459Fc2xcIcGI7Rf1eFTyjnKEwomCto+5Eq9O168ERFpInb4b1OOf028wf
yrkVzMiu8ScwoAw+xyME5QHMZXIyTnCrv0eoE5UtcKcuJuSR1KlMwL8wXJI0UiQm
Ur2BRdDwgPviOaCaN3zJ0HAyvFP/qb/26GuYGwHnYi2MSzgn/AYI9n8Ggtz+kGsZ
bCto9He1XdLdCRG5u2xMI/uRwTFLrMY4Z6qnLzff40NN0h4/aFX1kTfcuMfJH1Xb
zd0OhJzYNVCMYH8gSkxTqOCeyeDDtsoYG0P5oz/MXIDZOoBOIwS8pKLrln2iSuKy
vewsJWwKablUjvVxwDT9SyV+PfILCHoMYZ+vNE98DtKqWJAw2y96WJfGoIIOJQpr
MT+bfNiHbCM0Nc22VXBjYlrUD2JSiXaSWelAxP1YEA7TOPo2hsETNjbci+ivheSG
O+XY+6tfBZk6/s2xPHzoED6N9UW1wRoh7NtPTLdqlZ1Odi/CHcV5ne+Apl53cMLZ
pdlV5QgQeUFh/Y2nEYclahR9q36sLTzOGrFi/rz+RWlv+VSH/+ban+uYOX07aSx/
+qBQyePUJbhcPf9yjCYX1vtreIL4rkHBAvNqFtLf63fOkYfJLM/keE+vSuR/a6fn
dO02mk4y8IB+wDAMsF5Fro8Uf7jCEPvZtclFhCTG3toGsL++/R4Dr+RkWsuiD2PX
eE+VGAfy0t69P/Rnt82aSuje8QqAEabGXBmQe9YmUpnE3PqDcenuBCDtuRjUmP8Y
4ppzYPkx4QvTRx3wXynsESUJ5emLGcSdLgZVdcvXjQsMSbpY6Dqh1U+iPSz4e0N1
NaUMOS37u2sQGafxFzc9Ploc0lgbKVOYnQ6BFCyhBBePoVqHzlFXG23AShB4nL7z
gliFEItTR/hSq1s4FdIuKRKzPynvKZ5bI6M3Cqzn7S6HWRdo5Bbna6TlANXu6BBr
y+OgCRXVcWQLXuNQRh7K8+rBoBzw+jdoh+CbQ1kAAUgxgUpCZleaoSkyZJuISbqa
Pd/hWyQVLEZWhF4DzScbog==
`pragma protect end_protected
