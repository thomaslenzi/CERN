// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
enL4gH8d64zsR2gwWNmqXS+6CVj1QeJhq9fEafSaCpT86eplh2cwV9Jum21DfH4y
/b4hcl9/G9pf/xIrRL06Hw+i3izOL/LTE28XjLiJKv89hWlu+TFxqn6vr8GycBWQ
kRe4FIXgSbDKiH/zvW+rSLgaKFuGpDoTQ2n+6JAjdIA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 128720)
fUcU8dOs6pz14lkn/DNh6ajWEORkEe8TEBvrrOTwLXCRwpsje7RJgRXAMIDCTPRx
4npbgsQXYw8EUl9wtOh6Nf8RkysWUEThuzi+7pHWOWo8Xx2izkTV4SuZXpQ4a4Am
T15c+pfDhHpTIPqQhjR05ddb1hmWBo873B7/EFG8yzep3qzH61DUffy0gPZdmTSs
pY9V8butE8XTRBpJOFABFmkIFwl4NfNJP1B76uXSnXUOyhf6z8BBfO0hIXGrNSTf
TwPiu1aRSyAH+Br0AbvW8B5c8YBBb0wTAtIBAdRNi3JcGRZM+dGwHL8MQs/0a4lv
0qI80cS/D9tg/ifuFKTYS6/EnXi0gkBdssJHz28aDsLY8SCSBDGHav+KQoe+qzIi
S0a0EVyrw4EzcOd0E141ClhM//TiDJu/PQ079zSzAYKf/zEY7gV0Twxd+MJ9VMX6
fz+YPGc4wyWn8c0/PLcf99rxnGx0p7ER62+opZWZerODf5xSQAV0FtWYk8mDeOAQ
R/ikAc6yCVPgw9kVPSSzBkhwD4wpSd4nulymNPyAXHR5yao0olWJ2fLHJxaNkZ7d
rVJMUT+BCHZeJrad+d6H0D5vn10AW0KkEj03gHFJ1NqfM8K9lRsOcOIX9SluCJME
DVV4D1sdmY69/oTZEaTbexa+WihgRWEo/mn3hexit9jGYEpx4s+xBd3XnR34ikXz
MSLGOp4tLdNeqZHlNN4Uum8DqCiF4wPzqWSnrVJl2lIwMbIUvBkkENEyNY8L8ZoR
pacwCzDGvpvD09Le6o0VK5FZyiEo5tCdo6DjCXpQxOuntX0BWp5pjsHhmSLbgq/o
XOJMUHZSerPcoClJ/42BGfYgm7pi1UImRAiOP8iK8TFJyBPDkyRSF3Lkc3X+yJwL
+W7FKERVghhksUBureOiE3ZYRM8b2C4UI5ozD6oxC+ae19FX4AmpMqvzK/9xjHjK
wAC1uP4RXY1vnHLJmcnCaklW3fBd2OrfXiFAXWxBJW58xBFA8OFCD1FPmeaz0Hu1
MqpvI9ykGjfT69LcMjDfTeHbF5YxRomzYN3pUt7lOKSVSL78wxHnnJzuzywbb5/d
076tBCCgENne7TjOkMi10u5Ohx3f4tJ/bPP2Gl4fMO0Amdf9d9I1fPf2TBG8yVV6
9/cNJRHdxNLKqTYjqC4PkqpmAbgP89qF9bCpekT2QYH0wnFLR1fPSad/v9PCIpma
XV+INj1Jk1eXe/tTvMI771JBRPRpwR38WAHxNPxxN3T2DDeiy2mO8KOz2lHav2zD
afTi0OMhnENLBefK/7ZP+D1DndivOLUJdqzWhXisabIlV0rpD5w2VPOHFADIIFdz
XJ0GMon/WVMbbZeIwKih6cHUR747lvl3/63tLNWVZWdXHb9ui0xcMEB8i6E/ZTQc
fENhUOpVlTGd3Y/TthcEepacTICYrNG5nIsgUzDfYITNuuu4YVWRL676rRpp3250
B3PS2nUtnGZqdJt+wA1qQ7tGxZnlb8l0ECDBIz1glvzJWL4TwTzjnwpOzdoY6+h/
3fcyo5CLiZHker2hsIkTeB01N1DyGBqNiKtPDOomBc1BHllRBN0qUMbRmNK2zue4
kBQGDxpjnH/0SJ3M28rLPcZWS3DTgypc1ICHv4U3cVMeLhuNVQCdUjK6tzHd8Q7m
QNRrBavBbNzN3hxpYMoGC7wlv4ph8sbk1RQ1RMUcB7+RSEGzGbD2bSgpNpk5bGmW
bg/9U7uiezwPCL2sSnvYAwS83pysPUqjFFqYsbJ/xrrRRyXngoDxs+oB/jzA0GU2
+Rfg1kuL4bKHTf6aMeF/Ngdq+gEQ9xVeZdjAWliKhnfMf6ZlxQDGs6HJ28jXW2SJ
xjmXsDTnLY3cg2t7S9NxlVXs/pHWjl+PZU4Ub4zR0U47r+fr+c4/e3UeuRr0jEXr
mgMwfspN598yB12CoTN4hjJj2EF+BWH+6WGQMRm4CQkgxVT2z+PcPcNCqAfj8tF4
W96Ih/DbOob+pohLEGr1HJrxMgCQ8Sdi0P3MtVCIzf1gbtHM8fxrpeOQWGhw3Tcu
XDoQ/IvFQBq/2gqHCdzGZxweJrleVhxCZ1OsdYogI0Dmg+DrDrDzHQX4kmqN9Cyy
U/iI1vYl9OiG196DthD9CWYmb+9/wqNVN+oy+wghkXvAcPqhGr7sRpdcsDegMf4V
MG5pUmjRISpv6iTpujM1WOck/7ABX+Ur1fQ24mSI+965uN9dM2oq9nImArBRUCqz
gsx+mJo4J9kSH7ki7Z7IYicNzFfbk1H8+WL+rUs8BnY5JIrnk8prpEMuHvJ09by2
OulLsTcHgLop8C6DiP6pEnQaJDl9i3rrwS1S0skHSSm7h4a2l5PExCHRcHeALw5p
eT59F9I0KG8BhPJ9+3LnDYPP/WWg6eXfW5kO3ruO/K7Oj/YhfpVAUMSeXVOa0yTF
fcGgFGxEYIx6ggI9ZE0cRBf3Bf8H2q1k8EONzaWqzF+xrwGXkb8cWy9/RiWK5UPg
q7ufX/EWP+V/VCsIgxPjE782Ot9HSzQrIegaoo4RL5kQjqpUpOgZnGi8NSQeOKMe
7kE+5n4xXGsn/08t2jG4dLSA93zRZpvFmV+niREY7NwEl/ktUhDJnLRQXsiPgUoL
BqH/I8UJaRNhoodyXRbqB4VybCUpmHtoRvQ5mZKt2UyB4hl6g2ZI2cjWxEBylT2Q
p+iseavAOc23UTZHQdrvlTEkiQ5RcV09rn2AJtfchBbTXkWjpu6ZiUY6KTDfe01p
9WVh5xrzKrE+I0LAzr6iS7Npa0ZZbyaNgDxVphYfKYciVUkR8Dtuxlwim2qL4/ZY
ALEZCdlm+nmI5AJEwmAwnWriHaHWTKtnc6HfJXCoBTxzSNxoROwodX8koRdNCO31
VebHwwR+pO48hTnPswSbyvsiPPcvcgODvZboGISwtyQ+G7Ulogr4n/zJu2ERPwW+
n3mIcS67I8CHSAuo/9fJMgStsmoCoTAMolqRfOECtG/tRlqq526YystLdNuGCTbx
2si1q0umV1UIPI0la/rEsY02FytDgnDOHh83TlRwwb24DtdGQEUVOGTQYCsI8XsC
1/LaAojvf6XykvFgt6sd4cRKG68w41XmOsSiKHmWwk/wadcWMpBwRKLseRwUJqzg
5th5tr+AJDOHjfmCKK1qZey65QCzzKdyHsSCiDVNGrnCGCXbj0Dw/5fpep3yPqfN
ZKhzz78x7AYGG1JY2e7gsOYTAmdd33SKTudL8hV3e4aWT5K7omuBnwh363xFXdhC
Py8JT9rkJgs/adJk2SqB8iyfaShxa9NKtD013n1Zigtlq0iJWRlDpzC7GPRZ3rhu
3mjrdWzrPS00eYVFlu4yU2xxvIKBfTwx+AkelNIvX5LTLRT5z89BnXHdEhYtDDAo
NWF14ZeatAHUFgQn6kgkxsdKWW2kMtgyrtdFtPZUdM/tlkLWxBLk8t8zKTEgSBuh
L49TidAuARE2iIhrzL3ZgVEFSYvRkbSi8gkDA4OU9WdcNkDO0+wbtidAo76PEfZ2
dvoow9pl9HNtQnQ5ZS9LThfgm5q/p+OS3wji08lV+rTg/vg4b6RDHrLIwtM1B4V6
xOG0QnM5M9cOb2QcfkMbtYfHZzo4hwqiS49Cb3PomREl2o2tsdZJGJyz2j1sqc31
BmtTgN9G/6UAmyEiMSsZJK8Sc0WDcYlsv2se85nzjMzqZlVm6j3UTE0xgWorxxgH
H1qsCBisTmfs2zxOlCTy2t1y0qUFO/sEMIl19EQTD58bGredVskPFjfaJ50AJfMJ
3TpLrH682pykF2kuybD4pxN612A1kXXApnk5kDQT/A9Y5pO0TDLAvizSiyZN/4lx
tvQJuHVCsjjrXiajv/iRIajDwHw0mhgPUAQh+NSV/o4lWw287lsBm8STBabbH4gV
76LXp9xc+N4/iawFf+IwOHi75ox9gdcXdaNXZQsDnPpCjl68IrHg598caY7e0h6n
058XejlZ//en5dPeQUFgz46NNZ7Lqic4GX0stR0EVCpIj4tSI5CeqyTrQgX1JJwu
Ltr5sdjvaG/Md3zYIDY3kuN2tK648mlen4DHO8LDKUgWXUN9BVAH9a2fxMnMgvvK
fKc3crcJfHNNAdEs/Yg0s6M4GNm7wRoEdFPxFleytGKl5RIu9caZQV7iNJDk5E57
lSiiI9qn+WlGtR1GeLVx/LvmARarYssQe2zCtXj3Gs2x0IQQXHu77Tq+UnBZCzOL
vlRhoE3M+vyNa+8cB7sBLvSOInmp/KSZg8pfDkLXaclwThMHIkh96F9wnzCsIyw3
90OlaQK69FP7QBab1QeNX2WA5WoK2J17hpHUINR4DGoCaj8CXU5IazgTnaWPeqD4
hfImPTRVcmQiD6PlYuTUu03q2HxrgYqtn4Uc3wi8PA7R3YgvEce5Osmf5wsNF4j5
pAPQBFMaz1Yz7/xDk4LpSq1/IeA//sW947K5zo9/kqfZhNqdCv1ObNtPJ/uHYfyP
k+uimDxjoUtI4gtFKzScmfW3FI/6AtoxMdj/Q0ky/U1qTG8QZibt4VV4ptvY3Qy9
e0HjZR3BdVWbm5LpdtV6Eb3r6SjXHrVNNULni2/TZ5Dqg7se2/pMaH60RtWwPK2q
aHtYT++KbTe1tX23/sq3vA8itlncXSTac4XYqFJWaB41Jbl7oTQKCK95Z95R0G+K
y5TpLAuZlR8vbbkbeK37EdTwRFB6l4ZhA96bkvNCBaKSp9+SwIdMwy4uvDUGdotg
MfDnKwDYi1s2R2OnSGRhAcVg/f4o5h1/02a1UR3biAKa7W34KBrVadNqWqEwkUd4
eYiTKcHhKqTtO4Jd9MedCdFtgvDm9nLAw6Z5LrhsjqfvDKIz5rpHAcklYfPp8DTR
qKpWpOWn7LDdGD0kmb9SCYBsTPjpZV9NhOVF2GuMBL1FydKeSzMwMK9PjzGAkzlf
hebY6w3SYD94oyXUaPMzCoK3MZSurtKcurUPWAP2Uvx7dXh0AK42FhR9BgsqxitB
2KjYq8PF/814ul1Hm1iZCh7GxuLIqZlbuUr1WKYMhydM3bbzhs8VApZYgbkiPJwR
2jQdZyqDsqqfsdsqZLY6O9ojSOiT4s84npwGcsiNJLJlAn1Sz/8IKBIk0nFnfgmj
vH2VVkxUh7X5nAD28t8cF6Jw3dz2TAiL/T7t92OV+CeAmo26/NtyVTQEn/QsHMHt
UnZsjesGBfqv4e/u+0OdiQQFUDBH302r4Eeu3anJEvPNO0/ERySZLkjMju+P31UI
it+szAp34OyRd3IW4e68tHZ0yK3wdAEbhDRQCpbkL3dSibCyRN19Lohv+SgfiExF
YlhV2SLiZkelc538FF4NCzDRny7Oc5JqNDNgivVJTKKb3RHv0mHQKQigDCVygL60
U4Af2heY4UTvtHH77bdksu0MjBFQl3O2+3qpzNAIoeWD9OlHHwu17QVnOnIIZxT+
+O7foOKccbg1iIFw2CfwngPgX1s6dnb92dqIicj1vhtn8gRisMgpzCOhwSS9cCFi
8pzBNtkXH/QLvsNvXQHMoa1jcHXMEBOvnkTV9U9wvPinle7GRapbs4l+eKKCEk7G
4r+VRTOHeJXe8XPZjfAWHeVdpGQhZxGZg/AoIA17qPKcvnotb0l0atAW/HEObCcw
LKvDAzw9EuFgheuyz7TwPIGN+8vgmV3pdZswwRReT4qm5AqBhoQ6ECdF9AQgAyiR
GiJKXZJ5CBNnRgibm2Z/tTI1B91gvS3zhKm8VEKzJRxXXrXCfdlQmrDZWt44NB9o
T2pZdDT6jslALhWbw0EzydMF6XNab5H3MM+FrfbWyx5wXJv/upsVn2MnM0thUSbR
ZwRP1qzArkfEDIR08QEr7tnGleaNiVQznyzEdHFEAJSNsjwiE+gogDIAotizRpsY
4rSunhgqc0scKRPrV3nKQA/h+KkruNc4n2tjfXWmy7Ob6xJIGkBtbCP+QCxVrImF
W8T+QedzWiVCX6Kc8ID2cDTXPctdtqE6GJqztkq3BxCCatpklE8ve/klcDhWSSDl
DKJJIo9Z/hS+7464KZP0jAZjRuNa024EOXcCzl6+LptQOVRVNLJF+iVgDPHZo+se
ZpZ8ssu1D4MuRg2HmclMclKHylc9x8LDMmIOsnrtzwABPLm2VEeLTk2c4Kew7x2j
VNuQbFed4FpVmOO3Xc4SChRxcfdRKb/GhM8QP0/PfoDVdNhG7Bu6rKSq2AnPWfG/
RrMwAsHu2BH3TQBhGqnNjJtS90sX71xvSmIoLjoxuvCklh/1ru7dj/R1z52TfvVC
k8xYIgr3/hCgeoN93KOI1jsKE+dZP37HjCK7ttiruBCvXBkD2u61xJNEmVof18pf
4YTVsRvQCzCzuHQP9VyTCZPmQcPBzicVlba+Dsr+Lkki54uMuUJ5aPcddknNfLpJ
NU9FOPeqFGS9urjZDFBPojl+jPxYEyqoomRRl9rSEzcpc19TlQ5aKePGxM/5XmTA
juyvj1z7QQknTuvViaKf9uFLUVPk3rqCEsgWh2zrSnognbz8S9uISoJ5goEHmQTm
qlXtuBkdoWDyAD3iVJUJ35Ve6mhIitd/v4hZS/kH5gY3RpJda/QkdN05u2Jomlac
WgAXLkzib0GK8euvLRHoEnEzRsCuCqByoTpFVDNyqbiN0kyPC31+HGqFpVfzo6fX
a9KIomAxPigPdyqXlzjl8Y/trehWx4XDvy+m29el/dOlJdiuS1CugxGKsAbqU56b
LdUTwc5ajj4O0+EHhnolQz9gBNKk2Z2ze3tEADLxmv/BEenetiPvC9HZ42/rO2eu
UtA1XxHb8rd0HGnhlT0KiHMtQm1PqjmPvoG6RaFFK59GTOJxSpxEB3mOGC0H4i2M
oyguUP7XFUBFfykrmDMOOdtI+7aTYl8pZcxz8lcw1hjGl66m6OkpUnIzm/Azf/MW
PqzGSsmvjm7VxEc0y6n8BFGzSq5zuHONxf06tzNj5l5CY2tLD3snDdSfEI4JMYJi
kuOnJyXjlWtqs/zbipR1jralwpZQhuyQ16cz5bI0f2ixBP7tfw0Ht1sEMCBEw22h
O3/LHI+jY2yqTfSknppQ5WlqOExeNtgrm4pkyLmZvHbLdAOEMV9QCIk+4YTmLDns
XGXrZp559iG8PT164Ms309aMV+U2pwNBjL0WSCUIXZRG8611FvD80+0OnDMGV9+5
U0PfQwOTGfBqQ+fO/R0TQrPzfWoPYdmVXmMPd2ibZVjkSNDcFWNxpX3aZCpWxJRW
pEb6mI8aviAt2F61lAMgxlsqpQavXAKtgMuHvAjsySrQdIx5WmHloCVD5A7hzgv8
f36XVPcPDmWOdrL/ozafB72DGJK8zvp+AYmR95VfiWCxhxl8xVNsvV8eq12ExyGU
MPUvkh6WjsbBQEC4dSpO4XoDZC7+C0Wf+p/DJkHNmhCR2C4wq5WPPPv7A/ksYqHd
O252w0eULSKVMr80TmRPcPtjpXb5h2vtetnCw8juO5wPS6jXRo7ZphvoxU+mOwyl
pb591q9wrSO9XRTT3s0G6qSBcfVXXkHNO3gA/zp5FYIXFI9pXJzt2JIEJ9PUOBVe
DAzOdqafGm4Qvm+q/S2nRUwyg1mA6qIkw24qrv0jVPmv3W4r5jsXqdmpeDu5qFH0
3UPJsyY9rWMx95XSEny/ZEAZh1PY0wzWJTa41GkTtuMsETwa7wxE2PHK8zWvvwY0
NMLYe2VH0ejZ0jD573V9lJc1fBPYV1VHzg36aXntN0THMqzg353NlpiIEi7dsyGp
GDn7SETgZPGvU0ec7GGMplDf5pewHrvM2Fl05skxnVQ/R/w4858WGlt90rThTqIm
O1G3zByJTFC2/fK2UXlqAsOnrdgENsm+i/ot0uGBFWWFUgXZdVFvXEEBUBmoBvks
vA4cHFz9ySvslRJbJ+YSKzOGxiTLKaSGQfq9oum8ut0cBcywR6g5DcdnwocXQACr
yPz3Wp8vbSSae+T3beJ19wNZmujqUajMxgBQtdjNXXNwPU31NGBiZrziPhhpupdt
4f6mqCAjDBB2OBXylrh42ooj9ou8PdedZWBkzwsDVHBzci4Gc7u31a6tMChkSWjV
IiXJoQFtjTsu77q/IP5RooYnMXS3wmrWkSkwwk/OSBUAGU4o0s/9z/MX/y/iUyro
lCuDejDUY7O5OAuIaZzG7NycFhgJXayfZoVVdIRYz2G0mfEMF3r43icKzB3t4xza
NNt+ilcwircNfO1ODW7mhcHTuCQ98dMFrb6og6v3ZfrFZtasxYy8CN7QOz7e9FrV
H03wEYc1kOgRSNDJwTKdyW2YHhokCADD3hHpPowP+NbJLRiPLTBzHaUJFI0YVKVc
szopEy+L1OrWFWA4UtX4N8qDM/Il/IJCCVAv0qptzyGFxnKd76jpdzab1agiNVyL
jM/GC+dI+1iZvo7KjAIKGFIhjTxMG2TwPlnrrz83Owc+TG1kyEGOLkjmhMvumst4
Eh19QzMidG9vjJ3aDJldSmZ2+QjL4HdL6nxM/uBj5uw4xk7GMvo53WbmYoZTHc2T
1j4bbWxBm4t10IapkFTdLqMfH5Qmb1DbnrXS4LztzmqIf40cybEtk2cHsWBk9eZP
SjebXgBdKOHrdjlOGptscv1FsrcVqS9c0qtPRd9hazcbCSGe0nuSV0RZ3YVfQ4WU
SE2C3LIq/7WQkLJVVOVYAXOYYYk2TxyZAgrCG1PVkUtG23iJl/XwccptAn9/O4KM
IOcFCh5rfnEUrj86VpFTlZA1mXv+PO8fdLI6Vn+0xC6e6Kko49DGmW+neSSjteNT
lsxkUh1G/hqlpNR8hh+KUjY0JYDri8FUeJWKCe7bR1QNO2hxXW4L39v7Z8EQ+//c
4tOlrDgGodFW9xQQyHL+c1hAjh7bJjim0p9b8RuiRikHjWkV15hkI+P8M1J6G3tR
lbwVV3idS5ZxnIaGK9TIjVr7I6h7Ne4BV1tuk+EPGjpZEnrArBBCYdsDGkjKejez
1shVIKErzOPcv0B8D1QSeLybLEROV8nEkGNDQQ1ciLAYsZgTdT4A1MADxowd/NZc
4QQPRAmG+TXcFoyPr7TrlnYC2ZUZdUs84+TS0+WCW08QRhYGrCTHskXLYRBRUtdg
Szy4HAjxIWR7LWT4BFKPODM23zyu3iKWtLNDZNW8TncnKBQCWPe24/i+GE0Wfk+0
HFz+nLU4kRIJPlqZBRwzlvnKJc9DXcC+fIOtuv1RZkbVSJgzRDHf6OJnUJZxUbZD
IGBtbT/qJj2mGXBD+ljQcc73dre4LIbqWvQGKOaBABvcGO48jEjkcksysZR7V8vf
6jds7Yc9OVKZNDtO3DfPmZXx83w8/cdUsBdoZrwZc7OZMUW06aHVYHZFtp/WcJQD
0XN7cKD0aUlyObCYWBqT1hA6HlssNgfj6vPEeaiT8sKIoqub0/tEZFATjcya/St6
zDQwzLS+oMYZf3qY2yP9bG3xyNDpXzZ7h4XMqqseKjtAl2LDJhuT2or92eYTmuj+
TxidtUzoRnJ4Y/Tbaud6rfhLVqfE1KOn6kjnQ6kTmlbHclcs0SDfo2UZbZiywzl8
IxHy9I6aTh3HPTcylliT8A2pkxybU2r8lft4CsWN8xCeRO64dPSg75ztw8CuE6iE
JPXUqz6yV/frB+bTjcyxC6rtUif/PQ7AgitjfWwI1ZA+F8a3hdwF4jxM4OZqkh3o
VWLXNtbkzYackHxvTE0vbGZgErNx02bsYEytQS0WtL+Eo8U2HK8F0tKEhfxHbG47
Kx+bp+O9o7UbboUxZKSdT/NUo/auelatHZb4V9oNgIPsQuQQPQQ+BicaxPej+21d
DWm2pOIxOLoCW27Cwigg4/hWRXTf0eESqmVHz5gWDfDWeKgzBfAiOBmAEjJ4FVNQ
atvVAgCTJDp5JRXHF6bR9y3peQkuxJK/UgJ0wvCmEb1gnZ+5uKPrAIDoLsHvU/lV
u4FpNYDK8hSlTElsU/vkuxF57qTUOZcAyzXP+9PCmr9waLi1NoN2bFf9yoyrUKtW
mu/tY9EQ1DY1omJp3/+TNZIjW6AmSd625YcD/f9y5mVDtYUTBeMfz5/WpUqnsiV7
3uz+NSupOYIs6Xgunt5bNv7FN2XLEed2cO+9QbZyRVUmXYAOztfu8n9pyNFDRPDS
7pKHuPpVR/2fAcBzivFUYXbyGyngxCkVwA64Kf9YC9d9aL+VyP6YsqzCh83s2sZr
PIVMONdhcdgGI4dtKaWF8xhQRMmTyOoHjrmZ8imxlSOkfqQTbcY3eEmEOMEHT1wg
NhFN20Ina/nFfU/v8goFjzAtBpq1/cL+3G9wrp7RkgqWaAJIkSgItbQydAnnnmJ0
r7IZWu84xJiTdzvWtkFXqebIGvOHaM86DUHb6unRpUec15cZ5I5VGmlKLCHvRLcu
IfEH65li1lLJAk6nUfzW5m8ucoN21Fo9F4PYwVFMFKo31KzgrmJSjgxSCL99w64L
zzjHP9mdXeEqvb5s8U+2LomDAcLRTnupsZHuDSkVmerjIQFVVVrl688MB8ft8RLG
5IyVEDcrLWUm/gt1ejpHJJafbX+E7Y2VJYXTTAR6yn79UdiloNB8ZbUceYTdOSRQ
yd2e/MsqArPKuVdCdraQ6WBEdfh5hPiF5qteGShFgCp16uWsrQ2NSY1TLgd1Lx1C
M3qOPNmycULNepKXnO/HeLtjwMa8LkFz1LldcDGdhyoEyX8AR/AM5Kr7dp6ZKzch
CkHQaoFZGxCn6O+p6gmpl+G7HhqG/AbF902zt3r2sOInwtFEm2L/GcpvIG+g8YE/
fqyj9aIPPxBfPPKllxWOAxv5MtfwtNYXzJPlDuNzxJfA/SnD1AaxQ86m1fuVodFe
nYfkRJ9JRoC77JoDwRCK9LKxz7rQJsBt1zlhQF8W4v1RHjv3dLHTvgFQyGivu45X
b491wgwz14GS+7jbsbDwCSPj3mpTkez76yt9qEKorO4uQxYxtpLpo5E/H13Wi4VE
1ieQC/ol0dby+r+2PC01SfpMp9QB+OeYTOvHZlrXF4dJqoieGD4mkMxzB04ip3F2
8x9WwI6eko2V4TPA/5VJQZg5i4T5ppU//RUTqx9WeWz7409V51hvCT3yfnnIZUhn
gChkzNCid9H/m/WgYYpDB1cR8vPmlOAgNdixAqhOI+mKcNc8N+AkEvKVnq9Fb1xh
jyan01bOSBHkO4nDETAbi3YHa/7gHrlhqfNEwnZK2gOQpI0sOnxMY2pcNPyH9xQa
/EktExnRMHIC+LVqaYceL2afo0XbNFCgbqbg6HeIy+tNnECEl4vTXPQtAdH/Oo84
aIv/vPTcsX+4ewhAQgSsoJ4WLv6ApcW564iCqnwygc5J/kNF7hwB/ann7sGZnPX0
hWgUmBaZMyJjYbnewb7kzFtjgMKDK6VtGdvqy38RwQE9MyqMx+SvlzUxqCfcpA2w
aSAw3hklJtmKiYICaMWkFZnwaZAjoWWpHUD6v8bWBVvQf5NFq4ubU5Cu4HDNlyKf
o//4x2zJSORC1rWhirbbo1E2zQiczjcPtNqikgzm31baYEDbtJ8ZYzDIQtH3YkuT
ROyE/870uWdnuQVg4NUoc1cK9VyHUTnDt+JtTpWoQM43C6wWh7kyBM5hxvPFofmM
YTpVbNg2tkzHo6n4Tzib9ps06E/XJ7Lui3UIyitqZL7t8qI1jFttVmJBDQME//Aj
Qj/GlcwHO25YzgXZhUPN4aL7wchekc6nkOQSlTfy0j8/BrprEil9k6PykavoxiPm
rnIGHsvKafVt/lZG+37gla9Ze4LwSZCfWZIQb3MJAK6Gl9isAbElpqjiwOkX8cab
F+RQAqQmHPP/06GHG2AH3s2+oJeXM71tknhNALFsvEe60jbj4nfv6DV+pg6ugNFk
uCJch6vECaN4d751QtFJpjqLOD9pLI3fuEAufyLlNUPXSSGXDdrt3DRaamybxjZO
eNAWap1h1kfRL8lGPp+jT6lAWUoAberZV8IQyK2vHLHLOygVPS0aicNYL8X+30Ko
gVP988FqosuELXgsu8sBovkvRgY6JNc9x31dyw/0AfhOdTq8cR8yAZazPFrfE0IL
sRTEZK/aGLy7odTK+wvsbogmbq4y6GmdH2AXA0EspTETexcxZrD38RDqrXoRIhV0
uUHVRRauyunamN0dASPGwU9DP5ZkhhN7veCFO2klAsDahbXmNie1omGk9racQU4E
4bt0YVCzjvGtfJuHLH9uIE30L3sJk7i2yb6HOJGSd1MZZjadEwElS5nLwdeWal1y
DoGKDT2tN9O7nvlvzUNvY/cilSJeofMeYNtq/pGeWcN2lO37fXKYwzieBgrwDLDp
zNlAlp/VPIsk40tAOwxzi5XQQP3pvSn40IsMg2IZwnBb2KtBeH+1rhWHbLbm3SxN
opBD2csQVtgEp0fzmjByw0XJUGDj+IY7sotDMm9EENVDoF0xJcpyGRH1zgDtmScL
+kodHufIQB89Dd5kt4oqPyKhZySz4tc5v92U9P8b/uLVtYYOWmQXvZFvHSxBn021
ElV6cSKSWXLn9nzht5Unx04DPb3j3mnD2xHAwQJamdiQa2z5Rwxj9nR/8jIYMXJ0
vR0tYPx+w5ZcjYNnWjvAKnq6gTziSLdnQhQVgJyp48z/GKGLjQI0kwDhwCyMJJth
dmMJZkonE7h6pBrijraLygkQDlnzMEhgJEVkfRGkPta1yU68ZfOigNVtHrqvLRdm
Cu284k6kD+/qu9iScD6Vqs6ECr7rb8SemtH7Z/eZvGyZBCajtB2CWfKs9s0dKs29
xGIDi+HOhEJKhMywXss3BRIlCJ72KZhqdHp/xXTFqa/EvyOd6rIi9ShQYLDzrByY
tX8m2XmJbd0A5eXkDpUcwaSgGj1vfGVA0ez4UTZPQK6N2VsyEomK8sB9f96qffaT
x/Kg2FCV73mrjbL8Oh2SfJxvr4siruw3VTtJJlg7kAq2KldW+DiPdC00R7y3JBa5
hWj6tR2hhSwIMcfCWhvdhbhEtCXV4XUkaGkZji7J+wv6tvhoRpYqdf075+NdcCtl
wpklii1N6KsavUXI3hOGJXOso0UotPHDwGvxz0wEFmAc9mB7BQIyiC/oD/Y4QV9x
Z1i8YuKiNYMUE8VZrtM7bluy+X1poymzCV3RPdd2HywGMLV9XBVmHhOWzfuM6/wq
btvXE2phgTc2TJk6y4BLVQJ7yABqZyzWJCbPa7s4wu5ASIkUsfWGf/1wwv1qE7xx
moFs2dwHLk1J2jCg6IIoA9quf+DcFInuKF2czyoCmgLx0iRu7sxoymbfWtbXVMUh
5r77e7x2z4s4W8tsjoTxO2GUrKJW5PUcPfmZSO6pMb0q5U5/xqX4oKTmEomaf248
B3s8w8dIcGVcyiEF/j9MLD4RGOblgJO/zMaBmkvVcHGM+6ClIQpyDoO9be71Y+VB
IT2itl2q895mNa3/ah/owcGYnJNz7IJ5iObszSiJkPRgGhsjwGAMmqUvxRhFb812
JAneRNgnV/abO4pgdc50OoC1TS2jw6TfFGl5ISJcDC9EvUJ9NBFHDSWfjbEotZYM
gv14OWsZ6kqWP3tz7KlGG4zmHA16V/88JoqEjkexVBgtK4c+fghiUAhsBM++dzoM
FBCr6NOpngS/0aFRrqgCpyNqnMn9tZNWqrnb79F/Bek358l3z3OUJD/5h84+Mpd2
zN+jTLHbjs98ULoGorP8ZNi0io+OcCIFV07t/ni1wq0cQGoI4SP0GfPZlm2/e8k/
OoC74Qc0b0LHpzZxcuhzqAXvoU6xvjL6IaeMoJ5gS1hTma6fgOPO5tjohVY5XvYm
li8SAOGeNWb0sO0Alup60luV/EzqwiHnENbwDJ0iOas+8N/on8wse0EkAzAKMMA9
rS7yZegn+bX6S2uN0e7Y1Cvr+2PMHNFR6b2xgr5b6EhX85D5jqWv9dgm8UpZEnKU
pIaX9Fe7zRx9DETj8M7Fs7yQxCu5HF1/9gu/RA413db6ljoZEo1oxEbBh0WeVrBF
uWbfz/s7USsqg4JjJNYTM36aOcQzxlq+5AdU35tOtnuNapLAxiUBpf1ffV7rutuP
gN7Jpf8b+0QQB1Vql2jHNpC75Cw/r43ea4May81yUefV2/ytNrO3wXvcKkufWNRD
az5Oufm/kTATxwdgdKXRBvfSkt7wftxi/F9KGYCf3r9TdeH84vq4Xf12g3M5kV1l
ZZ42mrBT/OnbU+7na3IGyxfzLdlqjY72vmyWGNPbBW70RalyNzxZlEt/lJ0y9519
Xd1QPpyefeObzq8recwLrIIQ6YzwTgIGamOM7DwAqX/GuFUPI2J8DGZ78RHjaOXU
Gz40apRnT2hgAbTWDS1mjPVhMwS+pcqDi6cQamAXvKQXA7/1DXCvP39BOh0dzCh0
swSLKYyA0rl0enKUCNPSeCe3U/DkCTGWeJXm1Okq9ZFcNhFbyxpicCqECwfCMo3H
YArivcEKmwMt5e1n2IGF4dvCaXM6FpPoslIlW+7RgHZ3hDfIxsnudRAarFRyudl2
UiNpa/L3yzZi0AYYH1VJa58U+8wPGg1x4JR2a05EsKSQy3lZaytMbdVO+Nr+gcP/
csaBKhTW59oL2RgBgRlGLUD9luo/ie6Ea6JOVsEghGdjSkuwRLpZbohh6+WSYg1d
ggqHIMTTifqcxhvgB9FrWi+87jSxU1AzX7JINngOSGufaH8trjYERqlXmOew/gdd
zG3xAr2vec5eHZK4ZWY5X/gi2WhnoXUUbVnm7v9968oX/2xEef5G1s8JEhG6t/47
baQSmMFrrrWBH8eBjXeas715X1YSv8Lcm8E+saCdvFvZe7MEKTBhNRksQruusBtz
Zwlq+UlYd0Di0J3PDCAAITNl3lhGUAyx4o1rEr2+G/UWNhEcYmSe6wRKTuWnb9X+
K0uACWJDLGwVuF7sX0ENyLx5U4fHn+vm1/HIJ3kOuay3+pKXSRl2CX3AjrkGWTR8
8ckOHCpKzvfd85nej0/kBm2VlYvoOph81Br0XRobLkn0auZap0t6vyxKYiHnc+TH
6spYO9lmP8O5iBGZRev8M8VjVR81uek1Q6Z1y1nUEvmKIlpXs96q1Zv/EAHpDLVC
yZrgR12zcA95CqfwkaL44nbcozg+389etcVJ2cSPZoL/mWgc3LU5oW/W+8b1l1ao
hSE/Je1tmtXp0P8ivdsVtQVtw9ElPkWvJLaYHbczKKCZ6nVbAE5BQ9YOqOf0YTDn
x1nJ3SBKI9m2X5bCcM67xdxqoQdYqkaB0MoOwRUQAlB2Hrhh1Jn/uchRidv1/P7m
bt6lIF76VmAN3QL2belW7UUP9CC9J0BJgl75sNmDwuQX+fCsE6pa9gJusmbJg8Xg
XGYE+ZXg1jhqLPz8fVQfQcvFPWPivWnxR08VQxI/zARavgZAlPLrMdKttSDA55l/
cibOSPclrn2G1U13mUFPlaaxrSPj+RZcqyfZMlRWHYA2bZVMQceTky0mKAFd2JoR
GY1WFSX8QKZyrAMJAUBazc3b7+9WapWRA5ojsCvUbPW+e7Ev1foWci3SdJ5sGvCQ
sS2ItAfDGxeCyt7nA4hrUn5U/qtTQGBX4X90GkHrS3OfC1OdkmomntLBoPA+d70C
LSgb8bMAmp3+oeWjr3pv9bj6Qexl4gc5Zxk65pk0fAQLFkUFNBwBrXn0VBwZcvs0
ylO0nacQUUjTbnj4+YW5bNN27x2YhjUxk/6yK6HspfWaJH82CTci9lhwrXnzaotU
MspaCGpqzQfJwPK6d9DW9FgQx8qgV2YZ3qrhx+Kt1kWKRJy2j5lZH46kDloyysIs
WKI+U9aY4OV9xKvqOpU0whi9psNQe6avAL3TeH6MGZn42YheS9C8p/ApR4IDYHdq
I+P11buWQjVsHLJ6iBSwibh7PL61D+mQdcsdxq0K2ockaB5oNOoQeHH2C+50Qs1x
KIfeN9SFHOYs2saY8F00kK4GW43d70P5LIj6/8dyhdcnXaKrqdTHE3su/up4pD4g
K0endBXZAvyyPAfXdosW48mxrt0JBaVZFVbhW0U23OX7dsz4qrXEzJgDhPnxzShA
hXh7PCXZRwcd6VhqdrY5TMp36eKhXWeZHFWs1ALOzDPLEv08m2KuZor576NwmiGk
G7xki+MaVNvJEI05ofr3GtwF/8CL7jRAWm+8DSuu+4Zb8etDc1dRG1O8iKjo/MAj
tKJr/yrASGHNBTybJIpbMpFjjekm9VHAAxMyY+SOrtO5vokP/rITbrZuaINbU0wt
YsUlnICTd74cGiCvbvEil/wJ1+Vpvv/aObOJg8BMILSZtw7H40XUYjAsglSekI9y
uOYppbl5WWtJugY2iPCBUsTMSEB7hjWH1HL6bw0qKIY5KRMwgdTKakdHe3EACnr1
bRIOgIPkRatUGvgQyJa3IYe2wRaRDogUiN0hlqNmgWBi6qNqGuOJqzEt8e58Y8yx
EBfyNCuSSSzEstk7CgLKrgIz2w7cGMR7EVbZ8Zm89dYfq32sAsNLpWyaie4WAgNq
VBNV04+E6vYLxoHqrCV7RLqlkBueQpukdG1ch8tlPUBUaW4yz4knlZ/gvYUUjgBU
5l/2pdrz8g074F32rLnGMGNPIFEr1gc7QsY5a5SzmaM74QKNS3rsJF2GkEIRH0hR
iKXSD3CwdZUQxNflbkg2ZGmmIL+XSj/7JZWhWeUu1nAg7CXCs//bDe4rA0KrWm2D
o/tP7UK7ffx5N2RdCwzxHrcycOJwuHpDvRb7p+PF61pRoIv7nWv20G7ycTFADlIx
9SG5wdJ0/yFV0Vi69CUOaljTyvtYI36AmT2t9oFsX7DK+rYUh5xKW2ykTSFzBE3I
jQW+RnRYPCFE/O+lTTi1cC/tr0VoXB0kleUw7smenrn2guKGDdyHc5g0yglqAviq
dHcifc8QStaHnajdl1Ml5fZoUs4wrRABWCD4xb1SSezJ12D0AprIfarcsBOnFSJb
vtELVSZrAjoZDNWki66/KJxP+WQOi5VtYCgdTC954bdWMh8Zk0dD9hqreTcHpS15
q1REZ6tdrX+6at+b/udPmKWLkEh8n/W0tDzaG1+hvHjYEGZPHfE6C+2fIbDSx8+2
10iyrulFh1eNQ5dPs5abddRd8EHWaBd/o8+Qi3o3c+x/PWhQ6wlOTf7ehwM/1X5C
byeneODi70kdFuvHFt10T36dveGjr6GesKNDPECRpUuHOoYgMb3+CiBYgLc3+1LZ
ZwMjXBnDoSjmpfyhkTPf16Nm5syrJFuMAfUn7s14bEoYlEyszHlM9R/PZoJ7P3wy
obZJVxuW2Xpdw3KA2woC+4S3ZmiIYG3iQI7aiQAmgnNs+Yb+0jYhoIAfH5Pqal0T
3ztskXkSc9dvFFAyr/ScgVz3oVHlHh5kV+ilCD4gGrb9qmkh6qJJfpHeTg0BSYZU
rmIHSMRP+c1rsZlWh8UXuJKHgyFSHW8TaaDrANve7aJdXSiLEQwuZBiiS49IMWew
iwAEfqHUhRSlkSkNv9lcYxpA47WHUqeG9QRBCpgh6s2IZy6ukssjCx5rcFw9UfG8
MHBQAxB6U2E2XqJxKWMJN3kV1cwS9siHutkADfP3wu20WAbgmNVJkgGacCrIjDSM
pV4agNIHlxvKDLPZnKD86JG+xdnf4ZHLaafkroSBE2xnFFY49Y7L1lvLSY2+bJ9t
HY04Gfnlw1TswveIlTYJPrSl1GRte4wmaOL7kmAbv6dUmHhHsHZPGSd08qwS2LNP
LfNQXc7/Whsoar9vZ0ewFHZo0qIDD2aUf0VPnWSs4Dhc/k1tNS9ZwnohZWOtd923
+EIExtKtAq8kiD1dq25l6mkiDyOIb43RCfuMExrFhjdIbwa/4ri7L7ARH7UqS836
o1S2v1VZpim1QJ3I/WatNrpIZ5bjGlfl9gZnWRorVelLq2rx8LWAGoRwNYkcHA9N
tWIMCz9+G07bF/IuASMkaRZG3m0arkUarNMddFnfufi6TjB30X2eh7rZHwi/o7BO
1FU59syncQX4Yg0N1f/TTfxIEGNbSdl8NLS4X7oMjHkmBwS9i7vbTC0KEFAB4t9+
Zy2OVr42wFjGljfw4iwQoG74jPz5nMzHn8FKEVYT3UZIdX41jRsfLuGRntJuDJ4m
HSqDx0miT+ZjN+fK3KFG5jgfp5+Tz5snWSG0ckv33ZWOy3jyxxA6+eCg+2asGbba
GmIexEI1vh1Fft/Hr111R3DrqzIHHc7tMqIkLGsSHTwttlo7krx1Q3ROGI49r3qC
eGE87iy+57B5pvRhOcSh8aq2f0cFg2hCrNK1HTdeKD/hGz1hBp46ZpyIulT35EgU
MYcnghNZoVPwz09UFikVElfZ/1ub+Httz4I/R4XKxfxzaq0W9q0EQuHJmtCmI+Ht
nzU2F0hFAYx+C/z5Dp72gLKWQQfJRMGe4vbVCzgeIfNIUyDQpyiTY4IwjffAZcwI
QilE459tOMJMxOSoOdXsWHrjEaowkbEKRRhLZ+QWP+qiC3SqqxECLTvbHOluBiIN
ZxH2dzacPyomPgKrqdSSe6TmAjsK+UpHzF9ot1YLDSEezG6IKB7clYgfQRrTS+lv
F9p+H1YfnG9Hl1mzIqRmghHbHGCWIYk4IK0N2VbOfJ1iP8L2lS9XEATTb7t+ngM9
EY9adUcMMHrwHLkQC0kNZbFmS3aaLk3D1JegpGO6zRa1wx8NDmCmxzDPdUv6TxTD
0ustnAmpV+dVjzf3tC/+U/pWixyic9MvC0CNkKtsbydL57jKN0IRusbn2/KlpqXL
dNsWQR46oxcMVLvyfbv9aribnW+qaq/0+qwNkxiEJbz9p02neSoKywFhsyJ55V+Q
WHcp9Lj1wULQqvcyQruEOaLuDZEEnvA+9IPv+EpjkO6KqcYaAwRVPaiDKvzX0FMk
E3fCAcSCzZEFcQ1F3f9n2JPqpF6WVbJcl53QscQ12IMNWoOzu+PQh8VNeEiGyrDr
2Jz3FgEggQ/HsNSRqGQvC7j8S/FlbIsXY5MEHi48GqQ6GiDdC5ycTHHTHjCPBmS9
T6J/SwiybhKchFYcwe57IoDPm/Dil+aO0lHNX6FesFdtIdH4aR2SKg0FZ0dU83N9
sXovVQcaV2DphpSjwS4JlZmPyyS84rW1N7XWLpX2O/60YSNMWwwQS5WbLTyIlzhM
PbCOAJ03yWkbYk3BTXeztYZ/JeM95m9ziPHs4SHcOQGj4eYpRQ4XxyNLtrNiXqo1
zWQA3mwzr+vQ5m6t/KDnO3iIeQCBpHAKCf6v6mghgVfmrMaZcn1ZWFDHGKXKyXUB
sqG952X+WdmC8tsJx7JHn/2v8KYtIkjJNwVu/rKWw46tNugctHIq2R4VKHtEdxaA
aWvuYU5xa4mfqLH8VZFvIVHVmTrsgdva8wr+lmmZMGE+Mm2klanL/efiNWgRKBCK
sJfNGFwYtWRF70X2wAZaycH9kvWCWIyyUildJA1iij6IY73p+9YVuBhOKi4frqKP
18MAy/30YwufvE9rohFcpgCpSLtuADm1fK0EHyNgQE5MVyBCOvHUm0voecdsXjLk
l2868YhqcnP/lnCzZljX7wsIxuhoZsDAZ7mfm9F0QbrcJqx1Tw8h5ZMly71NzZ0i
wTDZ0H0K3AchiSsM9ZuM3cC+IJ5uITxvEB7mQTue3hu/QQdFmu9WjAjNmYE6eDL8
dSbIIs+R+Zj4twwdi7zm8zIpjQq2o0hH9GC6ot4fFnlwhTNY8+J4lkOMRdEQMe5U
uFyUcL4gOR+PKAW13IiHyHGqaJfaymUZtGwCnUGQJ5UQS79MRgz7oi8WgNs+Lux2
IWKbJFNUM1zaPGoAmuRgY+pVEm1oxLvqh9m1y86CtdyXvPmmeaME5En5BeyZ7ZQF
6LoF6ujbdQz9ZNYO6zYGKeOwbMDo2w4MXWvO/KWOinK0xf3bDXKQQvwxCZdQfVyg
P5GsH6KnTgbPtWdZVvMmanPChT6XKY/i9U+dNxvSf2iNLBRGNnHa709L0X6sQ/Kf
xrtCjKuWYPUt0VXWPLbXBwxgTfM7YF/043/hUzmPQOLSUWfY1xvlBouhuB1N6EvE
1djTkcYIDVs2MgQ28e0279/xN050PCTnNoAXOS3JD+gQs9OH7/G2OlokPHC31EkQ
fujXZ/SPRArVKFNoq6QYv9EhCDTSDfBC53JuHy3ljbT7vfOXMn5q+Iz8pKPz1AwM
sQfElhkiYF3I/Z2vs7b41Rv8Hp5cFDu1Ksk79rC7KJB1OZBO0pv5E+9u6ZMlxymW
OMovw8/DJ5TLKc5oyRhAWnyhlf/Anjd4pOTHxde0FS6AJmF7uEcyTKrcKWjmr/4/
jnobZKWArCi7BzpleacaPEno0nUolxDfrKALTCHu6AZ2zt6OeqDXg5DesPsnFfn1
25WZ2VF3XYKhEvrN2j4pXSEzcnoBPYG/hi7UpLexLa8xF3TxeL9K6m9nCilLyGx3
1FMMFh5Ip0axxCKx665KYxvPnjGlPMbWR1S0Vd0L/LyvHfboxYoE5ZpORx9OglK7
k8BFmgV7YrsTs7/viBNDO+ZA6BTLqnGu7E4sB2ucQOnxV2AMuvabb+ekQW/Q0KZa
eJDWSrVDUy0Ytfsnycnew6RIQbjUE6tZceG+IH/yWgjjTXBot+4crzPshHXecJsU
APLa+MrQa9XZvOMAxH1ejldvBUXhFT63/E5csCRoTx/MkuDWVcmRANLjvOKIEEHe
pIwRLlw4iPzpJkJae36db9Z1hI1Tgj7womoavZvpem0Ttd03JFVh0so0iTMkYu8A
bmAm96C9yjIsAkY6Tu1AWsPrhTqJO7AnplujIg40HBRu0BM2/4vXGh8l10YMqvoT
lu/7RuuSllngKkU7PO6eWKpt3AL/MZxEnLT4JXQ2chChXii4RzrJGpvY/ChUzjGG
ifrStuzvU6bDVzknZEmLob6GIfG4nT4Xe47x8E2zpNRQV+OxvI5vn9KGbA4k9EBt
Fy80Zut03UceJfQLCoYr49kXOk174qkZdY7qep2yGmpBhkOCDULfyEniwEeXaEYj
GmgYowh68q4C0pTDMolzrzJg0LefZKLqlflfs39N3u1KUTRl0GeOMmuIbR1ADKrt
1XI50r/9ZGsbhN/Stcn4w7ohaXGswl033lDGGcfVhq4In21z4E+UvL1K6kZyAwPM
uq/e5G4/yAV58wVYrRNiwXqa8/zPqvolu6grLiWqArg8v+QofiURZFK1WIt7G9ar
YF+MouuFIX1iKl8KbLZh2eOJohWVYlOqoEhe3je3p6J/ftk2OBHPi4wJqm9OkrtK
9QyffmnI4bKCVcIuUiizG3/k27csY7cIJKLplUeZ0IeydYw9olFEjUDHg66G02M4
1tT58ZiautOt2Fju4f1fikWQ2NWEvc6iiC8/etyZb92IUWFO77VkMlM0Y+3rMSiJ
xmXIPwFoooolQzWuBXSoLuAMSGZld45gmhZytLCDAyk2zmRYr+Fnb+cDJs6NU75H
LWk9ur4nf0c92EM2lvdaysWB4WdeAd3YZPRSl2Le7BFBUbNejhkmsSb4C8Dnmsbz
jkCPhgy7ZsBmz3IZYiY7sOL7mKTyWKHuEvlitEaSPgp7SIiz3z2+KB0UHNm889Ne
VebFwtZ8HhJsSyDM7aEnRpze4q/HdM/eDoLBVo08eQJehTy6qhN9KkONjUCr1qbi
Jxn0TdCXB1tQMZYMIbVBfdnIzjUw+dhVtcfffEj+JwbQlnrinAliV+MEnJ5kUE7s
20K3akYZI1k2N/7y/jMmfQwAcAqIPJ9ufh91IgDogKXv75uoX11qc2KzH8nLdG/a
s4J1SiZN/AY9UiqgtQGT7LEFAzj22G9LYQpFwpKp2j0MOc5MVCHLn3YP8mlWcjY0
vmAf4qJ+9lFYvxnN1NYyuEs9dHIAsBPxrAiMccAsAlnYOdDQu/VWRepp0vSVin3n
MsNWzq0jNwQ0Ez3pD6Yk08kMLJ7g2gOaNjIIoLzL/nFGTNJVsyOKgie7CClzB3f3
RWidp6uKYvl/0Vu9XFFDmKR2ANAfywjjfWTioiuOqBr3kVpHI9fhwFebSECEUoy/
BV9z3FHtwdzGhlkKrfzMYDhOldxDPteR6pZuNLqsE9X6DWhrXq2erbRYuD1ixyCn
tyG3NsC3z+RTmyk/bEBL01i2ACwQzlwcHCLkCOFXVRm2JOplzHlocerEPi7XLyM5
fHsavkzk2oT7saRjjrvBSElOGadErsGne+Z84wjnFM6gCGxSzJLUalAVkEUap/se
c3xITFNCqklpIqTiMYRCWjD5alV0xiOuvmWHbECyjSl/noabnitId/J+kKw9FxFC
VGpxv9QQwbGw/Us3bN954DY2diEY1EgmcXMBd8PW0DJt+ocaTHHXttaCXA9fYzAm
ais4MLv2IZ2x3TB8JEY2zPs+wdbYrZEb7ceEIYsA17CYzI/5XgcjvWxas0WYUpNK
POoasScXdYx1G7Um6whKUcvpyq1KkUfRiRbzFgr5JX63Lsz3j0CsYaXJ+HXhXH0T
Ra5NvHF+BtYdRMflRDVYmhDX9ucgbGGDETd3y3O5A1wMYwR0mtW97rWZbsD2nZSS
tnYrI/V2cdSQwKcPvWh+j+Vb46yAK79noXcT9CrsPkDiUeIr8Eb2SiG0B1y8VKZL
9YayCBFQrn7R4h8heZTAaKTfIu/YVBIaa/CAaTu6flXYz52NQODB4Ux//EpZ1qJr
AjVdfrnFZD9H4hZnvpvDrLPEclcdzS4RiGgU56ClsJimbhYaeHBMkHOQDhvfhVvM
XPNxoD5MHh+jCYR1TGm7G7LSP67y7NholBBdVzvO2Xy3Zzz/oQz+RScOMKupgRrM
L+k3zKvRsMf2s34dvlCKwFLTTysYrIhMo5K6czgcq2f7KloMI/N/vtvUs1SB7Gq8
BKglX+AgS4DaWzB6Ht2M2AiRhl3kjFF7oM/FR4iLU6RhmH2B4/YZ2I/WF4gCuSvb
MjtjVnT7zvvk8JuSOuAjJGeMSdcMEZOyKpXF35QRz3jwQomZibtASGs2Uk3FtJNi
BAsF9+8HA7gdGXL5rMO2oHLaOKNZujE3y2Z67gWOTjaWVEKUGun7DGkvTcr+BPY3
efZTSmZMba5zDgtnHwvqgDn6AFZpQNaCROvzQZYtRIRpXqb4GpIVun++RDgfYOaP
FyslB9YbY9DwvEGjbI6RJc68EMvWjx8JjwwNq9HGZXwstYZBFfCB/fMTVzqatzEF
k1nHlrVaTEHauoO4jbt2OYe7lrmHJkyGqgeXbbRJ3jc/kPLuVy3frH1yaieBQ5PP
g4hMYYHA43M8e3WFmEvBW5mbim74CI1bQP9V59sFtUIw9TmTyFAqZwUOyVb+N4wV
ECT3A9ZHkMtXln6NJ3g5wUAupCtDcYB6SCiXOkhoezfQoIbBPBp7D/NCywKBHTAD
t9AXOr2gnt8hZpRQsNuV2ipVRPFvOP6YD+ZSE/m49t7JkANv2tKKrJXCzUhbiqxU
zDjT5TRE9HfWVdv3YUgeq9J/6m2fUtHfPZ/Zu/mM0mFSfW6/AfqRnRdFNvJEpzxa
fwbSwbPjW9dZif7yeg7jYEfThHLzzyVcs4ldGhF5rDXo7OZJg8rUI2i/8icEv4k4
hszr0OJ41B+SaJQ5iBA554nq2G2kOzJH4vWIF9cGobX15B46IxUhCbP/N+apikod
9HPzMiqhNBjxeympRV26FA2UCn7/3Et4KbU1xtFiyiuAiCyk76x6174fEb70Tfn3
/pCqARHq+fXJWSGOMOtf9JBYt/43rVh3BBxoF+tXZkwEIgtMH1PnHqHGuGlxgk02
IpeIS5XPq/0rPqAxg7O/gVvEjcBSBUYPfjihWog9MrCgyLzraqEiphpAKnCea0W0
uJzxuWbyj7D5uo3TfAgxgqgB7HwPcbfKFGlNtCEmGww19vL++lCUQZRvNRLkkiDa
4yPrK5jOx2ekMB4BzTTb9c4Ql4kxxa1ntBG9L8nmasTN8olcnKSfFDUgH2c3nzpx
uO5vJnJ5U09hnewHRSO1FOKw1aylGKMpodQksh5Bzu/NKxc0O8s5VFnAVZjwHkXm
GtM4CNqMSlSUQeso5mhIcBjbg3IMd79DMmfOVzOIgEP77Ckp+goxiwF3bIFib5s2
0kD3DanR909B/n3UmWV+sXuRy6NEgIYUD7OebGeKuq5DaIa9sgXNnpWroEXPDHPK
npvY3q6DgsBqQhDh/kDSeEvsS7hCE7QSik3j9elw7zwQgi/vMqySZDhLdMG+/llZ
ouZZxFmtDbFIRpv650ZAAlJStBeJjOoHs7/PxGaNoA8fmPzOX2Tj/Fo6PYmv4l1I
TL+IcaQGJcYJD1K7M8LyOnxlu5O5pZg2thCfA732PRUGMWvkhZCeEJp3eW0F3cbM
BFaNo3k8W1HwBC6vdZfoRklUxb7BYl8FB7oDRbtNjg+KHVJ24XWTCo3ZJbd0pb1U
3P3zxrO+Mg5xMmeELKH5/XVtCjHvHyHLFG8L/nRJXwpXA2BtfQgby9erdMjusNdX
whJYKDHdiE3Ty1WiN6Omwhh4y+jdaofvyHfbOVchuAn7W6Hr8ETbBDGtF4Yd9E46
rCiI1gukMIloyZqYUNBht2Lt1JvnrtLqbmiBnHOqWm+rwnjLN7IfwfhXWsEv3j40
hjqB7hABGfeIrmtf5rXAlAs0ZMKQoIFsYDgoGbcjpAc+zoBHTMokqD/EtericPI9
1v/yHcGn3AOPurDFO9IXzTgQIn/Px7/bVYuqkWf8ONjZodzoaj1Pcd6cTiZDfHRU
G02b5Hz3q/Vgcq8z1WArD5WyvJRpKn4D5+Pm54j+2g9uz+R5VrzVd1Q+UCzYg2R+
d6SIf7WoKjWdj2mgLUZAPnkhEHWF0EDKYDfO6NckK7u4dmjoNTwjubnyE2j5d/p2
wMS+1YI+ZpuMy3Ym83yYUgJMnYQQ3EBUjvlFm71C46m2QNxE0YvKZrWMEWmVNZ6O
qVyziyzhg1pjyMqeD7MSPcsDhsfW2jrLqxYB1BWkW+OGRqeK/uW7wCBEFPujOXH9
ii2OSRi7+RUv3NrhNjr0rIgo8c72dx33TN++Y5QL/BjDw26O/bvBSxeUYF5U4gWc
cvP1HAfUzgo2BzL7tD97LbWqkbE0qbL/DDe7CwbfXrc40Afa9za/s6p6FJ8OJxKQ
9tjaY5x7vc5ZVwrVQVu5PatP4GnfYULNzg5qeSFMPuKp0C09q3NzO3LvaKk325Gg
nSUxPTB4qD8O9kLxIQmpWGVbdnegfAtWOMPOLELY4RCg6vHdu//c7wU20XGFiAp7
sX2WaoSWrSEweLXQZ3N3sb/oobeQ7NTZQvxd9MwsCbUrq8MAtRJan/LR91KyJcHX
MehoLF1DtwSCuhT6yAvZBhT7j/kNOp/lucbbJXeU87LH/7yEM6abgWPSaSXwMCFf
4ZD4cRSoF5/3DC6F0b0Iog/pL/2xnTc2TnoHFdXCk+8adVr8TK4+aqH1Atpv/6pz
HXZ5b+qj7HS+PxsIGufgz5HPslcjZOwXUbPgnrG23vN9dCY8404bq6v7WoHvcPEb
9RqH1Xb84YtyUXaralT+lfm74PrlO9GoSIycGS5znsCojF+GIfAliAk5jaKv8Tc4
K2hcQt3aI8Ii9jgemABEwd7qqBoVk7Q9/m674PzPaLliaU1mPgfS5Yd7Q4aTabiY
xWIR0JsH0AWwPFsEP3Ljjst768ljXPpXpg893eRzLND7+AwDZB/cg9S3gE5vV/Ao
Y0zj6vA4H2INeFwjwkYgIGrNT15v3VQUc2r0wPFvkHtWoQCX1eQ99DupLsX6ntd0
nOKiu6PUAtbA7J4ZGv2BOtDmDI6X5O75F8x4/+q3gMzvnbYnpAsuyaU9cvnMRaCS
Ipdz9Fy5y4DnZAKFWFYmU45EMQOnpU0h5hKwZ6/xnkzlmhk0w5Rd6XAFQqVAFPav
7sc/Anq+Zhvr79fsJUtscgSl1TR3P3IEGs+rGXD6W5R/SVf34Ym4n5MdN6F9RYtP
b3NGfvdjxfpMvLcBEzuEtaAEoe6LDyNMRvbjdfhL24gfi6hHLp4mNITbLH5C8Sqw
EnPyIx580DFWjYRCLF4kjJaAOWqusHeQnPSkKnBDLjZYnlrS1GYlNBw2DtY8NDef
Bc/fKGQdVXkDGB0yY+NUOyIIEumjZwvWiL1gAlWmk6h+to7JoA1Q/7JeAOPOOi9z
0VKAArHI14BBe1zapNNrF3FiN6oU1mb0fvDeG0rmOravpPqVlJdKcpSTyAB3cOOJ
UF7GjltNuSh2OdV+fvk4taspHibXax0BGjhIuWYXiX2PcqBZ66InM4LvqHDMbDbY
xpt+TYxco/BuXhr3/ZVNsz36bVa6Qa3dOG9YOnONIPwxV8klXf7uwONn0XcDAe21
EObeTaavHNlvRxeRppUeDmSMiZLjjtivM4tyjf78k34wD7z465ZMfNnH5KkHTTQc
jQlcLzf965zVJBYASH18fN5LZKOQnVz2NQzdMZ5nijRVhuZiFlPHekEAINB2Iq+v
QN5BOPTDAn5QFnzWD0OSqXVQtW+g+SJud046HI3OZ/5dy5lygVrIviQPMW0s7z7V
ugXrP0tfrA/RiZMFjUCIpxlr9nw7jrzST2CR8ueIRWa+TgBmLyIiG/UQjUV1mhLV
0S7nzrDeGJy54+hL7jCm99NEpxEd/zFPfQT13zGfB124CDjh4FKs05VchiTFpEFP
G1l8xctBP0riVJuE60krCcY7/kV1sKv2Q1hHqXCzHmIZy6ZW18UI/vMNtbmN3mrG
xRbwNKVkKc6/JcRlYZSj2xJ2C7bfSbpUl5Ije4+i/qKx87WkYk7a/TW8l/SLL3k/
JFsnSwuSLBHvlwl5NcWO2O3ei/TGMy0Xw1czwv24uiyE+GdtAim8/5h9O9I8M1GP
ucygvHML3WeUNoep3LptXsgMSbjFsOAVeEVID2oOKbMm02I9JJru2fksbaheQeG+
9uLa1uj/eNlwVwUlfx9EMr2veus8yo15ODMhZd1zXMNAOmYVexFUIqpV+J2itO0r
vnAflFitfWde0MFylkNtl+gsynXm8PGs5/8Bia9Atcogw87LGG90QNv/p3AYxWY6
7jKJLvjvnp93dpHZLSxLP5HfShOIfLIBZfEoIxiO7BGHdqRYxxmGeuc58kpdWEtY
Zq6ZghP6HlE6FpRDLMOhvjLJjt1ySUwTbgR7o5KcSBsacIgDpqiE6KU5L03u+LVM
ZrNdZpE0btCAoDv+bhMg28c269xixUAH+r4/6fjstsA2GCWl6lvhT8YHt+0VtUFF
hCnTE3rIGyMwVORhDAGPbIZi//rtkH7CVX8gycSH6YccvovEFoIabpu3q30gDgE3
lCdmJSlVxyqj9v1GgHfL/iuLQ5H10x1xVq52d2Kmf20fr/XCGd91pLRQlV4av9S7
WCixihjtoPoNH9dxi00DrsrGZH8BxKXQ5qjVwLedHnNEBnIrDuwpiac0lzBSr4hG
zuo+k2nnLZmTKYj2W30bCp8zWd0Dw6AYwXZcjzwGGOOCOZbmofV3qDCqQqSXIF7S
PTVc+PQoBCMKBJhoj3tahQlNu+Ju+bYJpKIniyWaD7x89psQaeXRxcyQ4x6necFK
atU7QolDKqscTRvBbsWjH9nsUUE4yR8rUwmkDHOWS/iWffSfnKt4MASJ1vHEvtsH
/J5HR1SyYHl3V7xGOlxaDPsZ0LOiks6585384mLjWN0kyNjq2xb2ZZott3D8po8m
s/vlJRlNOS+h0lQS+oyi71zWoM4E8q1vf2Cvhv380skXqqtJljW1OaS5n1jItHa/
Gf6csstkcTj+zbAwchBlVJvg1kaLdgpuVFN3h+NIIWsUVRIqTQgr3uelXrLVBsft
Gt5kMTQcKA0aaeHr0YfyuiqWHbTmFB2UuSh3jtnkrstnKA9W+dFq1NrrqoyKs5xp
w350rsIczckHHZlAM2hcFj1Aafni2Zc0kNdoBXGQSlTQvFys8izYIRvQuHK0VN+b
BplGW1dSwFEpNphCsv2PNJwTREkPkwjTlvnkkZ4AGn5JLmWl/r9FvN7kTWJkSP22
lzHv0VvskYbTkJSwBC3J1pu5+2YMyBFldgSVc1F/XWje83Hc7hAjZdF2a6kWD0c8
jJjQBj+Jg3IsZBHUjinctI43PnNGNiUHn3pfRx1wAULRxqSksnnomorqxFC5FpGS
GaOQo9CJ2Jezi3M9Vbwghu6zOkDMoErA8+pDGmLGaZlEUw1156laEk9DciNspqLc
pAHCOXb7JPauz5BEJ0XYQqwA2vGJJWmx1Am8J1rsDDG8LoipcNc1GVrIDPZDMOFE
TN3/AV/yrWYlbnof2OKoTORdw252faSwNZ7R/I55nhw6fYiPizlf8PDVD1g8ZSJ0
Yffu1abXsNmSYdTnfjryeWPYmUA1G35RA1R0/0tKs6hJ9FaNTRxS9BsldULgLlvX
f0uJZzcApvhFhR8QSXlBapk7BtVyL45E1yxKMig/jVG2vM2AyISZU6XPOTeu3NX9
Uotgq2IonxTdlE6kRVeUqr8rIVm0rzJ3AcPQMKOdgbSYNmNUfya2iLOsYc6Z1i9s
Q6IIZAjeafhR4AKRw5/xbXMa/AE82J8ScOAerMrKwDWql+MgIi/b/gWJEyuY+u/J
yKsiKLdqy5P5mg8LLASd9Bqv8ewKgHM2hTA3u5wBIc9TYKjaOy5yEPRC4F4atGvI
3JZfh+TChS1JJrg4UCVFaL8E7r7k7CgZdjJMzyGVUnkkcwv0cj02P4wac/yW9AI+
7L05nfFA8BI0BoC0d6aTQktpQg75f0mGubZgJ+YE3kAi2mFZYHFLDz7Rbk56h56S
ZnnybKJGQ8fnvG57bGGF140GfKneDCEiybVNP7ALPXJxxHi9bJlq4GRK5YX1l9JY
tqxMr8HS/BbizjUoPgYR8ko/R1Wd1i6vgOA3yQ4BzLMVqZ8Zd7Dp6UsxyluU0v32
pzOOAUgImb6e3xSHHWeicYt+3yNYgumPM0NFQaQccBzYBFBPGVip9LgF60bm226V
/9CEosF6GebJRH1ALHWapkAH3EJwImzL+VngEdIKlnL8Hjn34RFbY0Z8OF6qUBDf
KpsVX8BbaAPQVpr+xIBK4kUDNz21FjYUks7bOtjZenMURlHiKz7H6l6p3JUZHVVy
RQ9a8Ip++8SL25E23ObcPPTAeK5z2fuyAlbqwIAUVgHXu8BGXHIkfqWVMPTdSZ2A
yoKBd4OUWyNzO/R26WnwmlM+FcEquDx9oimjaiq11i+06NAsKXIPABWVq0RiO/YU
KMNjMUVJmV29XPdQZZj4/5n2VbMeyun2RZ/4098YWvAx24Oy7VUqGl/CyT+pal/V
Hm+TMzwsKh7JSyk3d2LyqxoYc/ZMV66g2m3q9i6umiznL19g4w6B1RyAnp9ZkmeK
Bh4wknecDdzfsMaAyECO8jTu5hhWS8u/8ajdIF2aJVrnsGLbOh9mhvuKBgdMZ1kD
q0fPCcA1mQhjzYve0Uj5j8xX/XSjMna8BX8ENVDvKuIbx7Qn9TNYVRg7Ct3dAiHm
FBc8UsBbKqFOKNIVhDAJ2PvJfyEwPFBFLwVko2vjjl6H1kLu3+WsjU0zxo8FLnNu
fHOwLQM+Ve8NDATfQU/BJIwoEi1J4dGElDkEh72hYOYq14rPwbGIP6+eyPSvHktx
KNBIwUDDJXcUSH5flJ564sUcKfymnhus0GklUjyYuhCVQJd2DkcLO1sE3Ch+SMe8
P1Wp6hXLEr+VQT/WgWz2FTRrz+GOReZrTzPtW0tazIuYTzxY0cHQxANT2fbu0rrE
jlFdF3Wdpl3POiSE7GOMH1+fnpCJl+EPYoIBAw09RSDjJLmQITvgkEkg7O0YlOMt
/78tCeMtT9J545kLNYTpcNZKqO0NJAyizbqPWUJF+FkEgTmyvZX7btaPmtI+A18F
+As3yQa2Mj2F3a3OFSgtxWSYDpRWFSGZ+TK7p7JK++OLhDNjLUj6vnXdCECeUbP2
ZoH4xowwFo+FeMFglIi4lAEFl0bMWeWhb0Z38okMi2In95E0WAyfoSHmnghKccPr
CE0zWrTuMdVFmUwGwOcSgf1PvilgtzHlSU0ph2yuF15u81nLCgFPS63V9Q9pwwjZ
SIeiZ5oMH/CNB+WIjU6ial4EcUekVKG28B3OOBljo01xEPvi5QEI9Ug5PStp4QQ/
Wpx7tLCTDgLWmygu/Mn7i6qeDqbrAEASOo2iHLPyB7KlfxlEvjw5lXJk0OMHc/kl
tvJuPEnKIn6/HfhxS9yj8FUWtzase4xgyrmu4injnfAP0N6Sl0oS5FNg/Z2Z8rNY
g8uVIc81p4SvV6v3lo26Pv/3Hm+5iZ5Ak9iHM7iz8Lnur49RmZP9C3pjExOH4lUv
9TLR2Nc6jP/C2iOSRVOUUiD6/Ph0GRnS7JCWAEAFL9A+zAjAozt+hxxCSkMH+aCH
sMPyvXb2Whhj77klFUhJck6S3vEvn1TsWWW9CzFqs2AaDcIVT/8yshKu7JvV9VBV
H1VjrcWPleqa/Vk2ELNdG1X8NVJxTUZntYtJMNBF8Xa/iXrbmgeVADpzotagbvCO
y/ouY/cIj9MRI4EqI25ZKN2zpmUSw6ePbCnpQRscC7m53PWjvu2q14m2qrFeJIlp
od+/wXH4DXCRemkwkARD+kLKYOcapsvUtvza7Fzu4yKGsv0Xm2YaY90UU9WMlrL0
pZMIztaH4TVgXd65viTPXhW8RFYGcMo+twFTdw+yd5ya2pLYRgN0/B0tPSWsXfcE
38jY/SJKlHqRcEzLzNmPh4ZkbsvNmSxopQGkloa2kEzNMF7AbjezQ80v9BQt3toG
ztKa/3MgY9JyDVWbAWUgbxIYhwUA5ewJDgMnl3O3PBA7aMUJxO6KGVU5cwD44lx3
jlIE5noGb7WVmn4U2rezxzzRUXjNrKTezYoyv3DqnuvFCyvVek16Nxx1BuWEh9rQ
AzIYb1pzdCDIF90gQrWJExT+JpldOpdep6gRg0sp2aWBjP7PricZmY9fBA2CEHlB
/3ii1IoAz1IQ5FiaSPafgcBeXgxLr0uXp8Rue9GWY5OQxlOzSL+uoNdAzEP+8w6u
4/czsTDBcwRjq52z2c57BYyKMS1sjGAwl3y0fCaT3vWI1YzJVek6uLo6AblvyD4E
c5vO+6gIY3FhND031n6GkFAgoPFmeuTGl64x960d8pnU6BsPf75tGUskGGW+UZlX
shD/PpFs2Xap7CC6/xXVyuAU4xWlcw/5t9emSMW6W6+byMYg3mcxO6Ki0B5+zmXp
M8uL8lHGRKtHhx5ZNJTSn/KcpJI15h+UYPAZB1yhZ3/RTx5hp1lRvtJKdRNDVpX0
28vsX60c6COz/mCYA00HkC1Eg16gtHEivghERUZt0GWt/twhyKa7q4W3noQkVivq
WpfvESG3OiOMYfQDjewSJoKwa1VjuAdSTlrXQCnpKaO8MrUVJzT4Hc5RgUC1gs/O
lmhwVbT2LAhpyaHw4qj1i5bI+AOvzmRtUXrwo2Q8FpMwMz3yJP38Nwjf5qlX7A4G
8gIq4dflFilohLURuxKQcqtVCC+OoezUWnfSIE2rYubpjdr2noqdEdkVGnwgvNpX
qluJGnY6Mk2YfV13hOWAmJRpzOhWjvFbEEZjJZqVFmd2GCHF5tBeUY4ZYliPeR4o
wdJoM9MEiM/11F/QWQNZCTm8L+VxIH5+g/7lzkDYLxzCPeChyG2D7E/zgrh5aoEa
45bRnkNWlnAoioHRJVYAsI0wbZUh4i0vb/XZN1IN5Gwfr2klauUM26VGa/F+ByR/
xaAFkuTpIzKDFAWO7UKq291M7TS89MaUOWnRXc8BXFQhlgKnz76BpeLsg/I+RGlF
b3A8TQdwTfTr14CQbvvvtmfOdVl7cVXCeaNT4ncOxYqAaN/rC0HSciqLr5xY1GxI
YmWuYEY4jAklgcOGB2yHPEa9DM8Qbs//C7gUmmpsrgUENaAeRcnp5iS5KTfhYtNZ
f5mQIvEBDhuDxRsBjV6J6SH6XeSjzMMu5xzRKsyccXzzkVApOo47UJTT9gC2BfeK
3wxxcUvBczW+WVErpbJIvagwbDx60xz8DbjGzt9GgbreaaiaSWkToG7KxVaAlEoM
sbb5u5OiSCi91Xv4Uu0HbZuKugVSNBKoJGrb6bm3+IiFCNpDcNs4f5yRA/IVcOTI
twq80JZxNRd36Wf96vmg5lxBDwnsA17czmPhz7mdralt9dnQzsRVDXWJfIq6yZ0N
6bLLw4USC+rGRwbCZ8GZB82ty2FOuJ2FDeYQ0gUX+wunhlKex3ck5g8jm0B3W4W5
w2HaqH4eR/+00v1JfKjIjpqgrzRG8eL9weCg9TJuu0yyDlnMsQrOyVs22hODibNd
mwH95eJixkUQdnU+Z7nF+tTFAVeHpKkLJk+iiTkz1LFCGVDPDrACB/fdfZrLv5/T
P3ep8xbbxAzvOiBYrzhMmWvfYTZofLhh7Ic25dqGbLaAgKWhu+cHBGscZtpRpj68
DAb5LjeujeBjZX7K3x2D7u9BrDzrHYG1C/XtL4XgjeBqvIrpGWj7ttTAyEZhw/8G
NC+42pIT34ZBHSetpyy9c4zlhEyl3Ks1o9YJBAljcAAOzUYECscNgq8E9TsFTyFA
mPG17BYh9P3kCgdeIV4tkH5ZOuK67OqQPD5PbGw6gZcQdVPZt2T5KFrUPETqjUrf
kV03/z5Ue5n3QLG601bpfyPj9Buub9czhg9Fqt44wf8AzprCs3lzsfuOwijBU9vt
ZBdNPpnJWIeGkt5J5Jtyg+F9o8aUExzXIAsTcB5bS9MHJdxIptbA+oviD0Q5wLpY
4W07ZFjoLdV17mBh+lKz00srGxxU4d0J146Rbszz25YcDJ3Svmmy79mBhpgQ21DT
9pdipO8DjNPe4X5uGkHDKqD607BmBvXvdEYMo2nBWklD9RNxj8ePh/fM2eD7nbhT
TZhCK+5HT1I7OVxxmsFoLX7Cuxl5QGv5vBqq+9ubo+S2wV6xS31bJG7Pwyn8y8F0
Epr3n38LxL4yTe6O8pyXjBZqyMelDrqdbLDDt1Nohek7s7Y6z83yRKQV8XKdeV13
2aD1GIsIltLTth1J0xhtJViCx9DbLf7/tXNNB/Hf0bO+tcIZi+sPH2Kl6LPju5rN
+OsOSVXZ0V19JhZOZr8o+ndaEFjOCYNySsURoh+Zz/AVNI7e4yRr4lejDKYHxdbP
OTBe0igGNZtxthObWpeHkQ+4rByQESn+26CDQ/POkWlxl9FdiTqDLzrJMG33UwBk
49DwmTqi3BGjmc6+WslusBQxew5TVRxdz2FQ2VNpy58iaonZicBlOxssAhKodwoK
y0iujb1hCWpKLDWhmM3CGEm6IPrHCV2skZbb0as4Jsha5CyokpkYtfrr2JklBMlX
RgD6HA0bMRq09MH20FlothqTpQB0UPEUerJ56d+Kvj5nel0J8m84a20wseln+0FR
hytvN1vgD0FgOQ9X9th8SLz0XoL1TwnIMAcWCm1n/8tqGlDyG5NK3x9ju3QiEHeN
G7BS/eE4IJq37Cu5kCsQ3Pt6LG0cGf0OLD7RVh4myij5/ggmG7Zxs++F9zLp+pQT
eYUakDNgl7AtZe7nr9T6CHVlty4H3pimY4SE6pgHLzvxoUJ5sDP5bYuhuhFuqW6B
THDPqcYuM8aU/6LWLio/WmkAhwGen9IP9QrJ4hn5v36o8nvXI7VO6TAJHeXDPns6
ZicLGbsCJwmtjVaYmFIaz1iTwd/eybpqnQIPs20Yim1+d5UaEKSOSApTGghdfW12
izhrfrDbZkrHcNcp5GvMA2c2KzbIGgXMiv19nr8FR/Ez3FGmCF+wTMvMFFMO/arz
RhKPwSxtqgCoUAM8/lrgL8nJF+toX2zpFXLh7Jpd2Wo2cmck+e91CVv6BJaLBKF1
hm9TfUEpTbvWK7c6nZQ+qP184LL5y9vYkdHfijbjR2yKsX57l888TVg4qmXdarlH
PpgZsUV/JDPFlEfiMTFVGmPA590uxazzA2sZYNGMsMRRRxhnxy3UNujcJbmZIoKC
P7NUwhCaPR7+1OmbGbf7yS0CB/Ud381CN3MWoJz5tAY6YMO5QDIhC2zwfsHmpBDS
CAZ9UPItN9i7yRPAfCf5yBWJdTULWx27oC4PbjrFVI6NIGAULcT+yAY3lGJId7uY
WMdyQ1q865qjq4UOrqSSfQznErSph6SMatYu+lKvXETebTwVWYeCB9gfyG7fDG//
sWr8Zu0hKvhVyQZwQoA8ovgEPWJX0aDYeELGC7IKZ+R1sTCJlP9n8651xisI+lpL
kwUXOsOgkY0Ao1/buQ2LGkFYJg5V1Gb2zIBm0nMYHikCZtRK96O76EgkxdGi/A4U
LbeS2ki1ciPzHQxHRYLve5r7cvB7FCobHno/YhLEgN0MEViPaQo8E6yNQZpiYqIf
iJSBv0rZ4wkT4E/XrAlKtfOSaUtu2Yyk3IapikiX7QKoe8xkO2HKE3cuDxzhp4UZ
VlsWmMpVy5flR1yucvUQXmV7g1jSTibQyB5HXdQRqSxv9ntW/BHRDh9veWjOOP7A
0bhjKOoCEYSLy9A8H9ZyO0OhI1IisNoAiUaASgzX1BeJzrAs0MuF8WsmRsHdSFW6
RCW1ht2W/W/2WUBfxtXilfXviDCBc5kOMFkj7jn7BLPsoa0JTqZ4IaZzh9oErth5
BMYbmmW8VQJTya5W1lOhNcgiTmIcXyFJoOzexwxUP5nS5jXQi/xOGc1sY/FBE81j
QIXJ072iWp6lCCkMIvXBg53FNChoAq4CNlppWS0ZSbsWTVKabrdekjsMMKFP2G2j
MYludk9nCDpEm/s1Rj/qpvLYuaJzXiWYwj97Qwx9h+w96Zv5HoyJY6BUp0dK3RS5
a20mAT/vNNQfrA+Izs3Nh+i7QzfH+2RwJzD8SgMbtNkG23TSWwPAlAum+xRoy/Lr
e2K79cUTw5QHecZmq4rRgwGEn6oA3omqosymglKaE4A4S11FO9UbYYAUcbwOLMvJ
I+v0Okzcmkp8oNL4J7/BPIiclaxswquetZY+tgtPwRGwkaIzpEwSEtWEuQcHYAlq
0waIOv8j+d88YS74y4UAIfjK7z3Tohe5ot1GGCFGtmkML/nUD95mCjL6QL170mZ7
oIQ0MnXBSsYATi40fsYjQSYxFFvTywsxvOrjzdi33XV1otO0dnHd3UwBX+AKTEfz
9NJXE0HSQOCHOPNkqIIb38lh1FqGRlaL60rr5UNk0M1dmi1waVyBVdEdSdzEJCt8
QvxLPrCZjI9SBP7GCqVuDz3kNWaOAc2tuQfzz1/6qeQjZrYRsd8hRqagbH+igFGC
HxgbCBcMgwYyWmuosKEpTbaprXkCexyJ/CDd3aezGSnnRsuca8t0BwEBCBPQXqUO
OQ5OzzLAEJpvgvlbRfCImYC4smSmv0K8A51ntJ7dwgxVfdmoVrbI22CBzgJ832fU
U9nXTXai6uIA/EWwZ42fvnFHPtkk/0eKdyO7GaVwGNmS4DO6cX7sc1lAl0wblnOr
MriHduDXN+0ChMx4AsDPRZOIABUnyc+W+7yX6sQtCC7Aq1tWpwK7LwgZ6eQTLbbh
F8iWmO4+Gczz1qOXSlbOBOc8aNlyQO7c5n0b5KNfHC+oC3bsnXJ5jLVOqwvCKwLT
HUqSCzFGaVFCRPWbgZ5Ftwmg/YM+V4Mg7H3P/Rt8keh0vT7qHN4MkHxLQVP/j1jy
UIdudfCOBUdMKoeOxo6558LHj7v9A3Oby21E0H4f+2ZhZHVDH6Gs3OrOBfYg9HKb
b6FX9hiTK8hGmr4GKLE0HW1dAmbOK+or2Uem0ESoCoMwOmv7/ZkBcnVoe2rFNWa7
+qB3FjzHeO5xddZTeLPeq2jWL0UZ0UA0b80bOKsThXQEdG+HHG1s2TyfwJYH0iuA
VwBCp/FjOxR/+NfslJqsI3ciVj+QBo7Rt5ufi3zpItUzjW6G8pggV7KPCkS7xKAz
zApVHaLB7N+UaKMhVALOtM2qTMucclu+zpdnT8JEQ8/OX3CUbx+FhEStYN1CeMxs
JH6bt02a6ykpU0QIq1NNx6evGcTmwx/u54Qz6PhFnsSoKGPqxZFtZTCy9ohRjSer
aOffZLpofXLU3L8isulrPWsylWiJug/W8TQ4gRwQ66wX60Tl6DXOcTxnXuVhWDcD
TKuLTp/VWgFbVuGklBNZO2ltg7OE3eBXFvkKG72H/2l4jr4BF8QzS+m/VsVx7gbq
5Pf8l8yUZE62xwiCfwHtQk5jtVE2N/r10jvUfy43mz3K3XUFkh8v3lxZPMLU8MVA
DwDVfCJJnz3WKsVr5fxl6IwR0j0hM8RBh21NaLd8ItrwSsZxLWfAPSYbC0EKMMXx
ovi+xx3dRBEIpgBuXLPmZKcavVi6IqkJNUGZv8KUU1IgcrEkY/wbENKyU1kucSoO
HC2id4Oe92/VmC/FIWf2yiq4DdUkRYF20H6kLFIfJIOr/PxXsaOUGxPrPJXnox/G
NqyC9PdvFPLUR8iuygIUUD1FHjwAjnzqyjw6Ax1UdF+0VNr+mlrBg7Ik5FAvi+y2
spodUGDHFzH78mMmd3dSpQVOUzWAkfii/9SKEweLl6baJAQKW0PdobOM3NjcsGtJ
zn8nvsi6bp0b1oRsPZ7Y7wuW2/GcAuwAtS4fIDs46alOyoQCvqDeQwqnXyijyx/G
xr6yxBebwbTfNQOYaY81NPHGzQmfexwq1bj+wM4pEl4qWPTQh41XWJrHUq3Bu6my
LB6SWpQgZWQC/bUzidl3MSp6JAy7vwc+cidjBtwj12eGwjaZQvWEdVgubJ/KzBZ3
Gz0biiOmQYGfyHLhZ2tUUMM+5DGdorJ3J9b91uhyP2bXSMpH7fgF7o+c1vXl2/jK
E+g4UJuY0waztbfQ2oBoauz/FkRLsboI0QiPjHAO9/p/jrpGre15qiW2yUoWc+mn
mThGPDyGoICdbeRInjzNZbjFhjezRmuiLWuxVkrHsCU4rhGXlMragPknql43+UcU
cUyck1TZZC7JLRqundk3FMsl+VoY7FVTQyOk/7LspjHFp+i5BahNEJ1S9t1uwf4g
4rmBvw3RfWg/bZ10e+nhMpFkhGvbtumVNClA0h90kGXYr+b4FznCQxV0yAdjScqd
txRvhmdxyB8pY8Wzhf/o6v+kOcSd3KIxZN4ppcuoO4UdoUGfeAwR3qu/VLhZ16zE
U5TjCHPUNPTvtCwr56vvB257RrAdsWwA+Wr+woa0jsc9Ik8pxoUOb9GOzTEcrdKy
rx6GqAsyxefHVyJKn0RFQFASu5XMZ5uHzW3LUr0oTppfib723F0czKnxolUkG2Wx
ZwFAQ5S4Kt6hDhq7xdOocdBluYO3VUJiNCOEeqnsJqp6d3AxQvR6tpsXAN/QsdyZ
/C+eyGwybvSsC+LJHiJ6xOZS6byHQflmLekZZS6J3QJZO+Uz2A1aink994zugbYP
M2sS+9c5XJsmpse+1O4e+jV0N/fMJn2gThlZzIYY9JhqdZUwAL+jNLLZoIfBFPHP
4frUFJDfN5mgoXvZTm7ZMPGPdQpr0MxXr7MF8ciHuPlWI6y2VGJpa21L14DA1sCw
EyqjFzJLNgXzBOX6ziPb2qPQwrUpN7ouhKiGFf7qTCrW+BCsb1H/czEa6a21oA74
0dJ2qSvzOtBbmC/W92caUOyILDjEJsGA4qd6kfOk2EpwTMYnjWrsHrhrxxfhzquo
T9Vj8Nj00pvWQgbmFnHQGfKxsIFa/FjVku8HlhEtukOcPgR5SBjysr/M1yHTy18R
TsrpcYF0C+h+R4XPYqOF+uil/RXj5Wa/loPXT5jUw1s4+cJ8e3t96BdRjQq8NEoS
FUh2Re968rKMgxlds7JT8+v0ExI/d69zCTSnTQ08oACQwA3EfZnNIH/ieKnZ6Gg9
AHO5+rqUBpPZRtErb+/lMfkfaUYDpuUzCkH0kLwCFd2cEk9jJAEz3wvSoLSMrirq
aKDi3+FX5wT+8eXqSx1x1TyhJSx+lZOXqjLHTaRWFvNnaaAkJChlGwnys1PYJfqg
xwdMxFzuM7lYJJczQzf4gXima/q5YPz77lACU3bjE/Zgx3w3lxcOd/7hSI51xtCO
nldyHsg57vzbHfEYXKIfYOBvuQ8EOBkiqHw6kQyXzGl0R1CUy4I0gMSDiB8m9JF5
DB3BhO8iJFRXDJhAqEn3yjA3zE/9GWwfPRv4qYYds9FGi6dCv9AiadS7H/cg5KMY
aLmsKKfz+x9UNXVyLtvSOtWb9SXOgjMJWWNbynW52SUAd1Gt5+EbL/MWq1JFOMnc
JhUTThibxIHrA1f6C9UhoCp7I7FCDLzeF6L3tFsxEqniYq9lm0aVU5v22dfNK33M
1S88kQvfIFngqfEj2F/MyHLA021/tFbLJoDyvY/ApXgKq6Xb+/2V1hXXve1B9Ujn
NdD/GLmS6Xs2j+EmeyJ2iL50NtOFa+jy9hwMW6T+GFT6ugw1zTNZ8Kx9UyQtPo6I
u9BXt2VQKz4shcjgML8uUFiWTiljMSzzupbT3dGlk94+7479i5YMUSUYLaKBKrHq
jSHq5eWg7nvMNEGaApVDTTyWhwEOITU2qvElRg6ADqw7ZLfkOifk5kN6Gm6HXr9T
nlG4vk7wSyTcmz6c76et8XY5Z5s0mHJLIO0FeUkVPDVeOllt/Ma82NI6qHF5Om5e
VxF7JfBpMYCcpougX1rdZllwTgaoHY8XeTOZmo2M/t3rBG8af+HazeSWr2wc3fGQ
cedjy1gyU0tXyTzGLXrZ2kuwIa9+TmqP3lHb64vJthrIU1b+Gq3b8h6RFbhu5/dy
VCtK/nQj06M050mSDMWocO5LsAZoxYVauDrxBMjLqhEQiBUqb4exzDTduummHP2+
EKaRmx+N6v2WDSr05O4WB75UNsFGJfqedMYLVTfhWuFBNmOYOv+G4p2iLAxTMEES
fKDENFavYVYwRsvmBjt8PoTwWDRZ/WHWjHuanyIQrAizBq2jXVWAf0JgphTnZnMu
3OGH2r/0/u0RJ2hiphk87LhFALPVch9/tkc+sQeYq6qg6nk5peUEpp/JTFcVYERK
NQxVfMCNfF9wo7Lmh1uaWtBEMixs/hNh52/u3h82kNGVp24GmhYfz4zmZz2aSLce
WeAW2Uic4yl5ykf/m1pnaC+Qm8djR5ctfgQTaJ3XQ2XaVd5hgvNXsIF2wVlWXljR
+/xKcIYQ27lPWNiqK44KccipgIR3rv1J0aCh4YPxX2MDrMpr44834gLe6mXuJjZa
Z62OXx9mcX3p2quEhwl3eE+Bt47p5GEhHWTyiznGeIr+hO+rC8giymLTvQ78qF/l
peYc3hiBbfbvD3fMaXRWaTYrTpk54iwWHJt/OTLu57bKgXt0mtOeh15uvY+xaj/F
2eLH/Vehk+eBP3wJ8ksMcOiNZE4hUUJ2UIG3Q4w9kc9AsmPHZrN6lLWsj4/yonb9
SUF95gJNrjklWR5FNgDBXGcsohBuh9ILC9YUANBtEruy2nGpkzQBDhiIHRlymjFB
TWEQZy3z2Z03e/upnn1MVZ+KFdmWuoBvB0a+Ik33FwNQyuc42MGACFtVuqbZwnrF
ZoDjGPGtyLZekI8IVH5Ml0oZtnEBGTpU2p5xgCzR5EK+4hWMA8VXIG20uUnwjjmK
DdDM0Btecem0gdLaCScAKiIsZ7eW6iKXcGrNLfvb0NTSnaqbeI21tgLsK9oFK83u
/HytwegjIqNJ6TcaLnK17gk0l7cRSdSMzeTprQGDDfPAb0JBRV8AUYpLxfQ4lNhw
4v674YjqHne9QqA7cnGALwowtzrphYKGPJPbaxjdC1HIskcw4W9VOTUuhIPNXMQH
hgbY0CUZ4Dog86zqZ1SlRYsDay/Nnj9yzIvIcE+18jSz4xeVpj2LoAh/j40oz5W8
QS7bJXbtc+x3Ck7Bam1Xx8mgF8xb+dlaa2KEX2TucjOpSJz8ktPz5M3T3do8ZtA/
VkNtwmfnlht56T9bfwrAIVRSrDp6le2ZuGBUqEBgaS2gbk3GARYyr8LAFOQLDC3b
LtdpYz4voaW+znUFRTyCrjvUVxMSDkni0HrkWIVhfcRIDRNtbSNm2KtZWkYQ3qGh
qRyYa9N5r/+b2NTJEvEfGpBGAo9KG0EeyZEHvelhK7hZsIu1QnmxAvidigTZmVDu
QI46VsCZc6hp9sf5rXZIBRZAuRC8oH65lbGbCadl3yDhpnfoh5Oe4LUyL1n4RDd6
rd9+qAMrsScHiuMYStbLB8WViOaFhNdk90vh+cMa8z2pn+l2nXk7aWrYUedQw8rR
BmG2ubXyb+PG2FgZXJb43xahJbscpfG6efQnrI7P1DdjhF8dq6dt3pJ5n+KsBzX6
lbdm+yWILeyTdU2CUHtzB8m/0t6fSZ9fnTAYvGlDgytYTkvXq3BnPxYUtpHu3fdJ
2dLUoIpwtQOnS6xiPtLNJ2J9Bcx5AmvZJaXOVWYUVN081l/bgUT90wsDUVV6jTCa
rHlxnTIOvZndQy17EPYSlIrCpvX8+fwqUtphSnmqpLJ0OOV3oqxtutJmrIjxRQNC
AIgac8wO9A9JcnGG7hYQ3AC1IbxaPUtha0fLuRdb+HmoykaTOXCpUFD/TqWAPb5x
654Ecjbh889FubqZBmfNNu+Q2ZlBDrKcWUcXFk/AFzcgkuz9M/Sc1aDDgzZzzrB3
FLCIFIvVb3E+vi4OZQ16beWIw7K2xVa2W9GwJKBY3OZ80EwYePm76i40JQH2/i9V
0tFzkPD1le2s6nV5+hQUyHX9EvWs1qzy2b6RJbacn3wDiH0dCZt8ewh2DrQ4QIzh
OwtvYqC7/HqRhUKWnuP/XNDJrBSnTLcTNaNN/5uECgKpIh4vaZR94/vAZ3OFTMmb
DG6Ig3RgLNwzE+oSuWHrcBlM/PwJWUVRjyk1EPw2BVUFxB/torxbkc4E9+UXtiJo
4hj0yHZJXzOBuGIFsS/IebBetH8RJLD427RsUw8sebbuQx7KvdmSUq1j9p7R4Vm0
YcUfBqdIIXyN9BCUHpw7JVyhI1BKglNAfmKjtpZ7nNSujEs2RixPyHl0As47F8Iu
FPgrvgRKmCNWQDFmCY1VfSY8712lixsx+ow+/GqfJagMFrsAY/MLpmqL7l6sGen9
644sx1BUWEtH3GmyBJMOmU9UEVFEH/zsPQGGBZ/auqf99NWarRfup9mK8vOVl8ge
u33xT9Fwyu75zeXnNlfECei34q650i/Pn4YGBpaGyw1ipT4sqPunTuSA1CV/a9p4
8T9ZZW/hfGnclsccKdbCQtCVi1rbFsRKQdR1ss1n64vng7qqXX9JJmEGDkeD1GlU
i/i/cAfjAZ67ouy3WeLeziSKYLQMxAIndZK6zGLIcgBczH/DNwPsC2M9Lx4EKkl0
vstzxefTvT8L/+MTcrbXqLoCjSpsgkiNcFmzgvE5ZegortcFVl2nqOeQ2rtueYC3
+nn/ZieMaeKW0/vneM9SyFvS3NxZVN5xw2HJqUB7o6EgtnaffS7XDIVyPknP2TfH
bQVHR7ejCMJHzUCc/dxF6UVdI0Ijc95/3XWj20EYYL86iH70ABJxoSKNZ3QopT7I
ztDYHw92LCxZZrU0GdyRGDoITpew8Vg80MmsWywk7WqcjpasrWNdh9xNRPiSSKqS
vyo5rwkzCCRN9OYa/BjsGBKNzCFOrTBEIaYaVtOOeN8XbVjoF3dLObIMSeiB5zl4
s+0ddkAeV2D8PdBFWr6WrAeSpsd7SBfoJGiBzPTQIMo28U5KrMUWX2d/RDWn9GEE
MmyEkNaQFAl9UwvJxv9Svk8kKIzm9QV1SvsNI5sTokRFKD4zy5pBu1T1EkiqgKa4
xmMRXbOT5qpYZseWlt/gaMLGNZ4OEdAKooyvte2hw3A4+WeDAChbvfCWZdLL5aOr
M1DFoXzSzlEI3gFuDx3DZy/+DM5Qym8hR13CgSBKW6ywQzZxulSe67zfvBo9Fzie
HO+0berzg1spHNNBz7Hq+Re3x7cwCkIEjxSBR5+kvmISooDqdBf1rBDlQvKNxIGE
+gT/X36v/0hqhCS4NMGjF0MzfBnXp1QuoxT+a2q1CU8yzFjU7JprDsu6f4fkvajK
LvrmNg8Z9UDMCc/WdgdHLuuHNetEwjlC84TQPlaTxeqYYu25U7xz7S3/7qAd3/Uf
CKilWxYY5M+39MexnuTfB6dUIZ6I66eT0xCqLUoQekQ3ErzSou6rGdx4kvkFZYpd
gOE1eagLzqOUr+WcYS5IUWzsj/Ec7bY5MyKblNmifSDts0udNq4fIfiBmfIuoWN+
4InG0hYd9ip2M2lWCLP1G805HjK+AWOt4++vB3EuxxOSfuCj0+YMVAqnnSJRMJD5
otQPYgDd/TtU/CKip3VL3NQAvkjfQd7aid7hJNqmgBWvcp11nU3XMR3Hb/7wQb2W
WEEXLQ+/iKb7YG3y3fK6EK+Tmhi4Ib4lqwsWDM06/GKeJEmSjxlaWhDCuXhZFEbm
wzwL3RRMiVYawO+hKgEXx9d5ofXnGFS26ixbt15CFiYfZ0+odMyBU/7pkd18Zi6x
+4mTAmEc1lFggf3tfTQkBZck98lmMOXppxvo8pO6OMo76/DoAEYkn9SqKrXr2WKp
FvVuPS8DKiuWijr1DSiYHjw9025OXlT3rFCCVkR4bopj57s8cjVZvtcFL1+6hYhU
nSZwPU4pRrruzudecTihWInLf9vjrdOWNvatGOVs6NorBw1yhHI+UGv1ssrsLg+u
pnLB05kfIgyNSsGdMcwRD8O8v79J5lqLGVHxByaAvkCCZUWFcemZyYzq18P1xS/B
E0FfRyg3d6qItwil/ha90Cup9p34bT7bIzELoqVgJ4Tfai4B8ythZJeqdkKhQI7n
z763avHXowSks+5cIXUjpJqnnh248st+GcJsv4cKBf71hyktJiq1hdhI6XOQVzjZ
Op7LAdbBBnveFz6qT3MW09evfLQi7yN4rgCz8Efjs+QN9vWXIR8riCTEgZPQdpgS
yIwSdAr11byhcLD25AlUzqjmQrwxHZJbx/RVJVtBUL5r4RO6DaOcNfQZMQrsG3MM
v3bc3B9N72XWxLtqEfZr7/hO+7JgNv0g7rUKKvRPjzXepopenAz3Li7fKsI1YhLa
cYheSE3z0mIzrstob4CPFHBvwbf1Q7y1gpAVgJJFKiIVaMJbHQN3oHkpZAV0TQab
w/XnFlbTOE4YidNewiAD9EwJLX2/AwqOsn9Y+OmmQCfIMW6Ysb9xw/7G9xXuwo7H
Ea5mhaKzSmxzPpoGghflWKz3QUV/pznnOudoVHaocPFVvb9Z/HI1geo0tCwBEkFk
guiVBq/CwDqsCMFwRDZwY8NMWj6nDdSRwXQ0LjhyevmbE6LBhEXs4Xtsyo+2PgpB
r3Kh8KEiaAgydwfNYOZj0BpzUs7biMVwEA9BYM4kxqj84XrzGUV+GLhbc9PYyLzg
9onuDGhk6uoPmqQ6Az3jjNEvoL+2PXsaVkhxOs3KLzGqnxXDxQLq1PV12QqbIaMM
dzq83In3H5/WE5XeL9azL8SAEAjgu/N5PUnYMoFFGNueXb3W0w+TVun1nwQspsSw
RuPFiapSjc//m2F51TygsK2BdVZhsEWl/PM/3uYBcqD3nCA2cBIz8jB5FvyDZR+6
4DEN3s3QcriKnV1j0bjan0lDq791tMBTdDVctYt7HatoodRDiFZMMYMmjddLwM0V
05RL+ayP21/wbQDQpoZtuhzBtY4kWumXq1FBQh9N+T2mnZkfEepx2eJ4IyivfGOn
PUwPKI2+ObzLqnqrJ5VVx2V5U1FWnOfMjFJXZdzazFU8MgeOocXQ5e/L10+1Bf5a
geBw1F7i8PQUmO134Z76TlkRwKnbwR/DkhfMNvncNHVZ4dqSkuXVBBM3nB7c24gy
4ios3XKwxrbf9fQBbrZEGD5fD8iY8MA892TO0pBXX96dqdzNIGkaqQL7CKpCequ9
+eMtcOe78CubZsEv6JWU+RDORpobP54cWdWkaW4cd0XPzTpqr8d+n8dTa7HinJye
3SKdNjo1tm3zF3m8ra2zKlZwSTXCDQG2hGhL9dSBHZ7jmZMZ/Ux6JoYqwnrI+EpA
96JIi4a/DI9K3VGsq+MAkMo4+CJf8o1PNEaxLeM3QjrmRThx6awVR6zzRCqG1DLH
YsleuWF1vuJD4OS+jyB91Zgw8PyWAmWBzhxoNdvztgKk0DnF2hVmu4bHnYLNyNjn
s/tLDdQhY06F6aT3xLwwdBiPQLNNeBz7rS7SglL6q1BfSg1pvC132dZKVkVAwPqz
M4wu0sPpq99nTRxhUKm5wDLD9PQiheqdw3bMI1Rh0eyTvZUPPt9omAF/vTeOViRx
ViJ3dFXXDWkmbaDceDwMxxq7pU9hmf4eZt7tY29rBrlE01YALlR00kBpOHLWKXOy
Jf86FbCj6VzmHi8/3VMpD7LBZzAQ2dtbvHu/bIwgsD/V2Ef40BT0wf9zQejOZp/d
BUVBNzEF+gFpk8hDNiqqcWCo9EkVaDPH1Aq0t7SBXzmzUZL16dmBpEiziZfyJFsd
eqk2K/n1ySsHKcybHe1BqtlR3x0I18L37+zotBJDM5Is0p+4VVlTmdht0rRl0sHZ
QLuo7HjM6GSy02qzyEadlIIwW1uK+khm+y/unndVM8Nlk8Yhxkcnd2/lDhPZBLcV
9KK5YS7UhziydIxO9OTAxhJCKzoGFzfe0HDB2AZk3Z+14BukFjXOw5xXBj0hvrF+
C9J/RRQOjpKCUzVbXjimhRyLGFuiETJKYnULtDJPxqEdSUlMTzTZxbTiwUFkgbFy
SNWhgzoOEeomadfV7AFJuJhGBcFzUkBTUA2zq1jcduR9Or6xYmtK8aDnoJ4pm3HI
XzqBKZ7PB+IwQR7YT+ChTuXl48RbckX45UbOeLQX6mGuVrYhe5ZHafML90+mGK+o
4osIVpmmHdeZG959lrirOZ6hvdk3oqW5coUxnwWdw14Cdz0+dS39YhEtFSht+SFC
7ZZ1s33NILo+ROJvmt4pxZDQLSJIpRNoc2/vpROEX7Leb9ryRoJ94dovw168XCMc
TEt2pDRV1vpMUqduTx0s6P3vYsPW0Q+S5lEycXEwimGzE/ocekARTdHRU/19q0IK
JJdkaMHhqOp/sULKvealfjazlcKliUJXTOM0+6jlNAuI8RpCm8oK3xKrLYAxshm8
kNpE1bvic9trSQAuNPMMIR52Gwt2egSMKrfwjRp3D5oT2EHAptgSbPp6VHPL+N1t
Ad5VvNAh4W3hTPA22fZuEIHDBmd5FFVtoGxupZhy8l2LohjYVoytGvOrxLt7SKKY
fWEYHl0ccttuA2EY/R1opLdgIbuY3xEmj12IpTXMdHETA4NmZgZIwa3FWf2VSQ3R
ykbz7+A42/4H3SQo4zD/Fzc5Re7RYdvq725twliwahvKi40sXeRtRQRD4tA+y8PZ
XYyc2PuzngpN7GWeumF/4u1Wx1uddUR3c9RhkZdzwYBRzZeukonztQqWgFXKjHu9
rMAdbIuTclX1Mxf+Go7N3Kyu+jk9jScIkYNeyoOzKO5uLlbOgmYnUEw3XmA8e5ZR
uElhWConeGHFzV2NCq1GvxKBzxlTgKdyw5QgZYQtIe/RW7ZOwRuMK0CbGfhaUUii
TMHSIgBaLTzgviMv4CV1XKspxSSpSr5Fw/dk/i0L5JsRnnLEtv6OAPzfHQpg3CJX
MAcRGr2sWIWkaMSAhmaTrzBH292gfQy1seWQ4+p4YH9FFAwWoJUKw0FQWL71Vim1
dZWIg9F8je0wPnXl7uDQBeO9cA204JEalDy4F69Pd82N9I/H99b/HIWPS7F0gnL1
k5UW7YIkMHyd63/cM7GqC3ckMPge8RRXkqIBLmqvswb/NFC9R2HALi+HF3SiMzfJ
GGZrHMC9zBZlBdfEMM28jeV5bKPcezt7aGHRe5raC/Jy5idqJS24NrB15U5uDzBZ
Kj9b7H3XN3yub1KBJjEKoWlaIvEFdTeuKvJZKdO45Zey76H1mq8JfFihCGenxnR8
+Y4aUPvt9RPw/rnfgrJoWOxBVKDKcDvbELrr3uaSonqkgEkZkG+XAbDKZLBDQk+8
PJW2E+P3zCXqizfmjcrxzaxgkE/c3lejJmMFv2jpGnbJQmyLntOI8JVu/cdz5EcJ
yWkpp6i0kXD6qoorvohSYuE2XXl5kHa4nCnq9Kj7jkQ8iW2Q0rxaaOsO/BYJXMVf
9wEf1dDnGhSmWY4j4jN+OW52BAoiuL70MTt05f88QQ49VrhMDKEW2IgELcoPQ2FL
YEi/j1rxuGS/E83qvuyBq/EhDPblN2XRrLysLywjGU43WNcesy0bNBY+egIhziWN
yTRZGmo15XnCasuxWmtsrh1/1fN9IiafGVkTDnjIY/zzdlx6dtBwl89TFXwS/0VB
mRNlBNqQ0ok+ghKETUE1e6ev+3hqm5ih1CAA/+5H8S+1z3sEhVG92CPVxFKViM1n
WpHdiy2GqwmcSkawATNhpXTxHxmu7cVf6VABYzZ65yU9mzQ4wUpaUPlcrQvMpD4F
GNIgG1NyhqJyINWk9QZPZVcXzoASEhoRre+FRjPDZNYUwJY9rJMujPzSrj362A86
4KOoIOtkQeuLkyGOtQ6K7HwzVmjVc3Dpp5c8cBDMEr72V3zj79nPEsNH/7pAngkW
IbVZeKTD+wU4hwAf9WWeRpEHY+V5FSKQ4XP2VZwwBqJGCwbTDzvCNQsqzRMeXLH5
rOvKtARYhGgel5PUDINlSal1wp+pMijKJhwgm8eNI+xLQTXzBzPzoPLwLyNLZ9UZ
dOGMV1N7JZVUoYPkA9i1nEmpJCXcmO2uFU+2ZG3yCseG1VFItMIepWFXzif2+vMz
PSjmKZKIQsWzvFxWuhIYGX3mpmv7Ah8xYWZxt9TGwiVlr4zRcyhnJfpmmqft05k8
vuG+qIqCkPtlUzEgykTcEKvPa4oBd3sawuyHJdiZCtnBHYwW5F+5uv5n4QtgVszI
D+ZvKJ/CkpO+ghFYIajP1ybC8LoCvUBplTOa/73kYyrMATvtAtLeHa1OwPaYHcoZ
CZ6cK/E4kcWq4OCRYH+4+ahMSKFWYtS2pOfQ217BFnnN221GFJsiCL0eBNynVxmR
RWbQk6dWLYjgAq1ZWtiBP+a85xaS2XAIdk3TU1EhHu/qf7bbzMXC0kmsPTThVfis
Z2sTC8Vg81Hi99+xeUqdlH+/xYyXpSM7va+mOraNNi+186ju7j9sPUA/D5t7tVUW
iDuU2jMGGQMxAlvMe2kFXqJ9F6UnfYn/Wio5KneX3a7/qak88M3rIbgWvUStQ8qC
+y0Ek5nQ5xr0kQjPtv6OiQAFLzD50FOitwbLjGac/bDP3MHo0L2itL8C7BSBw11r
QbZ+dFGKwIALrXMLrjbLbWvHBVFU5sY9oE6p8cjfWP+IEQboRjnDP5t4XbUuPGhS
ducDQYJZXZhL1Z2+4m6heYd+8q0W+tueleZk3VVdM4XkKu5hVOXiq00w3rFZu4/q
zg2KdV8ELK81t1Bp6wJI4cA7dVnqnNjqb8rLEqLxhcTk8FAMVyFwwK5S0FJmPC3V
jbDCkpxvl8BBbvFlIAPWtPqcWTzCpLNoETNTDmS8/p13W5B2lDWl8Ti1K628MmMZ
5+vE97McnItIy8l2w68+7cnQU19KMMt++YBoQ4RpCm3D2GfwEn1sENGPWlZACKAI
ejhqRkAMKJ+HD9Ehy+MTtKLLlBf4m/97hLTY3+PJaEnxrtZO5+ScoPnx92OtNKhG
JFFkIvYSImmn+R0hboyT4jr+t9zZpMXr+aw2HZ19+q3fL13fGkorBLJD62+ft3YS
mS5AdVDD9RT7VYHnRIvrV+jNZHG1wc22ZOPh2lCn41eK2oaOnGBev1tJjL1QtmlR
m9PfPkxFJgCFZGnmHnJ0fEMVZzTzDUcx4ats8pXMpo43H9rqZU4Wxh2xXs684tRy
l3eMhXv/cHg+YK/ygQq9aP48M5Sw/vaS+w8jPfx7RXNl+ikCwwr67VYu7/SIA/HI
cidNeH9IQUWpAFPA5/xyEN+D3yxbwO6bNlP1MzuMKEETFBSyMBVyVTogLQ2c+GLT
Gg/FlBVJhzna40lcD4eZgcKq3wG4KMtcMCSDebvxm5Jxn4K8264zH9C5ioOiCCiL
0P6YPq9wDPsETFvLiFjVdR0s1IqrhGYjTJDh9QPNG2FKPbC7pxbKuTQXGV0ZFyqK
3NZG6YisPbWgqJWwWM+vPJEFTewTfS6ySYTZCknTt5TkZgcVABu994z+0crTTNt7
yJhJ8Qlcs6orKGhiqgxXgoQ39fcYUaJvoS/8co78NqKK6yUJ3VkRe5KndIW24SRK
NgI+s3i0ODCJeo1INuIdSm4E2vKQydnSQAB7da6nkjCylQY53Ic6yK8z95HrjLY0
mzB60drRlXIpvrDcc9Tlxw5RxJmFnbWzIcdYpvXSMOS6o8tm8bOVh04XT9cM/xHw
Y3qYWan6sZRqn9+76B+juNEiW+wCbtxDSxPQGbJZ7UQMBHetlp22DI3Ua5/uhrLK
ixCYDgVvRxyk+jDWZjNTKSQoii8+JlMyH1rdMEb3s9CChiF3IfmqurTHdNc/0ehd
IBBSCUfHaenBX0xSsKbwhC4GOc8stb851uPSUe8FR6h4y0s6ThvAPs4CN0+FdEhP
MuzwTw84j6WUT3xjILEPaGX7WFDObu9bdugXFp//jfFmzh/7yabgmlubiJDYV3eh
J5hr2ZfVr/61Ts/o57arKJuIXJ8lXZ4bJ8rJseTuKzfI/atsW3e3CiaLcec/4XdN
2ekkiqiHszf9rT/af716qEhiz/63vLiNJ05Ez/UmUrnLOlFOtAlrUtLPSoKGY9ao
EPV78hFs0XRLCI0gxFtnc62sQGEmakK9X7PMolWa8xTRuuyEeiwBOon2EBwlTvSF
jHzv5b+VIZ/eJYwkFtizYGZRe6Ck1szFH7UKYfJ5PaNKbKzWji5D9zIea59U4j0m
0Hw6s/BHCPpmoHWU9MST3nPsDA6TSYC+05OViQfvueCGURpHbgCoFfLKMKbMzFIJ
JFsK8fIpN2eiWrS3gvrBLDI01vXSmRKRjHDiTP+HJRhVduT5DjTkcFUJhEetEJKh
J0DUADAuJmH3Q9TfMEVPVhaiBF3RwM0kopdKgVVXT6MaaLCH/szMrO/4u61WCRDP
9LP8ey9Qo3f++XfgMRPe5fcx/buZeQF/Vy0XilKJf7+COscpjWhw2bMYTu7dxYd1
SaJMKDhVRH/SV5X+y6pwzO7dlztdLWL3X9c0rSFwUMHWl4axV5YqhEDIjh7BI5CP
0N/UXUN82atO1qP5h1P0LWbpNXQwXbVpb73lMOo0125QYpvXhZViTZbGjwmOwIXn
tIWS3dpCjxwPBE6rPJYPmlpqYMT5ZER6evwglufqHu1XtNXCLcCwPCkIuZizHh6h
jWGfhN8aKGw1klrWyN5RVqRJeipTK5oRi8TWmeWJZ6qz5Q07PYeyFSQD17HzZG7t
svafggsBRlPwfmNE5EZJvQt8Y2LkeAVUZVpQChThKN6VTfkITaYTV+VxnDZdhETW
gqZISEGa/LbQ92DwG/yVOxljMBknR5TES+6XD1DZj22/Agw57Q8+pBzVHOw6Ui/4
VQXRYmmUenTmywhgcKAuxYlrVOc7Mgwa3NfjMXhUfhO/t5SY2ZXaCbKdaGb2r1Nk
vzyrnO8OvQLI2EwP66bjnOplD5pJjvI/WQCr+C66q0mawrzU7fJf9rwu5gvsjGkR
5cZKWnwJODXY2F3DuUXXnjzScz0rnCjkXc1r4/UUyTGph90t1/6nBTX2gVxOHy3M
BjZF2396PASiBpW6pfQOdsg4IEnVbVyIch57VgcEpKiscZiF1Zzb0WRXr5wbg/pN
Y/tjvP785nyuCtcmp7zv8sSgpfI31AkFX8v2voFkSQJTi32123zZC05KU29wo2X9
NlTn5PuUSzpiElLz3clDJuPZ5Q7gLnILls/qJU27KNmbjyaQ4fQVuL4Tdu0H+POM
vBtFbmq7xswRgeJT9b6jBWWR1qRFshN+hjm7ViMUM0Jy3jSK1jqmLO9ZoULlTkhR
cTS1vuIx4ZoVFuqI7hkXaPAcelIvI3qJHmOSqERyQGUeFBSB+NtgLIvl9frquYT6
ITfl1tdsmA0YJKMDv6tkUjULUd9QByC6fj6gSxY8v8KnTCAKZXLVMQY9uF5eR9Uk
NDqX9CBEC4yuIkmapui4urL3LcajXyrCv94Wx/q1qUtzl1QToof92yjeZ+x58pvl
9u22u0lPqodBETqnMjm4QfVT1Aqw9Lgn94npQJ212I9LExbLOg0Q9ehjaAEUPfzk
2oHVdi7ISQiN6Eot84tqSs/EBHYPv4LAj2LEbJYiSqEKkXjaY6RJyi7tJIy0Qyqf
3iKHAjkIVxpOIXAEho/mIun37pAU7ozPf7BaH7fZvbjfDYwxSS4T8y2cvpF9RZYu
uSLX50Z5Res+rxS02JwBMA7n/zUy566iRAh1xN3VY8zVMDTv4iM1DE119UwOg0Yk
ChIlBaTWfy4nXtCKXhXold118ctLKssE7lVu9vXIWB8VPwEHdnnSITxNhCj4o3AW
c1xKVT6KqG3VDOsSZWjqBvBDiM4WxuMSleQFQMd/ZWKaDaVLUGkUYT+b0AcyieMs
UM+TOn5ungFR7KB13jGNFgV0YfdvcoV83BibxgxtgAISN8Y7+jx6UJfz+5dRqIHd
YjxQRUmga8e/04ysYkd86aBXsRjaZNKfNMXipEsaFrwnMU6ldmAfnNS9WFT66TqK
ME4Cd0Yultks0uo18/K/UVEQ2OYCWu6DqrqjJIptixEdQUfOrcQzvbqRsvnTjTBO
kEKCeBramWK5LYdwGESganauLujeT+pz82b870NRdWnXpcgeCu0LmTJPUAgDXLS/
QipyQ+EZKSVm5EqBKRXY2N59ViZ59oFDinQ6v4iR3HV1ckrOKjAUsqDWdIWLoFQu
LUOpNbJWQU2W5N4oKZ70DOCWWLVcujlJrFolQd4LkledNLi/IDJYKBRc1VuROWnc
28i1S2A1kI2yncF0LRFVz/LHL0kFr8eURuEMWqsEBBMBVzIZqDNyNFmpdDGW3PBn
ETr/skW/G3McfWQpg+q+qV8yh6CRE9zZvNpkSRxqthXZytzjfzLzKUlXDj7WrmIM
eE57bzyIbC+R0KDtYTszLTSKKypvojS3uxZ1M3Axw16kVsOFhFU+MATtsS7B7xs1
8Ywyg5a3D75CMJkN/Pe9Q49av8IjDbTlddsZURPRGkiONILDFC2xPhdgUyi4bXDZ
7iGb+s79CGOBS1M6GACMZbVwY4nLHzicHBBxWl3Q4YXrq1VtdAuARotCSItJaAbD
ziDOKgiuLkFTL4Kuee+3PI7FTqgdgprKPP0Uf3VzvFM2v6+IPLfmPd6iql+LR2Tw
5H1qwvBWC+DPYeT+V/AFzR168cneelH8Pom0y3wSLieLDW5jmiH16vigOKWZby9B
FvUG7Ash+0ZGJim6OKnswrUDhhQwBSK/zX8+dQEda3/sqTHWRgS4zdaGUMt4ztWu
CTj3h59zYQtJbLNBAv01a7FQErKHBqpPbLLIj4ndwKSGKZ84eZMN0VZ3BU3FUxZ+
IMA/lgXqjU7haNcEIWzq6+1HQDBAGHnaRg0XkB0po9uwIqP+U3KHrj2iDOfSOvq9
iqvW+HwHyS+VGD8LcnxohBftIWAipIqoJhZeJ3D7mKyqGWPMJOypYmFqHAo8KxXb
5BuBjsQ1Cp80L8Umi3+W5xayqEow3RCGmvhYeUj/Lxx9b1jkrC8cmtfv/3XPwHjC
ghbmOB1MzTbsHacu7uKCYeWuBk2TKsm6vbMJhGp1IPlMtKg9hxS6iNkA67/nKmpp
PC4wFB5pwT9SJnCyk0h9YTsknLZTOyAQQyghGKT0cxASglZVh9uBuFeZGRh8jS/1
zsT90Lm1Pc6lEIJM1kfrfiqNQx3FaT2uo8OFaUDv7pflrdEkmSIPtwhDClodmXSi
6YHWjno7kbMq5e2oGL6cesDkLAW+oCJiKK8tyk1+51ENdlnuSNrdsC8Iv9xtCWRM
bYTg2S9OfaS53lBB1laIRuzCJmiR72n3vWpStEvOhRxBnCGPvaOfl+qYN0nhoa/t
a6Tamkb1CRZ2XRc1f6umegaW9iQRob5FJerkCPLTbKiBYtt5T+RpEljTkWVn5ObE
HQOvQrxn+JfvQtIG9GNBZmUOCso0uIPKpUFrtzIZPzeU9+4ex8n5xBs/3R5A3Kld
HSye0FCv+fqKyowSh842O5C8a7YGwpjG7mG46zhaA7oR7OhqsPoz/sswB3Uue7e/
+5mhpVq+MWyWlBd+BlC+Cmz/ZAgitGRJrJLzwNu54f1ye656s6wsF7tCdVSEJWOz
mzoaF9HHlATu4scvQAkfm372kXOQkpNyMql2w6hz5uQN09BMo/PHKSW7R/4R+iFc
WTK4MELoVcrCHNhPeYewHYbbo6IH6hVHjFFm6k0yjPejTxnh5eVrTCNP+guncYDZ
l4vJlk2wj2VsRcvnioObM8DtSpI64+UGKNBor4wV+OoE9HIM7LzBI5q9ehV48ojy
nKQjmj3KjrQqhmUPeBXk8b1t1ZZ71ZTb1G7Z0TKSxTBDI/ZHSIyZs5cQ8qW+oESY
YFfr8IR3xIrj+N23AbKxt81cLHAICXC2UvU2RFrDxxB12lV5nXZUsilCR3BibqWf
243irwWqrBhxYp4rn4ogwI1Lx9oKpSU8BtgWT7wU7sY5lvFgn5S66phQ0i4t/jR+
WEPYU/4QCPf9Xv8udOT2qK726tmUXvfuII71ghNEBlJtvQKMve0JkrO09sOPZs2N
ZXAi+ZXZYnQAiGmNbLUIJkzRjb8f1fXTiiG9QlfHMP0tW4ctZnrV6rMGI23cg14X
OFVuGZeWzMlUWT45nvWudh6pNz1DKAsrRc83waXpXQzrw+fKmh6yah9tHrg5bnNh
EF0oFg0Qmfx+1zeuL1qPLlJ1wUuyI4h2XoN6lpwk/JrkF4ZbdRs5yFydKrXrQe0m
nOdFp9vJCPWzirbvjesIkNZ/CIlp/k+qA57YQxLu3D99THSQmjTMfXyCZSPpZEYh
FmSSp/8p8b8TY+cngwKeCOn82lVkMPf1soFpOwGa8yP8MRwLTZnbuvG6T2hAqRgy
Utk1hCbXgjwAFrNgISjaAJaR3YZK889ihW1dCD85AJO4+yhJsBU6UewES7HLOAF1
l9cnqL9AShXnZS7UcQF2z6fYxMqtyy7Ergac4bCTU59Y3Tefm9AgyOW4iz7sP/h+
VW4HUW7SGCOEDpd1icidtOVKxAPUH0RNPVlkEv5MAPiS4u1taugEOz0pl/lXfR+D
plZlz9w/xy08qoparIKG57jw6QDzvOjszYZidqL+3KwhezYQqlBq4kEVcMMUOwXJ
/jrQWA1oy7bFW2IAyEQJnK0PtVLZGOYgVW06DkG5Hc8PfO6GGXuQm03Y5u9Hq2jb
/RZoQGXtexIHahmf3DD7DUQwxBGi7FeA9VPEchtAtxlWo9Je8RESxJjT2g5ZlfJI
Und11TPCMD+QKRFjQPc0xu9XFrlYrt3mebuY0KGoYygQSLWUVby/o1RID03DZw+O
uOwyBEtdurTzjPBC4zMkiIO7CiAiLDP7QxzRBmUygO4rOwAK8i5MrSwt3UfeRnOL
lLqI6nDNns/4bXqUDttKCFx1PxZ6UmpXVtWzXLk3httjPhUwPRvHxSA+h8Ch5Pn4
sEqvabs6mJ0/dhwSNjvGGlflC4pzQaJDhwrRN5qAYALB+O/jMOZzoFLejKw9Y/Rq
y/0lHUOQtJf26UiP7VCAcRsjPPN1FJNGn1vhg8w3c1+4R94lat5YT9JVwd7N7ckO
UndChcCT8//UWPB2rqLTzcNIhLIyNPxtIFbGdLlQrO6T2BuAps5Ko7IGwWkYVesV
wD3/tFLEzZkLPx1qu0zVBvdttPhpb0sfI2ONQ0YSeK2X0w8/xHK1M6zQXs8VJwBF
6akrU1pgoPAgamoU7C+5x9ExBa0ZnRhqooajex9ATMNgPCwUzIGUZEm4rrbYV0cF
v50RengMXmIGzea30qBM3HuztmyQTzqkxFFnn6GGg1+VIynUljsj3GWRoZVYMkGa
ByDGZ4qeCBMIdBKY+x54vQUcxkcQj3lJSt8URPycYvtEniCS9JDvAUIr8iBcYI3+
gB3gHhjgMK/yEEx1Rh4MErOsAV+JWnAxcoM9Sc27dHWcXglmQNkmVEQavu3pEbAQ
HyW1vB/jPAcXV2GLnrQKVGDeincfCDQszuhQRcSvJ42i4gTwOPPRf4qsiyb3Cngh
DvIbZd3p/n8NSymaRzpwUBDtg93C0EfSmhsdsG84qVVXiqX7/JHNnJJFsBAb4YbQ
c/RXgXkVqxuxDiLfGK0o4Qd+0aZHAyHtLwuBvy0opVY7EyyJ13C96V9/vvyjkY9L
t9HqkYgPnfRUBXstkPZC9Zove8Ns/1YfmjgEJB5htduWBNRddj51gSU6sW+ESR6e
40j4IpFyq5KD96TOxEvGYDiAStVt1Y7Aqlc3YPxGOtpbUBK84X+DjOVhFT7ogi7c
lbM9i1KaiIDSMiVvgIfr0EG0cM9KY6RG7I/kmyV/sLP+cLP0xewZvJKkfxt++MAV
IUsFC4jS+RmmZlvTEFAYhxVGLezvrmJmGMyisFfslWBuvFuBlLOO2jh89P0++3r8
6dQTKDCVpuqEU2/MIBlfXAPUYJl20aD4aRv0iHq5fJwvUv3+to78dzK7Qw1Sg1XZ
fX4TIplOYKY1IohjKgdbGRDWJ3g9vJtItOShHQJYFjlgGqhO5WElUNVRWgO/PsKx
XSDXCh+4pgF0BocuU/YuErKgaqp3UO7yRttX0leDfTA+wCJ/s/TTTq9rqPNaTE56
FRa9r2dL3PAS8NPWKDXOtbCOqaZXddFefUtlaUc1G0yE6p93zsQZO395LxPeqLsZ
Gh+XITiodhxT9adfmmo08dTiTpc1dtf5XNUpBYyeTtmp/curfGn4zF95veZkQE9j
+HKSm+Cw1rxJ0qas8b90iGIE0OT+DlW5QMMSDH7UfDJewvLdOK3QKjfPoazPfkMw
PPa5921R4Tu8hlMVzvB/K2SU54dks5duDhgkEblYhgFReAruhg+6ubWoMlecnmRV
PH1vX610qnd+7uJKE5EHiJNQQpRQy2PzvkcEgPq7N2Xh4kXDTZSQkmzH3sk9JZ71
rXZ+l1X269tOgYsYx+YpjsLI9yCuO0SJLdTYaPI7tWwdGdyL0BOFXPJ5d8RJx4eb
j1fgept1QDHzhBa6Ha3QVPuB7KIY52JQJTzUDopbbh2UVseuXehhf4nBtBWgos9n
f2nqvmjULn1brayVpmuZe/DS+Z+vqDOj0LOR/AmfTexEQ59ebSLqGMRzE+aNr4IK
InvDxqMd9Hqh2Gwhwr/TRr8CPweAfTJ17w0RRs8OFuJ+8sd6VebDIiSyeqdVm+vm
L8pEzt+OUxtr6fU/QRcyw4CCrNiDwF8d1ckGXiSxuk9zJdfsHE2ewFEE5WEdCEMq
b4UrgcOf0tPmY/Nf/rmUS9b1Jql28/gYMhcOG9A1JmuLg69WoE5b1J8U/McVBDw/
qe6BOM/feB9Qqub9LqG7Z/xwN56sNTpbCqLwvbc4oVQ65oLdCv3nV6fG7hFbaV36
U9vMNSKI1sRu822KcTHO5xy3y5s/aM3007GdTiIU726H3C1kywsYeM0zo0u1pAE4
oGXPXfsBbqp50UreXivguXqvCGItywJJ/+b54+aqB4odzkeN9sIYRdLhbyyc3Ake
WS9v540utPPOGAXExi++fXNNyayq/+O0GAZyHOMkYI8AYFwhppTszljquIuvnXhh
K8iU5q7sxGpG6gnGmHxeBp/LmMb+6UQgUOA0rD8FMSp5M5gn6O40sBkcvuXzjaS+
vv9fWptYSym7G0XQm7M4GmVPe64MzZlAlCMUvBEqIdZ4PDj6XbgFdlMJMo9UinnA
H5O7MzLvjO8kQySBBeQ+59m1pzlyydc8o33E/N99XYvZeJTDgUUjv5Z0pDF8LhIR
Qh4RlfL9i4Wm2DHy/rqdatEQoz768tziDjjhPMBTCVEy28Zrx1Kln2CIusUlFAII
ZHQ1T2bZ2SsHtrcjxtBC4UbRoVRquUfLFScdXw4BbISoj2tELKsOofMJMFJ6uF6x
Bkw65pHw+w9CCeUbQgDmFQ52YHNSTFMUU109NHCO1WCG7ZQGybzu9ABl649kl1fC
28ajmdV5PDe4kJfemAFpN6r5uOb5xkli97OhvfVoB8q9YYpav0Csp8Ox2S0oRrJT
QKOBeDqVCeGC5/xJGFEobFqKFXnspCHd2c+y7jMdUXAuFTA/OaVUPOrkRgKilMtB
xREoUHskE/qpbRePoIchwZ06ZUJ6EXa5NCPuMC29QBHhz1YCVbmOTSeHheGXiOFj
cGxJVacyb6zUQ/qR2bgCfuuD5j9Ht5FtO/YxOuwD1Iv2AlHF7U/y8Db5J5PGYLK3
XFDSPwx4ZT2qwpevlaDaviYI/3/7baY269BLQ0cmjor7zO2AeQetAP9BygFuykCY
aQOfTgq+JP1yzVNh3GBVLPwnign3pano1yLDWLhPtip03cOP+9riD2VRNsXkGfxE
rVxoSh6IWMLLj+bBuXe2xrhfxYHoL1oZR5wSUNyYhh7DrHTCrNq1ITJeYzYmIUQR
+C0scrGu08Qy7cSU6ZO3YscZ+yOBt6Cu+lg4pc3IATNa+O9XNzjxRdMdV/baonlE
t4+fyy51qezTwTvm67/aND3dKcOmkPWuChfNv32OykB2fm1yKcYlPA01QfwQHdAi
L10QVTb4O+CLZUgp2TpUaxCE3fdODQsdxUVE6JXP7cH+Lv1mX0EbUVfEmTdp5yZ/
Ju7PJGZR9rXai0/H6RWp7CcSFXsZRBbHyl+UPwd/BJ1O5oNhSCiT5BuRNfEAOl70
IURS3JqxltTNwcdN8cjVh48wcMEaN/xcqgxlshEa30gtLmCA1vTh9DdwFjkAv9ZP
N8jz6lhvw1UxGraI0E7dGzPJLg1fE6IL8OWKOsWL+y+LtpvDqzznWcuiOCqB5dQ+
g0AMEefrvfJL6s1ugQBWZrAG4Rw1CdviR5YuhQGgsAwbX2ztu7YanbfSx+HpX7QC
c0a7GlXXrMrjy0eXVt3srbyAaZUWx/NB9H8SA8nUpz51hCiQMK/XA7RcORPcFao1
FHn23yBWRNexUVSClUrV3cN444CLS3gPyZZdNg6FHxvtmNdlLyvJXW+tySoRZdUC
yYWfEIySdVldur2F4a15n+/BBl+3Mcjux02LS/ypdZJEWWxb2xxqaqqvr5QbrJnr
flkYl4Pwsu+RKPq3Pu9ysNSPGVSXeHQQ7KgL/+f45blEF+xntii3oWz0SxtWhFMt
hRhDqwLJy/nEEwm5/OgmbPf38UlppldJ2BraU7AhKWzIhX1+G4SqjavEtGfVUcpr
6+FlKa1NRH1zk/iygCI4GcdGZrFa86MaBhLPylVeDXL3uIba8Gh4j9GII6JTvj9P
enrgLe0T06X+7t7ODHyho5FsZqVnqW+aoFZTwRV9YXqM1UM+rRCn89cawk4RwTbv
fqYjxMNrG0anXXpC0O1NL+C8MbanB5qHGMtDn5y+OpymQdv1vgv/ljRLH9Zsj9vy
bZ960FEp4haUVcORoMrD8Hdx5dJWhhjflvUFrbXNBpnk0ofnN/HkyZc/MQ2EBL6R
SklPklwF1GHA97KvYqk//NpWi6I4HQVh/LEbsDm8xXhm3zmo0mG3yPzvIz5FaaXd
D2D3qtMshLCzb/C1NVAlWU7pwQL5inxb+eU8B0GHnZ7fIpUEGA6Vv0e6VUsg1mO2
x6gPBSyyEpTakO+Yq+DycVB6uRFaqqow4k+sAIOfdNHE5xMJVvBnXn0Q9SEE3lol
r8LPXdt96skS0NDWL05T3iX6hTAy7LdeEERX1t75NkY+GKVRJrN1dcHBufxRnGks
nIjidWeLTZts4LrDyKvClctI59n64DoXg0HYHWHG1MEFPlRTFGBqN63mKSQMh4KU
jco5s28DthwH3ovQcTi+LgVmZlUo5FeXAmRDHNwW0m+Effy5UbXg62WyjciUAdP5
wWA5y4+re2pGoXbkGZRt4CLx/v2oBTAGCnHWW58Cpq5aHjZZikcjG3jDU1WhUmEA
PTrcOgkQnx8OTG7wHBNPwcJ9bpeBIgN5uK5PrK0vR9ChGmbc2BMjdbqQm00g6ZQD
Ya5DlyQDpEQoFVTCkqxbShmmsZXI3iCCqzgtxSr3emkX7YHiQqSpkParJQ6SGdwL
+4YgUMf1EnmSoTvOkZcece/NreizdRhqR8LrXyHq0CEiZkjgb6P5ORGDIQyZGA3Y
J3LYIN4sPJUmVPtX7c41PLRIZAJO3XhxVLuA79SY8DpahYWG4UQh/ozmyPV1s1HE
qcVzPSlHqi7m5HIRo+TPT4vyT8EHVWEr55qwEdBglwBhrsgeUBvx++4Qyy4edrE3
hRIiz8e3xaHNwUVgTBUICdqMBBrhjaV4bzigS3jAFIBnrbK/hllZGZ+6gbzAbc38
YZSZZt03TesUkRXM6B0rtBO7g/tdCF2KcLNx0enMZmywO4zH1zbJuf1kHO/ZZLey
Hr6pTTe89s+nORIdrjyEFyKsYH0lcpCGoXbyW4XB1mzwAqVH2Cp+O5Iaw6UOQAeL
rvbYB2YyqSpTfbFtUBtjn/zATtyvlQa/UUbl1yp8VfYwbQyfzlozTXbUqxeUEt2H
obVekjRegYN9+YAZnGRyV8naLQy1O6JzNF4xSTCrFnOC46GlSkxEJY1U2gvSSPQt
JJywN9mkod13sXRQRKHoXJtQf3xGWLLoeGcTMuB9ugQZM2cDAzh2JaV/6WFR+BJ4
yn1imcc/u49pHe9rfu344exiJ+Vfj52VdknN8Y1ACuk2BXO2VbO+32jZVyx4yVK5
rG5CO+QIkSDyd1xY3aTFwQC5IM42xIfS0umEvYBR/InlwID8pKnRY+nhAdXJX0VA
cUFjKohZ0J30B9A9p/DNfi/5YueDuXCa7st6TiZs42QKKRtgXG4q92yXgMdAGt3D
xOYXC+d/Rpd5wff1qNWvAXiP3Hgwo0fP+6ug0Px6Vbqh+pVnEEy3JNjgO8AFrqel
pVtp6J3YasR5OG95V3H9KoGDX7MGHbbYgTpl5Z9bYkes1ZeYO2GtMDzQgpi8Zki+
VzjsbxeplRKM/erjaUHmTqEI0rHbKO/hHAAQf9r3smTYIjVxhx2yfLoE7QbhteIN
mG/geF4Wm8ftrfiFQwgrlRt+GE5q939qozll6b0edTOngsIFn49Kh+4WTx9T5fJz
3a39JOO4YGXcr9arF6M1q7c5kyad3RzMVJcsHaYr0u5Nkk76XRvH2ww9vEHSPiQ8
bqlN12lbM0UZPOQEN0bto3awu4jh6rQQ/xqfa8nQvvPCnYBTuzr7c2+r/LP9P3u3
YhvJDbQPW3GZPcUE7cd66UZTrfYXcRUqownHUrpHpNyC3NJQUK1/hLSvDPMhFJoh
BoojTmZGn8dQ0WwYVkBw8TZgo8w+BV9FVu3cCra/w+B6RCrax1/FoSUOsUS+RtPN
H23JVQaLqzjchwgrkEmWQMq1LjsMwb2ekT0mpQTEWPBd4EedAvSKvmz2B0Nn+ui+
WFk+stRzueo7n0pVhFOHWXEr1vSe2DkFOvegpM93T9xDFwmHaPhonh7/qtgfM4x1
5k4lBd3I/8ouRt1YUufHi/2aE3U0lTCDjTsoiFTuzsrjyQ3MGeqSUuW1ZBJjSUYh
QrIz1igluZPtIfeOfzGAflUsDTAZp3tARawau/Ffv3SY5OcvnGl0ar9MQ7ijMG17
Sr6Lp/F6tqiPb26TbCDKLxv70QHOkT4zXG4HGjFcexN5UGnqefaWBrANZQ/1Sj41
yX++JzF82WIvawBQNIptJGfzCkHeInyk/1AdbI4zoDQjQsgV8bfCbXrU9pRYmTL4
xmJ1JjheRf95acsKBCIvbYUPZOqG+unq18IrqMy0/fFMtRdRInUxuZchwUuYyDJY
5O755alSVHOvUt5ZMqvXEi1GCmeUn8Z14PzmQS6Im5Fyx/UYi5FeimTiZYhuFqmm
ORTOLktYl++1qM5QUpucccm6FeW/t7ROrJwwXwsbL0Wya+cnme3ER4DTTVQg5DFb
pE/UAy0Fjtpt4sB7xzkDYgXjeeL41FdhXOsCJgJLWDcleznh2BAgxvrp5SgEE4Gf
3SAjQix/TItgUIr4K34YJUzCPqVVXMew5x5M4wQ7ffLbFAqYMsC6xMySupuX2WBU
phiAUcZIYCMkoV1okrGsXZZkVkMqbUpnd00J+FshHvrELOoWMeWllE11d6xnwAVo
bxm9X53l7xV8RJRuZenmI+43JQZYR5497EtNmOm+CGPZxw0r4rSvTLob+JBXC7bv
6vmI0maqrQXfWonE1DrNsHTU/LzCSPddh7mSYKSZsO5Kxkz0iwTfbCJlvnVVMS5J
XYUVHphdPTk7T+ljLFcJ8S2LKMvkTtKBUGeV4IG5s+viZXypSm9cj5MbFPKeODMX
XoDrC1wFxaPzHdlpFoyfVS6TggtSEVgdVERVKqkJGIU22/1XbbqVcmttjmtXtJfV
SYtJf6J5HfBKhnUsKty+RqxsNcOnkuxL5qmbn+jPOtiDQcbYIlb0yKb+3jo9cv2c
r0qLpguwz9cQuZluEiUC4cS9rDS6b+BO1ClJUoLGNtMRgHEZIqLGYLJ7UlowF2j+
dLEiBNQaTFWbMCKabC4k3Se1EfVEKpWBiAtH3A7tgq/UjjM5mq6CBHKm6M6KYY/N
uBqTMEGXIZtH+Czw3t9O2C/DhwWDzsXSqygZWYs4iKAU8ni9KyL8t2oXYBYbkkSD
XvCfv5MmUU5aaPK9ajzGTF/EAr3ZHpN4PIjpJTwH6VcPs53hg7nqx85WqHeIooCB
QWXYPibMIiK3Jjg55ejyip6CIwjXzvYcqq9goSKtPPVGOfQP7dJqHCmrTRUOa2tb
qo0kt3zdQu1ebjZQ4wEwMHrezWxQWdJnFScPtStINDocwTld11jhNLt1ZcLc0m00
2X+VvT7NfPnU44wo/W8Zr6b/HE5qVLoG4uaAYMCznLUYMNuYL6UFyvrICzvQOpXn
lvDxkVBhV1lL2R1XodAYRHD0+baDybs+vp8iduKZuZoBNsJt89zvGte60obbLnSA
LtuuZj9d9+iFetGRBEeuPQNrUBIAiGaoPF0GhdXaOn/BbdyZG7jL5NcHCbY7N92V
PZFv9q4gtN3WGha13G+PzFUBbOKHcYLgRPo4pVoNHdIgkrMZZH9iRjwuzMRMpsDm
ofR7Giqwh2LFROStPwyI9aXxH96msJzyNQ0FtVIrXIC5MUihcWrwA6Avb8Ewb6ot
ZeI0D68Pwr9g/g2BtkR5pChObN7T6ZY3D0eA9O7PdB+UwISbJunMZm0Yb6gksuW6
E1aWIbuj21fHDiiAvrMLI/yjuJgKadUeyD3/LrxMxlWLpg7YLHo0JYO65iPHDjeo
RuH4ZbKR4r61KUOaNLpymgcTPVmXR0ePCCfbbtMe0pawXUCXCrn/0umAIsSkex77
Uk5HZIke055Aghx/KbC5oaagiuSK8EM8ljc8ImzaILGQyRUTSuCY0wgrQjnT9Rgq
yFsR6nFRzg/AstU4N5iel6ApEajzYPv3C0KJZbOFgbzY3G2UPZwhhSyJ3rliccCB
gY6Cj5HJRW/l2EcDbZuOz2o05uPngqicJpcEaRjAjTJVYyS+xwFjLvHhvAzj6myL
49qMR08FOom3yUC/OFcW0zoHE/deEXCfdDOfG6VKYx1wvFxkzJo69NLl93qn1cXC
NodmZVj9aXx5d7WcC5tYJh0zfLX6hhTF/20bhHifEh3yJpud4VU/4A330fQ40sOr
mPLl2IP2DNc5EFLdGzl0nG2Cm/dL7uSG2R9P+JZ8YB5vs6PHe39P5pfdUScO/HxC
qfN/17kKX4yfxy34mnr82vKVagbJm//lWa2RSwBTue4+THTsAU/pi9AO5+gOoSZz
z6sjMgkNA9WO5FxPxc5MP+vTVN9bZCHnnNiO7bNhCwOasDKBrmwRhxiXzaIFAzV9
c71px/iy6TLlRqz9EqPDUowrWhqqmacJSHEgKG5Ld9jTrKEOQixO36lKjH1A0oBw
vIYlUIAmtINOPLG3Pb/Av2orAfKI41XA8vI18fq2Pc4f58P0R5ZtFHXRhmlajzxN
PFAilTalsK3iUBtLX2zSzX4z9agSKk3Bcm7rLcKTCmF05tVtXfLsoTYO8++M8KLy
t2GhIWBhNHbcQyzZc+DAN/knnC8G9hseZFa42Zdz/3Wa4F0+UDSVOiwTv/qiDKRm
TAxmtjA9ZzmTYtHy7YZ0KWvdKa8Yj5nnnlFPcD4GVUl3qvX5dDuUNJ+nyjpldgs5
FimYChtVp+ywrj8pE+jb7LI8FME/KbwQRfHxVeRcI88vvrmAR/+ZxTXlEiIIHAAp
oshgEo7nvknPF98SngL/nV5mey2r5AOK/drTafXSvuEh7yFGYq06xNDoNO01Zi1U
hv7HWgbMLzOCiPwsUOYiWu+hiKIZRVEkhKI853dEKtcpOypxzFuM0B34iVGeUUpc
P8dqukvYXpV6/o/QKtTf+ooDnkFfuxU40moSLZ5V4pq2fjr3iL04QIlumiZvmZnn
5oG2yfp8GQJtI4XDx+Rem0bpCENXELZdItyP7iRHZpEZSYQn0nSey6Mpmsb4/PT8
RMuCSsKqcVVMjVJW3BUAZfSK6dxNJvi6sqRznJn/VIn9pq65+kvu0qQptnq9MqW9
ucGgq97dXD1ycnIENbse1fNTZzFzSdLpBShxRwRcPOGojmI0qt4O5xBoYTM7CyYH
vDtzpjKO7aZ2PbYGtXnnzDjjxyjKdDyFyv8Xo/0v+Dtd53CXRa0IUmlwK9i1QzJW
RwmcTEvDfop3EZVd0eLVMlRfCTlGnc8yqiN8QZoON/QxRw40hY9NQmY5zFYZ2ZpW
+qLuuynMWFqSnzyX8K7Rea1+vQO2WHkDkF+rDDc/FSuJb+ySvas0HnOq5ZPwGiT5
5Ni047bM0sWCSYPKUQKHJfEGh0Yp5ayF6aq03W1AfWzRd6ezBCot/wCYsyyLqPXf
MJyBz2UAx+CEfDP9WKHvGZNaUkLjEgvbVL7xR1UpkUqNEZ8igXlun3hMDDRYEHhY
+M/TW/6oQGZyyF76ZEBhAlpU2KRqZpxdRokqmlMw9gqW+b/EwxQInaGEPVJBXOP6
AAoznYNxlgJwnSZ0w4SwB3vxxmjkl3imyBNFzW+r5bXh6Ra5KEviNbU82gWRS89g
UsfnUhnkrqjf5jo++aw0pE8yKrWb9tplhy92sHF+oZstOhPBiDIJibh8MucHUhUx
2aNRbnGeCSobaKfYHoQiejHqr3Z8pXH1XLYVOTv80aWlrs/PySGwSFZI8gg34PpU
PAbe3dGYF3wY7tvIoVNM7fUYKQSp0RPwtGSYisfmJXLWa4Wvt+VO7hZaiMFXGSxm
8j51qOadPATktTc54f7LKaOI7TQ3qXwFcKvDF1B84IX6j8fu1alB/F0qYCiDCIBz
mE5xoGUKBW24XmSLjhRznHTSjQ7OMutRkl3zJ1uj+maAGymnzsydJOCgiF/MsjhZ
uq/0chgkpdjRY7QR66AXM/UEWAuUTsbBjKpmKkctGnpBet1hhvqyhUeksUMqe42w
47/jLl30UFKPzg8XQKcQxdPuLY0SEP0o/gdU9OBX2sG4IbKCfRTsy1Es17ma4s8A
Oqg7xWwJsDXwxQgN2G+XGnqSiu4UcVR4TYDWRd6VSqzOexZp6eZQ0lPNs05EUIjt
YJcmQsRk5qKVDbxGJ03f2EAyMlEgQGHX4l49gBleGG+0INsaYMkkJ4PlrBo8Iiav
o8B4nqAdgyzf5CvAj+03POoU9Po2NpeTHbtwMm32XbnHblPlOqgsCKGS/vBA7M3K
FSeGkCqhItEcvCdaZbJHA8AR/hXmQ99tC8ebH3csnppyVBQ7kv6zzXwQv402N+8N
TmlK8aACK58Q34LU8IF1JtY1rS1ktW9EPvZg+7HVL7aJTx+XP5g4yHqqms/xQsmS
pKWPlRM5rLAIWSqLchbnmA++5/218CXpywGGiegN6fL4v0sKsKJAF8UJb64TQsI8
X86nIumX6sMjy5Ey/iWq+UFeoD57PTEBbBGU1zxVUW3U8HvJELbBMUKaLhPI419G
L5cWHgs2d6stPbuskWRJSDahc4WyAeHspEkImUGxZ+H+nuTfQiLk5fZM/haypdkE
OvSS/Yegr6BKiS2kOLvwQigUl1IZR9YlR6gxSzAEGXWxlb51vbf6wYlAgXTI2XCO
7cAVABb4PsaM1E8UjFyaxSiC1fiF11vwxRSfg0fI/yzNhtxHehTCwZFYkak4vsLA
tA019gH0JHoDwsDrXWzb72kS7mtPhId0pboF0Cao0z1bYpYweXPGz0q49cCBnxUP
+lwYR/f8gV/lwS8S6ieaErhbh7qfFkGT1kGA1FK3fJNOM0Mb+iMZw+HQBU45ErJq
kTQSLyrWXVeL0N3uzQbSlsBopD8jnS9b6AZq/2dWVoU1tI//k6BykQdoAJlydzS2
4PmilqsrGdv1vdV5QbYzi5RyHITMooySy9wkmeT4dujR2aHyrGifJ7vrSou6FhOT
dkvNm68lxya2L5otlmX0YE+M3fXhI4Oxk+2WHsWu4106wzZgno4WCE2VYnyadNeM
/CM4sHCcM6Ul/zRt8Sa9wxlqbk2GuAOzYIVOizB0E5EAHdFhnvA6j7nJrjxGJ2Ow
wYFBbHbCJvffAimDKJiaN78BuY+VY1P12AcunEFvwQuv+T5I7xOAP2HqtVwgBfxA
4i64FeQAPE1b/Y5F5GcL/jUA99NpUF1u9P3P93vij7BlUVEdOzB57iIrxIayJ2zk
dKkRTnTnzzjMJqnfMYzbsCh0jj9fWRJo6STfViQn/o5VyYcrUVhPPpVDzxlxnhIi
qPGicvmxdHjMl48ypwJH0xbwxOh0Im20YTtFEHKDvqbbhgBYv7FELRytW/5URWK8
F3+vpsqhsFDCjq4sYZ7PBK7W9whWtmDmH2C6kCdA/WKZ8kQlokjp070ZkZFNmAaO
BpRHVy6m1v4wKpd/v4qf+QEkK/C5ZAdVjoU8XC0LdiTSXPSPrd5CxUZ213IS19Ik
Ywtu0NDjDb0I+PbGUKZsXzFYOZzZdVnKMXYMXCUtPRijhtl9IaZbUPRKN020MPBi
RYTax4nWB9OSxR5IUz3enV6q1HNplP+QznE1pi9nZWXooP22j3NbEWwAVpgIZdw7
E01ubbQWhxUhmpO6bXcmvCWLS//HLL+0fSKW8+8+Gegumv9xh4yvoqtdyKZYGTYH
yL9xwSQsK9+GS2BY/7UkqW5ulozywHmpcbSEyE0h9vmHyY+1yv2GoX63afkdQFLT
V0O7XgNF3Vt64l2NNbpXgIBopik1lPfNnCL1mU8Hei2JOOrKkRjm4yNATZ0eCsrw
QINfacqMqioo2yYrAtZuqjWqCa4zH4JekUm/sJvhs4uZ52Acq78LgghPz9v9NcJC
h+cSZpQhAQm9yAtOotAYIYKeAUJfp9sCLiXqj9Dz+EoRSx0S9EmdwBSsez0AQpKi
mLnhpOLHOePfRxVTnF/83BaNetfTUjnCjwcR9nE5ENQFLVWQ4A0ozblFkxhrYoz0
wdmssF8VcifuKhemaABXPN/XiVSL610HYJtQAma/HGKku8rjCBQhUNeh/fQvVVua
E08h/mpn0b/wjdL5wFVbsjIEsXtwtiz/H5B/K3VRRuTWJkpLv8nrUIPyGPk8m0bz
0+jOhPHkdXjy4ZVcwGpo0ZEPp30nDmJFifpSkgpIY68HFNMx8IEjqXW5z3Y1MH/t
gr1qxpaiYQu52EV9/Qsb/X5z5ESyJc/RXywb+kXNWmiIIBJ8J6pfL/mVii7INxsv
CXJYooYLS3lC0wFK+xlNGwRBbqQ1Lvupe3aHgvA/KygUbio1x5XL8a0yvylUi4/t
GYnKO48Rj/rZi0nMYHkaxS6fDUQ+siJTq79F2Ldzwsu5vsQ0+y1ds7sOxTNBbNxt
OvcX9lM2XRdewMfb+5tbw4vw5sni5sIOj13dhkVpmRRLn2kjxQWHates0zvrf8iK
EP8/2YQd1EjWSrulFkeWPDJC2MLqOA3WstlM9+57KMYjMChNgbBC2SWmK6B2fNb1
cbHsBfPeX75Xx9DmR7ejccLDkG+YOtdoPnyDcyNLBaa23G8AQGgBM8BlRCrdlI/j
zKGnJkQk6cLNJ49zq3u6towmDqbki3OK+VTL5ItSctpObGstbUuVesjFOOrPJyXD
G5U4ZVWQ7WW31tOJsGFTNSCN8PxewbtOZiJv6lAqxwLe6LRbBrZWg74IU71Kq2ov
P1pDjTRN8KWLD2qbbjceIKBEqLjX7kfeVYTOjK48yN9M/W+IbQ4ODQBr2NkmOCji
3dDKBT+DAyv+eaiF9p1Z+p66pTvwFYEOVuAXefvSl0DK3MOHIbSYb49qlV33kAwc
S2zuRPJi5FFXu/DHvPkkEQIlOVL+5W5f5CmZ+PzOfRyIUVWRGTA2qlHj1PW3rW5X
mIon+VuRr/6vOG4d4ku9HxF1JWZcMtrLlLCerFkqBMdSbqKfKObeKHpihZvZGk3q
5mYlOSyFVFEtSMtGB0pKLykU7ac8wHy5bpZKuKLOVmLNlHV96bU3o79pUiwgVpiq
ekLDRfJCoOHMFssV7w9RPzdc03uwlCXi2Ul7mlSwpb+StQp4UHPSDDtRUbFk2Cdu
LFgJyrU+G11ovYdWyPX+pflbOpr5Zr1Dw3UYN3ZPxbBZtZB2vCO2Yo1CRrLrJRgS
7kYa34zZqMzbApWTKZo8RUIuAZkTmHXHCF7fwAH7OboUU+Rx8md82j2YfzcZdaYn
fazxNl5qjq2sqbdkXB1RebFt+wltVX9LmsxB5lp+a9Px5EKu5h2f4i4HArrpDBBi
8mk2/2+6mpLZsfV6kHdECUKsqWc+L2+KEs4PYfHTB8ghZjZqk+Nh85HJha68AM9H
ZghdVKPx+ea37KLvyGKr4Estr5xqUiuFcOrWhaGhO84+vRy8uLEvtsdh+RFnxyrz
7lCyRZ9lrqdHK+HeTfZwRJ3Al/An7hCS/NamEvEd4vjPoEM2QPEHSfisFVKx18+r
W0pZ/jlFAlqQxwIP0snwNOA8RIoLnd16+V6pUbAlUMmD21OLKouQx7pLb4cH8X8N
XH214hv+0I2GOoilU4bUfrRkW/KT5zyKgnLppbpAKKOiiPr6HaOnhnO4WiYwWkTa
MTmOgPcZgsw2I3rrzQtnAznvBlMum4vvSLqcDrouQKqe6K/x+ozHAifkzz/+BNx7
xB/CXYwV1yl8hB0n1HehdYFdpOv7P3rBSZIdNjp2RKcRCFkHR5c0uk9p0x6VwnKZ
p8+1XFpnevIfxJGCfcsgeDWEzPZC44NA6oWC0nEU99OFV2WaIwbNwg4+eaFQankE
ixnQMFBic8GtcscA2opGaqIjNb0V3Yylay5CggCTJD28RosXEayP92Utf43/492q
k4p5iJAVUXwcC3C0mNSAkFy5Gf99bH6aSWl+MjmE9U1lHD2vUErBHZ3CaGMjrM1A
tz7zfiacxkdUqCrz2fqfl/FdZRX81LZ7qJTHGudJZJsaxhhRa5lrjQgqDdRyxIPF
BGNVvuL8MKjEbvyeSFBIh4hrVzWpDdWj5dWLRmln84TVAHRgmLPTf+A+5K6aSVch
VpaVCJoBtPkhROGEcOTUgBzJ4iyV0olH/uhLG2UupVbo5iBZmHmwQDRVPKVhvAKO
DLs8cr5CQw4jt3Cw5vlfn+7cfGcHJ4ONLiDZ1KoHdTo3llqMFOla3iEjv7fcTtFA
wt2JTELzitxdSRySm+yLnthLo/I/SK70C3mcPz4n+6ewU4VbTxjpZOVZHDv7Iq3I
1febvek22jx6wiMC9vNV3a4jB6nyL+4tgpEpe0orkdBi0bp/LdJymAyNkwqxAWzT
R80bPrxh6F5LKx90IELVGt2kfzNC4aNF1Fe6CtqCljoYRxAVsmDth1he39ri8hcO
ZQtwCMEj+uz1FTfsxnhWV+iJcLebIizUkbxQjDf9FecK0fpw9UIHA52ldwNS0oWg
L40o44AXfdmfzbFOWrtXxdeaDQ1M81jQVKXOW9VLFNwEWQBqrmGgNCp89Mj6r6su
3JG0YXqfIYe15c2jDfXE++4pc/RTlJA8atLkW/hQdlLdrX3EDnfZicuaDDp384Jc
RY5n4m6nygXRzzKGTNZKOPLLPQhyhTpj67Y/NT2vgHyBJnWwCW5qG2NCT5t652S2
VIFq7rG3/6bLqNF8NG4r075yzY/HAzitj/OfkkE3nRLHqskdbB3H4AfZ8Sep4lkr
EyEiMHS2wBDWCBMg7cxogpxnSdcFIyl7MxDZO3hIpIsQwo+1miysY8MpfJQejZhn
R7k/aEw8MFS7hjzB5Ex6VtvhWQLq3S+e27nPLomUQ6nRVsnLP9xqhEZEMBYEpmQ4
AerrctET7b2JSY8zLK7leIG4IOB89bDWckeanVEmYH1sfvblSz58CZOEcamMnFGC
MuZN6P99Af10hJchpDl/o464h9HTzoGH4lcpOTh7l0mRqiqnboreUsoQ9An1QdFv
7p32MfC/fyIFVPpvvmoZNz1PVXiVZXmejr7Cfqgf5QiLU9cFFOKaDi1HaCKpg/cN
MEnYF5BvMXDhe6tJpim32pt+untq2NP5tWZoMjET+Sj1JHo+mmvtX47RYr38Uqy6
rlZ8cr4OR3YLdWVUJFQmVjs4lQC1KMD0DAWz9fH7popHmylr4MJ4tdwVHS14Y3gK
5C8gpCL5NgrCDAfx/WYsC7R+Y3w5dUR6FpC7Ju2crM47xjTPNPpMyLe4DPoOOO53
WBTLApsPNtooe+PZ11chgf4dZekfiMhwS2Zl63Zwj+oLkuyYCsmh8aVUYC62FqUh
ieVA3fRszSOyJUVd3TC/9wGYtd7GzrhNDE0NArPEUMQr3SEbDK2OLnqb1L+irJ/F
R+iCdLKcxbeggRXDKfu412vIwCsOfT29cJAnCpAHIIyOiqbhmwazcJOBj4mO/J3H
PKBPEYgqUWOocH5gHmqsH/CTu4qweXslrybS2n9BizCBKn1PWWe6NdooF9ljXaND
7nj7CmKP63q7Iev+ZXTebEDZ7y4CY4TcvF8aI1GuD6IOwaaVhUU0vCTBA7Kj9tZW
53GEvwsaVdo7dCtMKvT33ruWhpk9nX0NFD30QQem9O4xA7QVn8QF9ftu256dLPOs
ZArUc4KHkRD0jkgpQuKskeDGmFeY0eH7B/qUGlUC7UjkpLwVdGKoZ5QzosdwnrWS
erGnU8X8BQkaqLKsGZ0CyNHPFczZHSm5zRbnKPxTs/vQPQ61NeXT8RdrPGG51Qsz
5gXfQ+P1yoEBya1E5DGn7akDsgVwJ6JbEFztjp7XSFvJTF5ZpIB9Ii/sxXLOkkDN
qFs9xwTL+WrJF+iaRjCkDN4484LoB/n3Dpzk46VLvwIUJMP0tKQO/tUTDf/PCaGk
uE8RS9hFKcetzLDeJpBZeeA0sx26Qf7j1IsiQor5JI17qUB48pnW6vPmivTaM9xt
8geIvwygUFv6M2K5cdOgiAG1jl6BcOVLKq6te+iUJFbLoB4aiV3+uNqyuRSaUWxJ
hHX1DcBx8Bwy8CMa+jtRBhcTMiG/7nMe2WKNs2q5slPK8L/MI9MgKH8Dmt5CQQGw
DfUkrxF4Y9j7708QzYJg+HYH2rZCuXxbvcet/XykunK+5+Wt36c74VtxeeI9DnAU
B5/yG4Bk9IKBfwAKTiGnl7mFDQKRhdlMuMh1+X1iMWxM30N3gctRSequ/lpdgD3i
h+FJcqPyXWlHpGFfh4gEtcy1WA4pD7zqNPGPDd3zZT4x9z+Uinelph4qAoGCqi9S
CQxCabyP5pjESrWVgENu+Id3ep2HZutnI2NTdoJ9lwJhC4JJ3C/WzAmWtYIUC8BB
L1Dsb9lxglnBJoVbSY6sIdlUgwKihjoWCUCD+sbLoWcBGjY3RgsDCWfqAo1b1yCx
FcpBqMB4gdOGeraKmNPFlEbxXqeG1OrTW3q8M5U8nsT7EhrzjIYal8v4s0vtKlGu
j6xHSyr+D7GvTVnkons8Rmk3okiap7xI23iaAIcWyxLOYHa8huxWsq0UydsoGiMR
JSBoHJE1AK8m7v+gr3KtawGTczyn/r8vc/uga7haCAXfiDr5YQdmVh8Leq8BGobB
MIEu/8wMfMaTwjn10PjJx6HVslJM6Us+LShyGVgWgJ8dn8f03JGHUqkVjp4Hn2g5
WCIiyiHzC8/8K9/20eVpKvcbe5WWla3xy9oSehMK3aMgYJ2ObiVuhERyQYUJex69
do5VDT778frOMJiEAsB1G8JCuJM8H3UKO5M0j1gOa9ZmV5miOOzDpdA4QlcIJr5H
OaMavahW4MD0joFiIZZnFn98/33nMsHq8MtVwhNu4WQXWZdX2NNrZQk09hmFFOJJ
Ng770OuU0ojVqN2xj0bbs7641+ZxZzeuiNDFUXos+V/npyquXOJpDVjN7+ZLSHoT
sXHnF8+pnR9+X5hcd1Tim7BzFpmFOyRXPu17zD5KGIqcpeHT2HldMHOEILO2+ym5
IUfuu+WWNoxIaN4uj6s/ilvcREbjawIsHzLe5L6e5kjb1IbbWLyA8Y1rHGLI5/dG
D3aNrryAb/idfRqWcw+AWvTKfV+jX/8iN6iQwiyckhq65AMmkAvswcsI30rxiP6U
6N6DrNX/aDyvew6m1icSp7MlYXs3dfT4yAKlNF7QBeu7Znq8Cd+Dwaz59mJIuPuv
Arys3B5qoLO/02GoLdivJgOp2Uo3abiq/L7k1Z0YUSlfAW33/kSaKj578b9wMld3
iuuKQOOcpA6gdYxnIRbyEfeNvtQEmj96jBXRgKa8pst+7yU55x27zy+y12dZwVAP
er2yEPZ3dLhaX0aB5buRvzbbhmnKJZIJsDJ2b6OX3oLfPVlDw8zyp7+pHEDnzyAm
/Htf1O208Rdagqvnnt3FXKUzbWEQE4Gs544EjVNsfSamrZnyCApcTqheHwInoe6H
UdrvAPhSq9CYMUqBN3RcrEhucx8mh0EFvktvRasOvXz03w75hgGs+79PgsNNgq15
cl32GTVEh60z7cyObd74SutVPXvJfvJEJYSEoHqTuvLN/LC4W2PYvzO5n38LsP4D
uQWG3sBJIDA2PQG88deam4ayshcMY5r23TSU3CDIxVhUN2JoKltdttWvojw2H6UI
Eow6IAjXKkY22ZjB2gbgSc6acbsMVhh/NKv1bH606G/4fkolBab2O+Pv+Kmu6e7L
66vcFLTrur3JielFJijLV7xBeU3qilBdFV/6CUEwT8Ipmf9kzR7RVMalKhVf3hff
tOBtsS+xcDpI03AptZ/1Y4R++c4MGnFkvH8q6Iyqoa5HcUOjjODFxzRJrLw2LRV2
TpbplbnZZ0Mr8sEspLIARCmEv1eFDvfnuleZwr/0JJP9SnlGDpMvRUyu05/P74za
50PYYoRv+5JsfweCQZz1112FKNZUsky93vj2k23QucylTv7YxCzd0bJdv0j4Gn9c
5tBKiverEHfNuDhEDGpqVmM4bsUoaQV6C5fcRn9B3ilyA8/DDO2H1VvghKaeUHce
VbxH1AZiPje+hJ6g9okMrvOl9SxNB+ZxS3e9ZGPJompdyUsgOOUvHFgtpS7mckFB
XWuNBaG/p6xVcV1J7vGLfjpkuuGWJB3fLRfqme6l3tU0sKRpBV+3Qdos6R76wVEN
gnjjPPMiks0kHqqwwFEGeXBgvH4phlfjvcM/wQ9kav6nD9APY7hmJxANRzFp8on7
3+vABIGDhFIiztgQqVG0UfDVJZf7F9gHHIv7OtRVyrV/MbcSOOC5rVo1KCGlfr6h
VTUQddQnoWgwwWth3j7jMZ/K5WB/2SNT7YLvF2f4krlrV+H0cKCETO9wZKaTAH38
OZU72+fe+drRpTjipeSROBX+smrWC+sDxNSklJc8/j+khGNRF49O7XQev43mcj41
y+MgteaSzH+nV5d+9jakbjH4rGZNke/WUx96RW4fOltrDztSDRgu3qVRVehmfBYu
NqQPE8wXaNwgFBLFCp8X9fU9eV/HIsa1e3sH8emi8a71N0xXyI8e9BqqmWEQ0Z0S
qoE4Q9sKDTou3Djc6bVp+NwsKOZ1A5/j/Ft3gDt+9+8gPBJCnMru3CyPKtOlnyvi
NfWmphdlkRL32/r7vbgj1KoPKszb/8OIhYYUZ1cZHrOaSVtRe/tdPlK2ZYO1ug3c
8SUE1Ey5YD+GKLmeTXdksfc3yqESvvuUn2uoq7mu/H0VdadMz+G3phoxtT66s4hM
7eFjcqN6IZZxVRqHupVbDhZ7HDkg5lChrZvEYtMYG1ic4cEVV6bnVoiOwg/1Jf0E
Hq1USabe8O9VHpAU5UD4bPcFI2vHth5bXpTuMbHMz+zPXxDrWEFwiJuGuNC3tbMu
+VwRr+UsIyW67A9TrpuU9jA7nnMCvHXHhIKzAspTV/2eAO7Bz6raU/w55ts58yzV
MXySDKOg3V63PK7f1uhdAFikqa68iRZi/AesJSrW/FdLDNVtTIty7Hm6eYeXjLZl
mkmbAL+VuBGbvXFNtg/V/bOSDvIT8wsRGE7Gl77CtfAUNdAOmyjMlf3kPHfd/NQn
3Wvhslm/h4qh+rJgpBuqOw7AloidLWujrWlwegllqWk2ZQJ83034P0g3OB/dMhLb
0kppBTGDmJDpYtb8UBBk8XNScqK+gDi4fQeCVoO/BRABzAgg6x635JEB86Igr92c
gAFgr7y8aQ0sH6TK82OUco/ACCRadUnkt90sEBOJC0DhzJDNbtmtTooUHrNJGvN3
xyBpP0gxWdVLzWNJVZzLFJpuaydgCbpIY/Wk9oDlRDS+18CL5HAIsmTWViefKr8t
2oxVhaUnjORt+v0hDntZZ8XE5Q3QLkCRL28HM9rwP+Wo0y9m+zCR2lISh1/axxqF
I4b5bezseRymsLc/z3tj0P44jObV7qhifvtMhUFGZpWusDdIzAOBtfvWo1GM3k+I
O5HBqSTf69wjQ2Uryj+3PerXfoE79xmHsSx9wSAvZw8TjmRpde+uh6yc9e+Lserh
C3TbnpX5t6u1c/jXAxuTvzxW8QqwUvTvyEUqVvyfxYm3UYVZjjX1tUBjAKs5Zwbl
y12vhWKS/5mLcoYpN0Iiale9HfaVxz0mI4vohsAUo5lE5Y6A+S2JFxG4mqbjGYZE
uQiUt1QwKW0C0ryixIL3WNvDLAZzarwEmTavFHGgmkOOBIk39wW6sVt1QlVN3bw1
j4lhSbUVQpVeMSKDlM5HJIYksfct4SqrdDuwkB2JqV77uM8QoV7L7VRcm0T8a1dI
mM2X15CRducr6aabNuGvyoHBoxDgUj2XXm0ifa9DXV43rt8aGoUuGKa8oPs9Q51k
+gg91svBUbf02bpSrhefW2K7UvIrYPjGvpj4jM8Ya59pf6jpYd5kJ9YfrtN9nkhK
/iH97AWSl+Cr2xfPCrb8BfFCqIdxlrgbhYyw7hShheiKbHHt9nJWKvuI66UD3Gp6
RtncuC2ZoPMjTVXi86DTLqv0Kyvxgy02lIt92jJ1gpRWGuzJfi74X4C1NyDL2o6J
CAs6x0XT/Fk5dXXrVyWTOKSucfhRaQa3doOugA4CAq4h9AbJ54ryXP/uni2gZQia
zqwYEFPm1rm3BKhWNGAfMRoQ7RF/xRMFA5KvSWM5y+X7E6653AtqvXd8u2+Q0TCL
Cjpb80MXA+ILfd5jdEX+e9JlaYnQO/ynfDVmHOYJJg6tPEl6zQ81+r2l3AyQlLAZ
PmlEabP1yzAGnvrX3PnWt3KKG+CyU7T7XFLYHh/Hs1yQIoRXOttmB5CzZrvbl1g4
FRKALJtprTGnyiBu6l4z1pgGX0jvPrjKcn2hYKKiqmt3AMPNOnT2KfPoYxIY+WyK
ty1v7IVgXZ/uZ7Er+Pr7/5jewOD1oHNpZs5jkS+x3wjbWcgs2/mpkgUPk08Nhtw+
d4jfobVeTqCjF2aSCWHuC744UmxCiJp3tj+R2opPEldWgDTgUjxCWz4baFVuqDgr
J6/Yk6shaB+1ZGFlw1yjX87TybQ6alRHXQ8B/Hv/N9hlkSzap4UizCv27/tgxygT
pfLPSzGvCW5UIbsQJ2Te+sqG8YNRTUXefnnJIj1RZR5/gsGwY27igD+61FIn3OXo
wsIwPUebw+dA36sm1UqMo8ljPDQUMKb/7dSTkGDZIGU3LOnORrP3D3CDOsPOaRmr
DuuyioY5jyuIKeczZRGprTapweokirRKbqNb4A8UlE/IhbAVs7mfP5IfXwRcKuYo
PUb7y4WQw0RsZ/1TQGMSiuOG5MGJKWp+EckEBekLRKueO9p9F/vWCH5Gf9nESuZN
GybJU70gIimuXSZAi19grkkqkBUZfOO3LXUPE4dUqzHrMD8ISywCQZ/asvmP8MG3
eZ0i68qaMsHzqu5WN70OnOAYyqrWBv0/Ia/HIF28yY/bmrAY5yEoxoT3kLhNwe7f
nOSFo9GlnRl7dIvyVxglpBwbfncToAaKc247iqudyZkBi+A+tAjiniBVQXrpnxW/
P8izvcgoAKtMImj80+fxO7sNWzhdJiK1ttfMP6aFnqJiRBaGUFew1YfaRYj3DKbB
YxUa75JBi1duqe+d8lVPikGFmsUasKgyI5HxF6nF0v0+ninL3pOeCyzpsDZhGSki
MxqlQSeh9dJrlqxP1w5KqtwrdsIzi0G/BbxjDhXguiXDDqMXydl56pdoBOEkuRwq
3ITw1677JJtL39/VGs1B28PTOsakCPcc1BhiNvn03bt1AepZI8cW+x9oI4gNXajf
qIt66dNfINVL58pgoDrLTKNB/zeVJhzclAdlJwflj6gt+8YCL3EuAPm0uoYwQ+dD
MnYnxm1JjZeg89VWf5l2yIaPMfjcbujvMDEqRl2CgWzRlF8th6zKO2L9RyRnpZIt
BzsqFKSTKuhZUXGX39rDTNIhUkVzM9csWO1xx+LF39ZNvBbKg5GLQCrP8fHp2yaa
9Qsg/QXWcIo6wF727dzlbStTd/4Zy+Ob/b0NFjACC8qlHKK7rDqAYjR/XqaYudok
bdzCbzzPW2syGCxeugui6thORbCuWvnnnCSNARC3Mf3oXBaJvDTI3NigtuORksiM
gTW9UxB0j43w0l4uyfYBVrmwXVukWBxLEy+m1g20T+etHq/wlzjau0voSHrvQRec
H1H1IlfC15OEYsGBJg73UgLrK8Scf49XeH8ENTex7nPsF74OiZKY93pOOjAm/qhr
M1Pnq+S3boXkP6bDiZaTtF9dkeh2+ADkrCwGX5M3geaHFK2Ff1dDeI2n7vpr2uXG
oqbl9c4waoBB/3uZdcUcKVyXZrhUXtHn28gh7JXorTho6HHJNHzBMCozZsjZ/zFQ
c2p9kwQ2tzQLOYGUkR409ukoCwt/vmzCuHd4TTNmO8OAxJ70ldL4LwIG3zwi0FUd
cT5J//MWK07poeIyCScorRce3zRYZ/gOZ6dsqQ1rAtmSAB+ECVVkb2EiJLDCd7Qf
Bd9KjY1FCO4DxtQIqaDMZRzRoxSTAluXSe3BiTPJH9JVpBCBWLIAptx7HX0U5VOo
UwQlb3E5LzB6MA/kBMJZhImjBouZdOqNuvoABuiso8fu4Kw7FxXwq7xG9Tqc6P04
XSdfPIcG7lZR3ZoyozLhRHZ0KVAYDoFi0YdimSp7rnMPyd7Ni/6ASSS4WWf3/Lfd
HQSks7rHQ3e1IbrsX6PKih7KmriF889g8u9CbOo3QjPNuqJsvgI+MO2Joy7FRpO0
lgKlrhlWWNv2ya7BqzH9KT2PLnErRLp/K+djkayYm3SJyQYjlvY3mFxfGTfghsas
tdmaN8JHmXuPZBpY/VexmRHYd03KqBI3hJ/2E6mAKZPLH2fPw1XKWuwrLRuNlUeR
RCnZq/iDbEfCq48fQxheMHZdY7/DaShFyrHrvJ7ehkcvhpkUl133uv79CHSsB+Gk
lMt8MJXNractEarfqwcKxoMeeqsQ6dyeklK1bgiHiBlXJodXLad+KbzXMpNOJNfX
QF1UcWx89iCDjG7eOQDaZ4ra5I4kcDP3GmE804HkJ4eQ62Mwfwm9CX9xCim7vskG
+2rBw9RbV7tQOHSJBVIbhD6gmQgW77sMWLNHFuLjGJ/6g/vZ7yld6qwydXBH7yLr
1hwExlqrIkXR1SqTcZdVK1mIhxlzxIr+W5dbuabp6Xj4YsLvugWNOcEVUTsB5kA6
N8A3hGMqgZAuqpbESrmwVnWO1cm9kCMxxN1T9FmuKL+xTJQQ8NmGm+yZbOqg5QaZ
GzQxY+UUaOdJtbccLTFXjrRUXuhD6mfQUhRbrRmW5Wns2LVnf38YEqQjvx5ewmJH
YxmS55AVijD5qGWWCuSwSds8dNgP1IZu3fwzk19U1fHSTroYw4m4gJLa1VaSg6nm
6dyyock24JP73i7SBpbCsJj+qX7ZChSpDW6f/ZDZOAp6Wk4HPKylkySKzpDip6OJ
3p3gVdMApsgWEcPwhXNYLfD7tgQMD0r95z58jSiWg6gktJZVhtHJTNlvxGGP3YYr
PQvckNT6t7ZmqgnIorB9tiZHXESaxWI55LTqWnomLacsqDWHtl0CneNtJXsvsk5B
uWzfgSnf0j3L7yLzxYUnuaajdF6Djy7ncHtcy5sJJb6c6P+ZQSvGsWQ0V9dgqX9P
tEcvHm9y5AKzV/EJq4vT5ZoV5HYuuQOV8isv7heT9w/hedQ0lDe99r4jMzTAleOg
Yx6CeQo1YArYrLHnQfDKNBMdRwRRWdNebuof4QY9kkVhA9tyx5x6SWYKpI7yA4Yo
bQoBMWAE4kvIf/Y5lq2s/B9pw11pm61JDnH9tlKJMJUE+TQVQRd3W4OFiU2xqlST
jRNedMRNPuUbryKkckIFvORUUmEa7zLaN11vg3YLO0ll8MAmIA6DNV7JOcc8sm93
Axw1kYacWkTKjCDH7UMG4CJWFMLQxHbSxPchRHG6tXKkzLKdwRDHjyyXfymVR0E1
pxFmXisjgdBFgJIGQtyXYMB5u+gDDB5nLri2Cgw12Cvvehs6sRJIIXykmgooMKQq
i32yxM3p6MQ2tMePrgXJY2BdBkFwGGlSRPh9t/3SloXiBOhO1eIRBrQ80wfL3EsR
D5Vz0csU442K9SnX9lkuoSelAEinkqlNqoFhSTbDNo4NpmDTCk+ssds6AFR/obN6
bavR4qMPd2xG5IBe0IIKTrKbxpIJafYoF5Gwt1wmAVP7s8hHvWH9jnPzm1lVDXjs
PyhTUWuhytYtk/aQSqypnC26xxCbFBnwixzV67wmFw2gnlOCMtB83B/ASJcRh9uy
AbsRz+E2QcLhdyY5nnBIOILBGsIPebe/8csuLqSOtXQvtddt3OiUjQcYRy7SuuAw
YlKJ3eztIoYk4TXyM+AqAH1RqwJFavobOhdgQxXY6JCgV8EoheQPxEhPI0UpFLLD
XaRoMnXdQBbrCteo0oW/fQ4SjDcZR0iMUoLOo9YBjeYRxDibWpVFJIjchFtEr7fn
TxBluT6+v4Xfb4YXt/ySpsNuzkoGYYeE6HuyXC97gc8mO+3dkmB/2vrDp/g63Lsl
3aSTJLTp6MRu42+v42+nAJW3K0I/xwc/J4Fk1wUmuk29hxSdMN+EK+yqXJyYZX+u
alIQV2gI0IRhp9Bha+4YedO9gane8+nNsdCiU0cXi8JxUW4ZNDI/QwGUlcN0brq4
0fxeNAkiOOBUS11itUpCJOui/FmHYH3xwOumVzp7pYLRYzJIVdBDgxSmEanvxxPc
CnE1CcFRKXOa5CCmx96GO2/xBz81GoQ/Uy7A+mmveS2MysNIld198e7QMOST/ffN
FTru7h8/F5XxfJzmFyVUWbFX9DpBcLClQ06/cMzs0ecJLrfgIX4Wh4Ma2ctjSu2r
RXpQeiAwfVZ8unsgYX9V7U6hVoRrysndMD6horrdACd9DgIVEfwMPmjBDVoNoKaW
EEv8KGDgi936+F0wWxDgkYNBNXiiiqIiaKBFvbnHF+MYkLGjLUS0Tna2jtGypB7a
/TQH6i0Q98Aov8MksrVTRIVaknvGiO2tBl1/rH+CndrfBAZK3MlMnFUTuk2AKwQR
uSFGblK+Vh4Nt31yfgZUkRS1VJL5Y0RIadtSIN3RRC4wBL/UjdvqsWJxzvX0t93o
COvYCDlBRLObEEPDbCzhrxnvomUJvjWEIOM+OHDLmrOckT6F5yr+TeRZToPfk8M1
ScQe1FZTctsw/0V1ZXcATvA8Z2/GpLKZLK5d/OP/Q4Immfoi4HvoDrJhLWL2ilAS
uUUdICmb6WDXA0+G2BinVe7sAKElDtrK6SyngjMoKJ/4FGfG3CPB27plFEXRHTgx
pHpV6mFWDXBO8ZnySdtj8xd1wGiiyxE2RmhaAbmcWo5CvFiOSPqCAd5fJypcaK7x
Vq3nNJPJZY4c805TNKIYPG4VzZslFP3i/fwsIfCKK5FhPNuw1X1a73HjqUO+NbGb
miW+mCUTFWFEUGQtJj8E/sGXPRez79142SBCw8sOH+bb/BHXR2DLoz2KrI6xCZEe
JazYR0YPoaRfecS2Wy4eJJuZ3Zj2kUmjSW0LAzp0bCrG4rz0atjyFIR3hMXV0lKR
5VTyA3vvv7fFFFuoqlZTz1/0JpuN6RvudA7GcOK1ZmZKdDgsSTM9Zbpy0exK7Rgs
aN4VXyhitQF3fjkgmASYAk0GPvKU96qUadY8sxUMHb7p3XvdXLJnqPN5DCtBwhNX
YsSYsoudpnQ9ttgq2Vqjd586DrwCpyFKwiFf89Hs742Q01Xanq0iS7cB412XF01X
66ickCuTjo9zROKBCV3WYcc1trnIusVmgbX1w4dpQv2dnBgAmv5JvWU0L6K8e7NN
3v92OV+nB926tfF6Sp5a2LdTVisUlah1Ip1xuo/O77eJqD6st2jMx/wMwE7RtZ5e
1gtBZjKhsuf9+UvJ2SGLpA+0jQT2I31C9ckaLINAiZHxMrCBXo8wrZkGmpL6iHyp
Jb/IhjxW1/2tgzdQnVoA6a5zXuC0JLzzfK75qjK3NA5oHbQvk5JhbThjrNyY5jIo
SBZqcflV3tx9YCeuYd+YHMp4QdU6Dw3fRjTP2y9uAcK2ey8uK/qd33HpoLZgZKlA
cEyxPh87vZHp8IZiQYpl52RFEzKq3Z76VgAMGh7ot0d0+W2apYsUMSlkGIs1V0vL
ADQWBf7i+K46LrpD13nSTCWU0wVwEkhyKBaclqEpl7KNCRQgMei4r+Ocm/i6NCdB
ZGUjC76XM7KUGWbaoGzZl+paCwYuUYyp6c2lumwUoIVwXMAzP+C6/RcUZzVRybYF
Sa643beBazSTnM36SiXn+5KPNb9Fp9n4eB9PK/wEp04pIDNz4xUvgYSQRFGEqcs0
c+RKwzWRkCKcbLNrJFJm1zyZJXGlRvTXixu668Abqn9SaWXAkI9B6nEJG4A+iUL6
iEKRiG56ytUVTYXzDG2ltmSk/nccky0bM5EYX7It9UA0XxnTECOWYSc9u9u/Zd41
llM7Xi2mgT8ikk9Czfk1TG/5DPPazG3VV7H6qWqELd5yqTlM4a5RLcm9ZYMBTiR0
KCOoebH/cRCRlwRUTNfpM81YvOWkhEnq24OVkfTJfEFEH1wzzuqjraOZxeKJ4DC2
3t7U4D/MNKv3AO18nCbxD72kt0ppt5bOlnGjMfIu+K7varZuUbpMS95hF6XJFcnj
TWDXKI7rDCJhsWJMEJmPH6M2c2N02XuvjYuKgUjQUPlBYRV9qUBfepfQTt/TcuQ0
NuL7JjmXeUoR5lP+nOtHMDSiNdJOsWFfanzZfVJ0YaRs10NGiRtULleP62/KXQ7J
VvuePUm8oE+Y6Tus/dODb4HLfWmfaMeoy/fXiW4Cey1QWXmLFaf0QFudlQqnKa0z
ujKfQIF90cKkBZzlKaogtlseL74KwxPDthXPK4OEnPwrEDhuLyslMYFiO6LZcqLB
yuz9Zp/eL/aF6D1yItVcqSSlXrBTIslqOA6CYnlvPkphhhu55jvN2L0gbd0g7y3q
sfykOnQukPsu/xoKW7qVXiGgUqNHAqi0h2+8XMuTd4/3hm/xLm4JU2oBDw9RNvXN
T+kwK9Ho+j4sfZubPxWkxLnVsjKKEzJDpYE3NvQ/Il0Or27tQ1yOkUZf//8MUd8I
7SW8Ee8yBJS4lWpUFhCusqOE/IiqPwM5TvnHKc9Wj2Zet4IqXHiVRC6tifDUfM/O
EBDEZ5sYyXjsCjz2586YZJdK7Ch+XQkFZbKqY7vGUDqrZzcoZbbAEGIOpp5pH77E
BPfOJA2CAp4bd4HlrbOXuxVVWcIoX8siaX93qBq1WCRxbuV6tLlojd0qyH4rlwQE
cSF02hqitmq2XdQnMzFAai1w52TjL4hBxdhqErQCqf2T9rBgKyQUAwM+ZcoSvV0d
LaBkB966/2jvV52IGYlGbGTTlIvvJPSE/keobjIbTFjeF/EbUbdr7Ri1TGnEsy6U
3mLP35hqIuQZi9HVKgOwwRTmr/38eA6pEWSfE35Pb4yQ7LBTQzbT+iS6ndGQGgFG
IsHiA0t7mHLnWT1C3PMW06LIt+uzuPdDkR0Vd8DtkDV3BndTfQ9ce5fhCWn31lUC
ULmQQTKWdAXTKwqS8TXnUa2E/Nxeex3JtWWB4UumUvnB4zjR1Rq6O2lNe6Wn+mN6
6NoqIowwLMXKmVD9pIz6K3Mywdh7pTiqWLvArsTvLmSlrTQyQTm82LpFlxkKWOV4
hvQFWOQOZYKFe23N+0hT0OP9LYFwh3iEH6QvaMOK6Sd4TMyqyS0XExx7IFacOezj
0x7ySAAYY1DX/PecdHeOqveJNuCRlYbbz8v2EZ400703gEbenyxizaf6cVvy3FHM
8hYnOJSF8MKfFRtQgusndC/W0BMu02H8CLS8PV0DPuJQg5+A4tbzwd+ccyNXuE8E
DPAVH/84CnXYTq0iqINRnS51ntjiAISRIwYrjUryrYlCNxHdq/5FJ14WTP9Nnc9S
t9WWYBMVaHAlh3dcm4LqvhZ0BATOIY+EpK+rs/YNTtm/ZG8NCDfkCB8YJ3xJPzdi
4bVwPhZvdznDGKpoHBgm0UBFE3uOOLV2g7K9H9nqbp1bVvn0hLY7LArERAB82Rk/
9yuKsfxjcJdpWWlNgKkGoFk6jeHpUAt795t+XNg6/BVHCydS6Q8AshG789hVIREA
fJFW+SMfN1NEUiY8H4R791TF0OoTdERITdrYqq+CiqaTyXFb/NKG9kbBW+kmpjU9
6TlHRc55bgRkaLCi30DNXrX4XzUjbL/0PzRoTaGBlwcrykxnTTgMgpr6HThDObCK
MCaTRAIyyO/RdICo5SDVTLklsUWvc97x7/P/7hMs1rbecq8Tw0Q2GXBc2P+mC2kx
4aeSDweC2+9SSsboM1ua+QiAUC9RfcHjGXwTb/owgCsoA/IXwJy47SC6s+S54owx
zhAQ+/AZGw9srqHPw5Lv8qUdcYqqX+0GVppZwuHkze3+fp8w0rHFD1hTiv7C6iu5
AVCPVwmP1eABEs7joFrvXUHMv1QzkDMi/5/beE5fy+yWP2oUMps5Ux23LMpJsaJI
PtmZUz83K39RfCoDAP+W2C4rl+D4PozlQXvRWaLggSCzMs3iFKkXo0IRVNOGAQAD
OOnXCU+7dSbkbNj7tG5MNMnexb4NJF2vw/cAMuu7SrM0flQoCi3TntO8DlWJiz7N
UNLbPIIa8q1ok5tEKY6eYO1KbwtZFtSXlENaXN8yuVvigG9trobyqUxipcDJ4U/h
NkGyvs2DHa6UyfRD2BVgWc1gsNN499N1YG1iJBwixPtxpPCg1Fa9MF3lK2g9cbcj
e7CoVXuSldFVC36a67QkKaxsRyaTBuPpyRO8Oq0R4uxDaOqOd6PrPmsB5JTmv2tm
LBK14x2Y8s+wSE42zboHLS3ghtxe9VMAI+j2jbSyRlzDwsGs5xdn3u+W7YP+KiAm
C60wMTbv55ve0fp6ZOuF98iJwdyrgd9PMtATwgFcmGnspD98uYCx14IhzlFWrW0J
+APpGG2ZgYz+cuBiNS5Bm7/1dwCeJTgpnJr9JJOY/0uYBnC6BrjZ3Zp7DEUD8HFL
lftsnKRBXRJJFtXleftSxZF6257oeEGKKtMQD4lFMxOlxlmCr1ztem1phHpVFBTJ
UeQOS1D4XsqydRb2MIkM+OMAys2O9ArDR+3LhN3Ue61Mycu3G3oKlIj0pXpy6XS5
C2B0gXCyRjaSeOXq9N844XqOADpW1bGTohlpiP9MI/xiSZ3SO1Uto77LeFgGNyP9
DchP7M0wfwHZ2754Rg4FJ1u3zECCeOyOxwkqnsN0adWg9AemDWWuHu5dDWW5tYJo
B8JhHe2MHkTHd/ar5n+hVDrBU43G/TUJp2RSELTGxaQwvWKEJnbVYFFZHQ+qH5sc
BnAZ+DO4D9wxeIij+Ah8nhbo/F/7BkZfZ530UDzIvBepc9n+v2eLBKKI0e3DQqnz
lmOc2uPcrjDIo0QyJsqFZveyHOVRBv4Isk2WwKBCxZwEgeFz3kYS4bOdox5bLR9a
23Rq34rrQZ+sg5HKBH/IfQJ1PibjM4fR/LTcFQIJLlyQw/5UWdFCQCJKN/hJYmi4
6JExO04elOr9wiSPM/4Wvgmpo/SEok0zOdguiuIRvbnF+jrkG7Ub823rgzyZTKVK
qNHxzpd7tuj94zeUzLDEP2GTrzMCzPAL7R88iYuappozI0fHY9Tnys+gynOReoQS
wc6UTyCozln29axsyCBUMWqjpwW2nMwUIaR4kv4fC7YVNkk65bN99mzlFDELLyfS
5xERBHAFfFlGTLAUlVy/l42Yf4olIXT1LtludnAYmnkfugcyyTq0g0hKCk6t9vup
kCuLXzvdvNwfjhVw9YiQ7nLdfOYpmNjGhodZEPRVFaQZtjwHijZAqK4JTmw3iYCJ
dvK1c/F6ugigxPWLZXJNDag7MSfMvH2KunIroXrkAFGwdjyuhcTg0HTYAluQBZOL
TMT4trFw5EJKVOGH/YooS5xbnogBu62ga/yk8zzMDUIwvHLkrjdEqxDom/LDUg56
hK5+TPBqYUzykzp2zEtAmrIJ5iynuM4XW5Ajb0s+VcvktgjA00vvLazmdLx5AfWM
wDL9wVH7cTEv4Ig4XcTHV7TSWJT0wmHqT2WYfLt5mcDGGl2JAvxSqTIBMawf82nV
ksYE1hb0gWZp5bv8RG5fNrsH+aibs9Fn9SRSQXbHdGl53mLPLrqOnECZ9wBWtVru
W6OlqZBA4/wlQ1MCDydlSiz1gPfHnWcMfH2yhrnlho95BpbdJviXVbU6H77H6oSW
XY+sqqcA21sYU2/v659L0DJZiyKYTAqZpsMtSdm5TgwXJpr+D2vtyPazFD1Qhrx9
+wPdwl8kCV2CE/wQQnDet0xEnNjEFgxIQISIxSRWa2dz17Ysx2JG2bsloHJoolSd
v5xPEoLX8ubOGrjtIJyUlAXXCgt5cjfc0G/bYxTLb86rtDoYbluO1QOEoDGqjGQl
Z2+OfwrFNjD8P6dRgZh8YULiFzG1CeWI7sTzRRG7X63KEc2nUyC8Kr96gOMKjTO7
hEflTtAvs+RJojTWdipJGv877pxK1UxKAZGZSCw6SssFojA+l4z8YdHL4r65dYSA
H9IwuIi7apQsvY8y0/pXc0mI3KJQ+zS6VBk7QUqOkvyNHtgzNM60+B1A7fRqF6G1
Vw+AJ6u913X9bTQ4G/fkaDsnjAH1FueOKQ298lZTb9FLspiicmlgZecEd8C7/Wo9
DcEtKAH12RakbM4IwMk6Uskle4kNTxmkyBWconhf5A5xt0DLuAAtLtffRyUHccgo
oPj98SGhWSbxSs/D0V0aa692PtqgCpTSQR1/iGbtppaso9zwvAnAO0x0hqJQxPty
GfeWmB3Mg9FCC2B+5LZj3H61jfb0UDaNeoMT319etxUgEkbaqn2DfhHzBqtKx72j
YGeBAo6py389d7OjHnWm32GnDWd3Ogcz+XnIcgBVznxaMoE+7RieOaOjo7NTL1ok
9xUj5Wwm1bBsbemrM8XToHvMVsQmfb0KwtZzFtI73hS4xmcUBCwQLTLrrC6q5obF
YOs3FF/eSwRszuhPTrtKnYN6uzHjdte0GZbtGERN8IIdngEZ4CCL7bpUGlpQqjK5
vrb9jYTKqKPlpLkcQGAvl7Y10aVXhWXm8TWZWgw3HKQA1/Goah8wny9i2WukZc8H
Q6ub08wWWbg1l8tnHoDmDyJ/aIiojvgowUqLogn/PdUJdjIFW0qY/8Cjs+ok5W0l
zwHu/XL6HiWNmyFR6KOCN5DZ71T6Q7X5pRzijtes6MUKHfZUtewbijgh3IL2pAMI
MiGu/1VWN9pzXEgXMEV6evyNVUOT/eU+JvIXxKLUYaa5rpsOlJFZsG+JlrBE6FOT
Fo70qDCslxzmTItZXcWspISu8Y4a2uUqyrL5xN61l+TjXQBKo4Pe4JjnAfrg7cfl
ULGBUlvfDYPENv8eG0NGZ7Z1ix5NEquFAf5S0U2uvY8Hr6mZN3TqGzLtBCSd1GPx
fSR8Ht/oCpqdP00qPempW0hKqWC6b1fOWiW7wl/U/6xxKuLpkAjLf2XOi9ylHHL8
Mj1UyyI65uMUbiBEebQ25slBw7dcadBE2394h8kJBYLaOsjhMDZhoYypF+NAu/TA
5QdIKsHeCYdzEm5nea2yrlLTA09P4Tp+BGFvZc77C8RdHPV14TSFDWdFc89Bup7/
gX+ddyXp+6C55itkeL81DYA4ur8Kj4uhN660URVp7FwEX0F//DAM/LEAeg7fJlJq
NRuBMJwClQzfKfdPPA1MkQ+ljGHHt0yXlwiOW8hpWG3l9MQgdXkciSBITOFiv5Ms
oYkFfmBcqNWFs7ikGw8Q1R1y/Eoiy/zOmcC1iMMHKtlmCXEnTNfko2IXnHHGEsB2
YYSiwTQR1UZwzylQRwPQxm06JSBTia9jtYG394VRDRFgeLITSk0O6wGR6A9gjg2u
MSfHab8lmpv9PX7tUmzHH3fUkTqP2g+VwpA98NZt09UxUn2OHa2Ek1Mza4hKTFVY
Z8+wvfKOXNd+W1Uqdrmyxh2NBIv5sO2Njg/htpR4WmWWVe0GF+oPgKVnIvLVPj8u
Pq7EmidEMSthuDEgwlw6kGlpg5Of6LdI8dMM67LNeTtfb4xwRsnvrMrgsSPhPJxI
n2c362MN031AYBFJM0uJ7VoUbbpfKkgWv9u3KUE7uxm9SmzcVHPY+iof2+vzSvos
s1prh4rzoUpi5JwfOxJXQePLFTYzMae1F4UVdNTPtnMG9kId/m/9vcFb0D39YOOe
FqwkbPHo1olslpajSgKcQP945szyGxSdbNmn7Irj+IIBZwYYI0yOUfi4Qe1ekpbB
j/FCAQUIcUSamh7husQcyxgbUBB1GR95FYFj6jXbZWShml+VdZ86jZCJcfS0gWFl
FV1nPYcg9Os/Pdw/bf0oEEQIK4SciW25BIVkkxUs2jfzkm403r/IT0lnanUWL27i
c3FWKFyB1F+MhBxlAuUdW36ZpmFdpZin9B1xzxZWch//AbcT5bR6QBUTwB3ZzgYm
t8RbdEjBweQo5agoHKcjGlQy1eU/0bc5gAxRJmaXK/jWizMMDVWqBTyQCWM4A98f
Kdy+IrNHSre+6UeIL5OFSGAuzRB5RhIQvMueWgJBqQ9LwqZkgy41qZkBpVDkCC5r
y3kO1DQiBAOMzuF9BwU9bGAe6qoqeLiluIPTjQrQ/ennc9495nGWL5Cm+jrR9GIc
eyFZgM6emjhFJIvJkZSQGjLwXibbCvYLj778HFrysBij5QsT7kGRdahVJnwfSZ1b
OviTKaSHKMCkJPIGRvzpmtAX6dwtswlDuqAeTzGYxmcmZ34I4slE/pzIqFT44aPL
jS+nWJc+5+DasWptWx2vnZ0MDzRF8JuT+TG06LK44mYLpe67uLDEsf+D8AhxeEek
pDzCZuXAZMbnQbKfT3pVfB8mLl8orzTF3ZSH9p3xQctbacQYR2ddTSfBpSc8q7b0
WqB99ZruEDjWZclXQ2NmKC91FnwvTaONdXsdc7UmTvR72rsosxgfPADKg265zfHs
qbj1RXhoLQoBQJKFbcO5DTQyV4mcvXvdfoqeaq7KVIrt6k1+oWQmQR/MA0Fpx9Tt
rV+yJQ0lJBvbUfyc7wY2e6rczhZAMwF4zpe1sNviC6lSSJQzZC2/T8QR3vv8M2Y5
ldzpWfzuSywQzi9iHRufy1uh+1jlQgLM6ZL+cOg2YYF2WABViIl9Olkprf1AYZXL
6jVYYriUVQ4pDt5LioanuDXH38mCQhh3syV0UxyCRfBMZLRExOX+oVAHEihWvhiB
oiTVbYNH90AH1vKt54vX6aj40TzT24Y2vHq7SqapCsMmTNq9SV1RUoFsSGdFblQj
fTRBg3B/4LnQW7VrIAqvGGOnHXXF8NtLtAKX+rNU8pRxo53CQLhyOZbkIm7uG+ia
tK+xNfbV93uuervKinEVfIVsS1dXmgos4y1iE4cIbHGkgaxnePGbGT7uiRpII5bu
WkfPFfvZ7mZAezKkArdxcWGGekdu9cySBKKNJcQLn7SpH8X4ZNtlg6OsfAumVfo/
utHC7YFbhlpAHSiMOrdNjMgf9nuAXjBWQbahbQ0dLz6COR1/tpNmXlbPWgckD1Wq
VT6RonNfshQguiswlAGyMoqFT0fsILZSXtGSZe4tfC20A822cJ+08bNEyn9M6UJb
ZhsOQOfH63Y5wmO89z2cEeQsjLzzoYvhFqfYEUPenhLkyRASXd40U9om2pE8KhgR
zqSyZ855L4MFMc7fWZqy0Ksn0QaF00n/QesIhIG76//ld+Qx2fjz8cAeLvG5ep5u
yCmwq+bRw4PgGPjufj7vgZ5ET92HDW0/5fBLUhyka+9n8c8yxjkPyVwK+7VGyggx
zdulF2kBuYf4sWEzaZTQs1ZWZZg38y6YReR8ZRk2eXY9YmfozHTHIvaXeCBjY/k0
fYDfo4t0jGo7HjMrEtafZy5CkYlbzs5OGg74wTORX9d9xrnIICarAB008a1mmwqt
I6iSeN9WZzhMAUYygY7xan92GtlkdNUIBDWR0pU2XOu3rao9B7YBLG4zDHn+1I9Z
5x9GyUvxbCaiNkx3i/d/jwJtF+gv97ZpNSqPHyLuFVlndsBz6MVJCUhWZ7hhjOFk
Iz7cW9FCJcfx5ql4baear9cGuf7tq+2ZoXCt5Q91JVV8Lh5U/RGdxGNSkWXoereZ
OMa4BLmoMcbv8X2ZIa5sxiY3DaaBKlqr3MzWh3BTqHErKkMwdZmdIddT7K7KQgGz
iNsYcg2SFUkFc7acP3gaHYtF+bD470e0Rn4ECWo4aLTTydQNka1cWxZqi+Vz+LSW
RYzLeQ1cUA9zoO2f/n6ZFl9pPRMwi9hh03JrxERBRwjg3w5QGIh5C+SK8ErQZxe3
1a65sw0MNQiiBenXEMMnt0YQDnJDzuOqLBLOm7RMidagXA9vlhjrW2l5Y7Xsi32A
GcDrH23B8OF/PsvvefU3GXrDbgPcC/860N8/Dds2d9Py8+Vo1CtKInJex0vWSaft
0iHftfLcsJX0ySDTCigXirafIcPnyChrKeSOM2YBseJplT3R5r6TgD6FKSYe/+Bo
GQsy1oKcWKwZo+UeniAg7aNAOuDETL2UMoGYdJ8je/DCtFCYtwsYzkD/PnuLZ17c
oMnW55NN5Zz6xRid4fxKRbVobzvgKovnbc43rxQ2hZRLVpM2qFWIMrr4h09G8rv1
Y9QglhkyRw/czYvqsmYx7ngZsphIAnPq87qLY2k5Jp/Se9ztXvEAIgIZ0xtNX92Z
JmJh1F9dpL4qQ1UePPhbDmB2AYIrFuZJb/khDwWmczyRweMUmZ4qcVxhgK6Z2SGs
BV9c64IbgkfcB7VRzNTGSkfsxM7fhqBaOMuZjehOpJ2t9llTdyCcPzCNX0NMmGkm
F3OWOpFvRSozq5MkBv4CM9yNy5huD9kkRAylLd8HDBZJkBfxxyGeenRd6XImEshe
NGG7RUAQc0ruVG759yRo80UfE1RRrW4wiMHcNfhWvxwffPQ0xzSCPWIfaC/GPj4o
j/Nvz5bTUfCq4/U6GiPP6XwUw8iQogwqI/0UeyKxk7Spog4KTBjnK0VNoEdIWZx1
1JX6vbNvd8pq5Qk/RBPedDpWeKVwZC+wS55qqd95wN7SsFyB4YTztp+JSo0Ocx6H
M7o4LDAhOYbmZRaG2iRIuDlRo7Dmr1yRMwZ/kc7U8gnv6L/nl0uMfBe/6Jvog2LA
8g+FqdjSFTizNge6mbVwb2SkujGECyBX8yKZpAEOpJ1iYF3R8FC1n5H3Q6yk1QnY
KjLmFB41xNIoM5RRbM+z/RAKtDsQKeub+Ji5M/n2nNL+qQ7NrNmZiIAhGghTk47z
DYRpmDd+5b/k/5jojIkXtN3aUYCNVVnww8QV9EvDCi+6miypXAZnUcenIFtEDHIY
cfNcK15w/sC7ZbwdLv0ygCMGJCr9X1Gjp8xSR2nXzu5UrhRmY6PtStyFDn90CWLj
FZacifxw4WbiLU5pFrZdraNzuv/4pG8RAHh4tExNAKl0bceBu0Y+hS42+IWpKqW1
pTbB4dMhMzaE4J/T/Wqqs9Yzd5OJjOhFEsLgyjT1eZwIxQ2MD9WmgKNATW4atMAX
wyi4iQZwPgOWAQycUD7hmd7Fx5RjUSjUXOwchTXvrgvfzIKE5TbndyshwURoVLVu
SjabZucG+VAek4TrvckDmcHb0Pfir8Sio4LzeGxS/SjjZTEwCnyLjZs9CBQQ0UOK
XhSTpOEsQFbpZZx0oHmd2OllNiXGDxMZ1pWETVciJKtnd1+IBS4wj5VeUnmYRZie
rAQlfhlUC009oE6BxR8i4EkaTGH83BnmnaxRehAR30WVTzBOIxGxshmQMqb7AkaX
G3bAOJmFLw5Ck3AS/XERPeKyKIsSNCEx9xT/PlnpkMdDiXfuC3o15aDKgWRlIBEe
sQdiYKQoJ7aU4ti7rxTiIZXBXek3r5mhyeu0VKekhGSUrhvWhtO9GJKt91FSig6d
WWu0UJE0EHFxo2aMjKOLUuJPUx7QT9KVyv5aV7cKDoDGvkM/zez1dX+VcULESe4r
lg2O0O1xu3mnL/DbtPNt2cXgsi7ihALrJW0YA0bsyxW9JQNfxP7E4kysM/bgBW1M
1hkoQcLCKgqOP+PR2dG9AaN0SNB652jCOPdoUoxRq7FphHNhELbTPFsKy1w6Iq4/
cTngn/fcV+hC+IfKFRfpajcQmS01fc30jCzRjscHBkIsx41rLg0PwfjQgXMiYINT
jgFMd6G7HAjhx8jST3YnjZns3YLzOhXJK+YGpK2Soc4xzP6dyHTXQs0lO54uirhj
Q9hxb971QJMGCrgi4Y9PmBnzafb3el64nlOhJiOpe+WkUYCz2gWfigeNMWEFNgt3
uelrcYOJWbTbZd5B2CgIGoJcdHfqzbfktu+Op4Rw3ibq/gj1NBZPYAbJL4Gf2wRf
nU1hkFtTYpLJjui4MNDgQ27PfoBwo77S5UMvJ9jEPhZxV6yNs4881L6a2lLfIVLy
+3bysUYcYJqmWn5J0A/jq9k1qBbWn3fPLZFTyeUaQMqn4AD7WdUsQyrjyAHcyZZf
FbqC1NYpUS1C2xQYBWYGmPDigSMRAselfOgf622f0V+fnBcuSg0hFjN51GHl87xZ
tVfclWxRC+dhVSHjbDVSJe3IiwUaYO9FauBCLRreK3gOkZwVAbYSs7MrCdceMVGv
MI4wB6N+ve7XCk1wvU6KTdFpU6oWMdqST/bmBK31LNBea3TXvig4iSzt0VSJwrk1
Ag/4z5fyj3BTkYsmFq2ALvtyewFQDp/SWaChqx7Iuv4R11yISjdaKt9h7NIxJ83R
Pb0XOAhZHEtX1Xlu96fLvcmpeeuNPrC3zuPDKKLypIMopJHYXCHvYlz0bqVcn+wX
/JvZKGeEze8DFmNdJHKWhRwQd9Bdf9+J54SEEsjDZEAFoiWGaliT7MX0RD7r2dIC
T5N/zoqoBX8WcYz+BF80v53Z/e0eh72wuKZCxZsIkxcm1oKxAh0vkn99ucXQVYvs
wtAXgqR7NKXdh7F8valBJOAcf1isjElWoXkEBo/DQT6sCdcYUsul1w08fGx1NrVd
Z7qM2eDrdcWSqY/Ag57cKg447/Q+Act19bZr+L33QF4KOm/wLuN/l4NRdlwyrWiX
kKtmW7SDV5B6Ivj8ui8itra5zrGz4Pmbh2Q/Bl5qQCBxe2ixUTiWVgcqcBQGJi8K
Rf2Ig3n/dA9MDKTgjWf42uxJ2Pp4jrvMEnNKLvwvYILorOK1PSb+7F4hb3cRiZwD
czbYSHghNL0uuzQ3x1SRKZSbqUWoC/cQuVNVM/bOUuhHFoTrDxFYTnL+yiRnEk3i
QA5vTthbDkrTiMrpJNy5g3TEU6s1G31oyqppV2Apm/St5m+5z/FH3vGSKMRjTuBb
PrwNQWcb9lXoPNKsENkXvzXqD+Q/R5uY4Kznv8miVby3HbymjbXLsP6PBykg+9Vn
+/RVsRPdhOueq4ohbPJCBqOg659tj5aAQ9gTTDzcfZEo2bM/yWcRM3ITGTq1TAAm
U9HxF/f0/2R4XFp+rr6H2EgSe+k059AbonSfIE9Abf+F7esG8pvHzoxLcGrnJJha
QBN8wipjX6pNpO7OxuzUHl3/joKkl18tbih3+ApQ8LlkCviIVlBCPH+JNU/ftUIY
wAJQ3HF+F6CB0xv+4x7J/FWaw0NzyUYRmwTtzYzBBPvaJgah1tcfDekJ0/4YTryX
xZujXmANbF/fG0+y75IYzDdf1Brg3iGELUypTxTTX86qvnfisIfdkEVJlCxFh2HI
o9jGZT9hb+E5b+HtJKEatacXYGDVCSzdfJrhoH7GUgYHeAGjFTCWahGMjNsY6c20
CTJKJrXI3mqtz/YQtCF8ACO0oX1I2iK/IHFNpnl4zW96f4HilJdvaMxdmN3FD6/o
dNZGWrebwn1I6lXBzXhsLD1ayw1JJrDzkwZ4p+C+j8pKkwNMlGudxDZf0w+DvKx3
JSICj7RdUMAIiwqaX/fYBmofMbNIeiRsQup49g+uPl82KcDFI6hpWwv6+UzaPjpW
J9I4ZOub5uvnMEn1DnddJULd5mpym9v/BHK73oA86EAFYjQ3D+qQguoOoKGE1qs6
uuGh2Ypa3yAy09fFBGNBSW4zceBD6DjH3RUyeqynRmgU27JoTcU4tabTkqnN4rc5
lOvlIk8hz8qosfrRh7cKnfePprFBjUM9bcslkC6cv4otmvnNiCl9Y+jJq7O+m5Ya
nodpPeGbFuv6bezfTjMF3hb4HtbfftJeLrL1OK/Q+fDGLeOOMIBnCzGAVUakNa1r
P3mUeUh3Mf7F/u4HZNCK4NB8OludTSvcXjo3aoKruLAy5q2eWiInqWPYX9UcILpK
FoPTJJFXnIqmgCVXwTrFlWsCTjgn+Cz9CinmlHMkFZNMGIZQQJqSrocMtSl94WLG
pKPLy93EJAR3fc8+KQ6Ci8GvEjGDjBeq2IyF2R27muilpBuIdqhPA/SO591g6axe
3xb3gsGyXKlbfV3QXC3ZCnPtWD4PqoM03FVECDZ1y5AHsqNv/XU7hkxDAnTPEk+Q
UfrQT30IWppgRhT8o9mATSJyYLX8gAhnqpnK9bfqyAbFxTPdINzYIWGAz8cJ14Ac
vaSplc/juyqJJWoPFfCdmgFcR+oSOvEDYGbJPIHcOlvPfVT8dju+CQyaP3m2Gngn
IzrHXWxwiMwNpTTJ7YimE+KO44VmC7D91+ls6eNnkGS22b7JkA+9q7Q9nu53w3+4
iMjqAo7IzAmScUenGS269LWtmWkoUZ25vMVk1pIc7foQS2r1xOjOpOzUWWWwJVl2
Rpen9uYbT8GDdYKrqSWn3U0cbIMdnAPqOx1/vpS5JIdCPWjST4MVQvdIgTcMYvwK
c81ULMYqCFwBt6eJjbUwGum28iUN1XrEJJSZHCrnzYdz86xgI9vIz3J4cunGuCSR
czabby6WSCf6Qf2gsuQqJ6AwnMCIq7ty6/WA7XOuoh3TxMk6MLYryXomhLP+y2e2
Xf5hBdxkaL5q5cNizlHAiJ7Ikw1bOtatXqEDVdwMN5xqBVnqVJeLffVoqWUFEySn
ho3DT1Si41i+1zhUxYZUtpx6QCsyIgnjpDZTadt7yzpNGVFfJJfIxd+UD76K5vYt
du+Q2FRq/6QkELr9ssY5OqrnaPHNvHZBwverlUjogF/LW5Zn3/N9u+9vJPs3poGU
mSqhDGiQKQJqx5T5UQGEe4Izn3tfBI/H8BO1v0lIZ8YDd6NbHpNIe0B/e6eRzPE2
yQa4W2ine1xM9+p6Ms4eLGkAtAt/0G1U9n6x9ywUWLUYsASsqI4sCZe9gAOcNuhe
d4bPz7lYu+nxpO5NWzjVpgGzuSsC3UpmEb6VQsH8HTLqOzEMvTA3dXnZ1uF76Hj4
F6y8EXi4O8xI8KU6qwqptBtrbN1bN1XRH6OeLEdLV6XtXnpzhRTCAlvL67IAYbbV
uOtPwhxtGN+HMV9z5GiVULE+hSF7kHtI749u+bn3o9pWEkxSrTMNXFFymqvL7hpR
MXwq0tBWSKR2u0GzB6DBgREOjZySgbs9f5ci6oErhC/RUwfDZYON/VYedcPPZWih
k8rv594q6CQni+jclOhqxnAgwr2jRR7QVbkU2KxzFTQPMLXTIs0ybZyq3Qa3qcz7
PTVbXcPwM+tWYA+pGAJJv4BqH93bFZykQY3uxO1Yufk/UwoaPMEs+zuD+/IYMfRL
Tengk/sLAh7II7F/bj49zFVvi1qcx/iAoHN9bT2BxSwDWZiInTKpKHFECk+BJRAZ
eNXKL/Y3p/ETk+tNZkQz6GALq+tIH7m9FvhuF6dKD1uEvGO8CyHD0b5icaRJRpXW
IdgJfGINhQOI+6SEXPaQUO9Z9f9IyLNcUBLftTC+Qj3JzxKFz8U8lSFyoJhGzD0K
8ke58jU20ZkhHcH0Zx5bbsJ3xTX+Mk5CUUXgcCGNLaEqpBovej+tqwDrBv4SqqQb
z+bjGy0Lx9dWiudipWmUF+cp6k6ye3xdS6t5wbtBpqb2GHtvuLBE/3wUyj+4b1aq
Si4tZZto+ZQ/Sj0hYM9LAhny846025Epsgpfsom9UyuRU9kJSmtzOZHGcGBR3yuC
KiVnNA3FIyqnu0rPgRk+gk5X+LjeXSP1Etkgv0U5MVh4hQJ3MlDqAa5UIwaXgLpS
dfFn6TleimQLpow5n+USar8bXd/9YyOAwNZHJWqK8QDWdAtyQUtadu+A17Vw95X7
ZSUQVl0BEnaIISGbFRQQ32xPjm1a9RuGnZClL01W3998Ij6DgKWfOLtpI55RpMZY
z4WpzeQYwQ3NqGyNCDXiEN3kXzJE2S8Zl+1xSg6+Sp4+zRptYcqD4s6DE5PGag+d
WP+M30aIuTU/r7p9PvOZvcJKfvU7r0X7enETzA6yn9HDaKVYeAP17Y3AitJMr1TJ
3CQqRLi3rkfuiGk1rn7AL6Q29Imd8XJy5UL3uooACCQxaFYSoQJtkMO7i+yJv8VW
n6ANXmFxbInxNmXf8mQKwDjWtF8r0YMzbAMuFPya6kSaHLDW5Oolt6D5SiwZ5Boa
rZLp1zPcMBXi9FNk1oqrmU1Ov+N+UKcRwQaea/Sa/pPl0bdM0ZDPg7g7qntPDpg5
XXmrgpcmNmJ4XUt3jwhV/6uNJdJ25XFWNr5FnHOMlNBmAfWjh2RKCeM5lYJyVXg+
TBPsXDUk57ywXT/Pm63poPu/3hLFLMqROiCQLPBlL5gMy9zOLhWhImhyVH+Z0Txe
o1lxxmiDSnI9xS7Xl3UY5ufA6Y1eFKAgUHl3vr0SMX8bhW40SaOzWMFl4ib5JfHM
G/cZlMXqF9vitCQkzMmHOpoSa5QCdlT3Xw9SWs+wVoHpTwpHYkhXi6xpFNYU2xc1
SNIlObxbWB0x4b7+KJOpN4smLYLvLR/lj3mF9w5k+6IHlsUU4S5/N0nCw+0dBm12
Q9EHQqfBujeADlyPzJM7j+rPz24RVJMb2PN0a3M83dLjLevfE8e8v73Ztcbw5Rxr
hurQac62hixhTV33uDj1Z27vq6gkh7eNL3Phtwo99xr3qhhzDbqt36un8C77znEO
/vQBtcVH3rcgt54piYC3oWEh43OotZVFWIUvJDJ9Wmn9bLGzzdHXnN0yXIiz5yoH
EL+ttyQkuSb8DybjOwgplr34jurBXsd2QzTz4ydbmaaoR62EozpI5mLXtaWFSG3Z
r/b+V5+HeEFFiflJP9tr28wWynObOn9w6ZrityYqIUosR8qJkfmzoqxmkL+JhvKl
WHrHCUAPVgiscB6/DpMgWIcP0S7GT9KqsUw4rq1kPMbPFW62G3pcOLz8yvIYplZL
Pis8eOsA1Q4wc8BNlOgEgmrKXFd5By5DiMvSlvFgCY/s9Bz3/qMRf/DQm4Z3LiqU
whTAu7IgYkB4+Nc7AiD7tIC1tPeKhb+j5FULFs2OLq8riKPXSJ0sB1p39BkxgKJ6
F0+H50mK0nBQ9C5Tun8lnzOUkvKoAJbW0grC7U42mUN5qNWfQcNLeM7OB9ZjlJKY
QVyIwQbZj8gvxAeHPd3Y8vf+/M4BZps2ebknSIzvuT99FCvFWy9RWwv+VYD1fSJa
sAlMmOJ+BwGQlLtYKwv0urUBBUWJi0GB0L+RU9XpGZLt3VCLYYTLSvRJeKelaY/k
HjRLBZVcKJaWBNIeqj2Jv21CgEBSlwvw4y7eQyyS6WQuqFv2jwHhJUAg2VncN8px
NP38euPxcVxnMgxIp5Rs3a/KU8Ml+Z9X7iSl3doAL82wAJsMSvCnskmSH26StH4Q
TGoqcz+9ly/ID43WY0cSHBzjYe/2xD9jWAXFqjo2Q1dekce+8rV/momBQ7aliXJK
EzZy/r3Ly14nK2MjFOpOGgctpVpN/xFggLNPSIg/6AVH8dyHUfY376dzJG+X4KGm
P8u22MiHWhuxsIygxmLh99IUKF/pruhOVipP/pkwAj854CYBhnTQgzMclecG5rS6
fs1GUPwgWvWqR1mcnN8VJizlHyZMz5NE9dgT6oEuQynQ8rQUOCDCrWTZ4t9xLKbQ
TCkitUEqK0BIY3OUNUyNlW5igypvILTF4x2eMg71FDxsR6F2+qGYcvzjV9dJ9GMu
IP0Rewpa2Y/DR6LpE3ce1FeF7aJ9EtWL1QXNWzPDhoe9xsaE9ssvKWcKQ6MMBxGK
vaJtUDdwCUwYpBNjZDggqxJ79IvZboWuYT/uXXEI0WaWlVqgXmLXEyt5vvRIFlVF
bn1NMO7UXtfdmSviJklVXNFDkuUSb9r9C0WiaaR54bT9opS6vfnbw83VlyuyMOK5
6zkTPyp37MSZsiRd/92WnyLLsncBYAtj43+i3qrd9JyLJQNx/Db8YE/l1h9Z7157
3KlwxOvvNb/Z/t/PxWn8w0CBPgfYRIi1hH6PMdL14DzFaGjGrV+HHkDoBg7gRcli
J3C6EId+a7r/QjdOyEBV1Vfc2jtq6KlDMqSmjmF+DQ5Tf2BG6mJuhsByng76xzvE
3V2CPisiXNUISuJmPN9vA/2YnEvrSEH9jJDejftS+jBIsUPLc8FqePnVFxL8FJIm
xNCZuJ/4dfF81DcoXe1b+DpP76GE5NgZrRzhiWVIU+d1kXfC6huWV68YrPixo3ue
0UfLexj1BG7JgF59Jmdqwh+x+eSTvrBr+tFlUz8Zocw5MuNrDBwWTZqJYToXyhTj
Axia/tqhY6HWlFI75Yk3gueKLENDC8FbtQcNygOALcPUNE5x4dCtj2ocSzSnYqGw
dmA5WIOgLun2G5Putp5SwKpYSECxpNGxQCAjluHHFKrTaP8wffBu9tb0IHZfA9I/
+v223WWLYJcpbjg6DVxlbrMJc4R+ABsiqONyxe2Vqtb9dv28S0PG2YqpDwNUfSTi
JtodTmMZHXe+XlEJ9WEb99tWVpBg2LjoF8/b6puRS5Txx+Qsmr8j3J8eUBQ782B3
XTuhPa5objYrT6TS6H/aGr/UGcBX4U+B5/VaHwYxjqI8ZR6kgX05/i+Xx/x6yUEp
sCMQkREczM+vVuWxtESYU/jYdMo+BmUUq/RuvQ6X7YBI1mQwVVkCFFA3c1VaZHnQ
siktHIHz5Mf0ANTZCQe0XQH7X3MEo8sCX4S0FqfBW5CplZe53MwDOWhL3c0H2T7g
R6vB0cKlIMpmso5ZvKyKInOrazzgSqa4lICY2N+ghV71jxW5xlg1HzYT6Q+jRNDW
spYuPwrds862Cz7a6ofl9f9l6EZDy5LEJBGEL+rUfqWeK+PTj90YvQgJs3K5yujB
NHYRnmT76e7hIK+YnBfVwWM9g2Tk5ghksQNnANEWihMm8+5d+LpFPsgXoCwSb9Yr
6GMndjQby80zM9sHQwkz14hN9GEozGec2Kz1MhrnRt0r355XTHqeAoA02SSFE+Y+
KIKzfEP2+F7rvmAJIJczm2kY1bPc4phWEeopNukOVnC3DzUKutZItVdxDwVM1fnw
TlbW+pJk01o2RAdB4ltLXxiuIkVV3lZuhth5TNSIiOJusabwTXJsEVfplMD8rUlK
wVcuQQ9Xnp4PkNRPxw/K0qq4+V5pVNnO08WMlzMMQkY4UET1erLZTh4swtxFcpZb
2JnIFlfTp8uuYvs47PSLCk5sdxwLRvH0uPn7wJhysbohS1Kl2nKGLv19ydqNWb73
UuoTqcF5H4JqRzYVnyHfZxMlZ1HJL6TvUi5vo5KrqAgSyu9real+rnvmnGT638hC
Ne4hmqiheCfCEeguPIpBs4hdDa8/2XxqRn3P+yhCPdKLYao4Ijz4AWS/5RbbxxvX
ScjvcxZBKyNw2aPK3a2EJWQULbB72r8ul327R2UVo6x2zjyYiePtn2775Ds0PFWd
GTB/Hmh624NKS2juXeUaLhfIseqmJTIpQBh2TKtAauO0iZo9XVKEXWB/SR45/+Bb
ubURol2lijyvhgb79RLNvmlvSBQWhzY1hrlcZV2dtqPoA56Oi7OyzEeN/it1BlbP
ALeCD4g2l9l9GZJFPBwbygCh9DM7ltEiAJO2IE0MI+JFu1N+BHGi9RAY2fgWVfHw
QVGKL8YB51JkOKbb8Eej3eJkA4cOJXBCA3SLGgW6HN6kAr7h/tBSFoAaJjyBxiYr
CmFfg4trJhetQeqMNGJYirSdvn3cFYvQbQNU5iI0x5BLdFc/ga8kpInTaby7R0cY
48go/O/Aw+oMjWwPlwZTc9zP0oYbUgnDVNrRKGD+iNvHWBbmVnM27dIqI8yyLkdr
U95D8H3jLK9kIl7a4oe79Ssfb+0T3vAM+9ocw5NkPXE23u/Hnq4KiyzvLbTz9sgT
6jpQuJef8sTg7KXAT4HCGGtHX3UDeHN9n9aoaeHx4mwnTkdCgXxy0soNR57Yjtyt
DS9EudoV0Z/So25JpDGMcWZu8a3PYf28Rspxrcn09/Ri/mt+JhFaj0AqD73+dohS
joGDZAXCvq5qQ6pJ/cw7163kY3EHU9VhP6CQsP1URUMDtAQZucRxD1tWI8uqMrKS
khg5QkkkoxliQPMRgzNAQ8FUmKsvI0KB8sTct0jNxS92FiQ9T3hontuuzGrsF/rv
a+qJG0pI2TGJ5ljvbeSX0/bfRV4FsX28no+gC7KMnM7R+fwLC4DzJnDTjO+xW7Ix
nuAFuGhjpG2uQCBhfqfPopwySa7zaVczBoHaIVmOMnW5P0YlbRIt8qXmahPUmHmw
kEvqrUpfvakSmIFiKNsaW3DuHnMWSdwU1Kc5Le3W3Tk3/TBKG8+scvrWDFE0UAWt
9CSSo07pgzEndduDZrY5WowkhHOk+6X5a2nHMSzuktcRGaXksKYV2gsr5OhJjYfX
YBzXQZAPT96gj45H9Ahwmvtaiw5vGYKd/zbrl8kl9b8WzVRMC9Sh6rfz6ivltbKd
/OPc87bGrRhTn+RxwdXM9J3IIPo7nAZUbkj0P1TnfnzcFf6zkX63b0dmCkC69AJ5
kQlyPwg8tPCSgDDaHmXrFqsAVdcfuwGdRZu992FzHumZa/Ru/si3FwiycbfoBF5T
uwu4hTLsP4dx6Jt90+9RQBFxerRGppJMKsF9n6J/0wxc42Ii8tuPhzkt1WAvHcPS
CZbOVoyIj3/zq7uwV8n65K4AxGe3n4+pLKoxeo3Qgeuo+vvZk6BthFEt3e3QSQy/
JEgvQaBEt2zfE7Jz9BfcGNp5gdvODZBsw175yOraCYX5OhfpMynLLU1CPugcbQ2+
GJOJG5wO+38cEOH8W0akb6UyVYxhtiglgySUfgs+5ST3K3RM9QvlPjzVDMml2Irl
d1WPDc1cUVac2OkasyHF83+9EruO20VF9cgL8cdd8dwfUZ2OP8excYPBlvjlRVYu
FpbjWHx7RvF5Al++y6NoAaJMAJW48SaiPHQOOB2yvqXYEJvPXKXb2hELvL2+3T+D
bKr9hbm8i8+xvMpwI6Lk+kQklt0n8jaXSJqWdzz1djOINErpSpPgYfoTn7dizImf
L7Vm70Fy1BOHkTTQmYZfTO/292xaVxZfja8w63aPqEjsMTPPg+Wqbo1UZGCfKEkI
HJJLKzvE7FbQLdikjUQuloK50ufKcJZDleNUYKZmHBe3yYoUtiiwdSSaQ6O9DLll
YIUKIXVd97meCV1VZaoeep/e6Z1Gmg1oKxYxIPFn23IzlmimFRNjbQCyEeZJWJMo
A5jrLRhQPxrvh3fp8hiDSiaKd157g6f3lIFojjv6iWiB6ODM9LbRke3+gbXks/Gg
j1p887JFSKrAd1OLp3dk7SsscI67tILbPv5NiF0F1ylqdxhhH/8JJ23ZqPq2qyqF
isXOnPygyWVdNbjDVqc9jk0mAL0ZNNJ8/7N9Lt3TUXGSHTwYoyUab03B62/jfKrP
E+emXK2xuu+6NzkMCmlPDoqmrf1P+KYPDd39tv+1yG3VXyxwsSfZLtPeBDXvhfZ2
Jws/VTGvRFo2aq89aKUZmKLaD9s4OYsTtxo3WJ88DG3W3Gqr4PcvXP/gyJTcezfO
H0A9AidXOGqG8i+WvdSvc3mh5saXQfwJsp2WlxO2t3pHjlZsGbeBzlWaBcqZ5TrT
2bioBu0a1YcVm4VvHwmG0r9Uk+dEhF/o6lgADnDvJirlNyTRu5F/COu0xdNpTQDT
a2MhJqWh0le5yQkcrw97uBbtTZJVP01QQKMzmw6quIw8isNu3mRG+3FMWEhMzZzm
uB6hKIrX5eeDpsue4/8ADPnKxbcrhRE6xw7lhcGrkPmkP/xbW/V/NNXOncHpD4U7
NR/9GNyRzOU5cco0wR8khqlahwEduATjAQFno9LfO9qja412Tl8ezqEYCgSuMl4B
Cn6UYBojGhXilLJab/VAjzM40GQDEfeOCAX684VqLTpUoSxHAvUEklyTuNXMSQgD
eNlZYOX94ENuP07e2KEp3dGYK4mRdxnjwOxW7MGl1iiVNts0xE72JbZnC4GZjQiN
AJdR/h1/rOLwh9ZR1A0c9etsmwXl4aB13iXzlxayW9tcQY/mbQfNqqvR0PIfL7oX
IJogPbchU2uGFRfQCnhMXNmpo2Rr49hD0eI7A/uFDvJqhPAhDvWcJjEkpviX4Ch/
KD+Eu2YSV6mSy5+sxAGJw4ntVFYVkNw0yG9eAMHHnf/V6UirmQpYz48vm3Cc/H+T
vJWjcWEkN2MW3QLf2/W7xXpZrdbGExBMoCtuybaYLvvtJrokGvTg63U20lTx6+nU
Mk4Xztn8yDipB5VRhVcE2J5ce1fkNhCJgthYCPktqBiX8xFVFGU0pD8AuAM44BM3
0gGXV8tQDA+P4vZVIXwU/mCma7QyfHTuDwrU2uNOvxgorIxYquPLth++me+r7f+1
qbeAfab118iDMU4ZTv4Doa8jJXIGjURPDaEh8wstefaWhjvYf+DEZsm5H7iWpLrQ
L+JWATYnTc+/2LlkC8zWqZHfdsHk/J1b3d3NRg4ft285pHLWYdK25PID05/VItlR
rz7lXSClJy54eUpjx2VPoRsLipcDymDadKLusN5hJH8MXzz2arc7mImABIEjeF6S
Okjc5WZaClOkKfuO72WNlftZcvcRQSsAkxsSzyaEeo1HzVYiV0IfuQYmdAJj8+E1
kWlN6X9XjQTk8lc3KKMaMQ97q2xRhPk0ObilZD0taLywgtB8cOU5leQJKSdMwoV0
AILG54i7aZDz67EhGeAilhzOOM0FBNRMu7QiJ81jSi7zk0Q5D23jcFiWsIgPTSWH
5GurfUybMcRvAz/N0+l7zHlsDGcK2vr8qgTHWqWCKxCNQF8HVEqL9wN617HEscfj
30tINXw1yNIC6K3UcztP9ow/bqFAxTrO1F5v6OdYDm5zkMPoC9/RdFNWjas2Iip7
B0X9I4EPg4MKlpAq6fdC1Qxqfb04S0S0YtRMIbMCXCJllIX054sK4B/EjIUtVFIB
0JhnqwI47vCZRlH86nFL0QUfhrJn3RbqBr/n2qa/y/gtJM/8EnCqtZ/T9vG0FQ6l
Ev571lKw69KdMfiJUFK4PNrH45H/XT4CVaMM1fU299pTqGSXSoJRHE75nezH//W+
QPs7k/Il8i/RmHAITnU45FBjkN9wc6Zl20C3dOPief/CFGBQgxEz6Xh7KffPyaBn
Opk8NRwOUzyib1GOPPgeL85fQzx+REUwpyJInUo0LWxxbZ2pFGXVrlnYrlMKHiCM
CHTzoWirWUeZ+tgSy14DM0L4bnd6fv4zEk/7b8gPEM7oqQb6aVsJtbElSyr1bTG6
hhDUSV6MsUbaOKYH5NsYbBesc1IA7HuUcQu6zMbGH0VI5XdMAXT+ZqKanegI2wjX
Z5wZ+6gQqoU8GZ4Gpx12VxHvQhDQ95e4+c0FLzjHsmmKMnDDcxMhT66NiYf5ynLg
el9SJ7TH+ZnNTJwMD5LrddItqZ6JrtH1M2DzwxIiaPBi47LiKJr4pK93/7DNMwFP
pylmd6d5ZAQ/Qax1HA0xq+hkuJ+Z2fzADR3KGgxU2ufr+mQVsOAvIhOP81Ze7CGV
eOXTKOHGPPa8DUrUcq71zS6Ij2PGS15yMTQBrenFvFD9/zM7/mbjhBDwlwhxSuYj
MeRe/IV3kKLMydqYbsN2EhGpfdBNqtpfX7EPtnqIF/1SjqvaqyjwxpSmjaeOupav
Y1spypV7CrgeJLCs30YZwGdP3yNkv/uJAQiMaFDMGlAv9bfeSJwx4TqSaCbKRUu8
QECsOfbsrwLCB4wSNB44sVpukM/54RKn7PSRjOvlB+w/hKUSdsWDJnPAiR2aBIRb
URpwlgiUxup/v10wS71EKz5K+Onzl5HtOKgBswYMgUT+s6EpDnYGwW74ayQv8D+6
i+NFT+V2Bd+y5bGDWGu0/don3p/ixZ5s36uh9RTyzGHGXqwH2WoDCNqKybRCYaEu
MmzXmgrFJP0ll9qOikShHK4dFgBZ1+eV58g9c0Z0fLl1skcpdsaQGe4ffKgyYY0t
KzypeMQhPuLxWRljdKywmhAR4hPSCiE/s+BxIMMr7vRkhTiqyGJhFBXaUArnC1ga
qVL+OEBbFsMk0OWh3Ez+tW3YtJusOYMDSRu6AfJkxjgWbQ5bc1DNwAF9uNUwvTXN
mq2VHI3i8cmukfVNg9fwhfflLe2Fna34XcSzWDmOgQe+yNalxlniixXmgSMI9POV
uK6Bo0WQPvcietCe+MgF7cUHKwiPi4HyMDuBNszmzIFwUeEm2N1c54QDlSaxkWv6
PGxABtUTC6uYGjI8mEC2gluRN1YaLEoD+ZM+2f5xUTNFNt3n8BAyV1pRs58LKdfs
bmSjR8oKODwzSZN7emGINF6lox6Y/GU3Knbp5DWpISWAU/RW6b9FEIaOqj81I+YG
mHri3+XcT61eSHtB/GZtaMxLiXhWwRiOOv5MYVe1G9Q3nwro1LFCkbxuBtVVtpgK
D92pV9iVXpuG5R2BQfOld8lXX9mYCWgEl32EdZzr35BELcHveUBa25ZS9NIG87kh
22f9+R0Za0+wQ8teHU6vccai5bDc3v/mPXGtrAPBxTtWcQdtHUDjbsfNVU2fwDxk
MV7wqKIIj8MOjhHSXRbTvrcVIFDC51E4KQgoBa9qsgp8a3h/6xvJlCSOMS/3ta1z
YuqAuC/M7ucm4J0knlTZyv5uGW5Mna6A3mv0Ups/BIJ4avkWFOlnfAldxed6Q2YC
JVaU6ctU8jBRyn3u035djgmcFpUtRnENkxXLwndolYh6ID1Oy8R01hDLrzjuykDx
OksO96RqfhjeH9Zc5MC2Ruzrq6WWnDF5M2AnaS+ET6x1zURfhHAWYaLCn4C7nYxg
3OABgzo9dF9+XZWnusP7s8bnp3hWCSiSQqYE81QJAtjL0AjJuRokXuMcgqn7kIC1
6KWZFI5RlcR+dqIzagnXQSJML/yXHmTQPizOkMdX2BsPhzMbPxpNK8XhbfUU+IRg
/bTnt5Al8ciJDgLF1klydR+DEggLhXkE86mswZ+FXt9aLsDTZbbjsTTPGFgwApzS
jjv6naeoybvzsyWS8PA7J839fn3HCV0QK+Z5ZQti0ucLOos5VQjYf437CHTwd+EA
QkDP3nvnNGZ0k1CcNUQDLf7jtOIvCYJ/AcWfWHJwa+d4SyhbGszd0vu14UsKR6Wb
iHk/sJ8V6ENUDJDzjIht3dMFTlXPdlbutrLtvTm0oXclKU8ZRZwSOWVD4FGPIXk6
y87Kbp7+rDJoQlnCz/n9g5CaGal+0FwOyPFdzTvlV2fqHOj8Mmbo5p2LqZno8SRi
C0X0w6mdsvktg8PvqqO9TJu9fI6PJHipxJGHDvLq4qcwYaEJ/jttkthvVkQGls7V
+1Q2P6m3iVfV9nx74I86cXlwdn4G/SV1X6aZ1zz0tE0ETC+ok72u1/yl6YXKl21b
kF8kQHwRmgv1JRPJwOu5f7ymG1f7FIHsKQICwpjeI8a6cWNwZp9MvgQGfR/jNv1E
0aDhKa2TnNPRxk1EoTFW4foQlJhHHkMBVVQazqhKOdu5EUohxk4pVCDsjreErvtJ
P1DJHgf+TUf14+AvDRS9F7xWV+GtyvT0qGwNrl9XdwfZvTe504X1ty/SLdIHOtWk
i4T4kdsOQ5svHB4m47LMsIryKfZqQP9h7SxhHaFtnlysQbuRK8+Oal/GUg5HSd4V
bC5IwEhvM5iA2bRiIyz1GReiMSDX3aPYH8w1eR00HpXIkzVJ/u2QMLSzSBxfqEIB
SQVQJ+Wjz60/LAckUXpEeXJj5JkfvmC10rlo9+2HXJlirlcfE8igDwjpkUkxxq/U
3D6C0U2q20MNgCgsTcWT1rCkOwXY+UsqWyklNIDvKOYrXIAOKgizBpu5mBxb8pBA
wtLGk2NhDKuwgNz7U1skoGaPkle0o8Z8KE9WsRVvG96YKCyUQCwJ339Xr3U7j0jM
eCEGZKug4MJ1PdmZhC8S581D7oFSPpUHQQknpphuyiYlOEbW5COPzhXBUXVFq9c/
rOhJmT1THBczYr2RPE8bK+uWFTDvJzgXuPWLGKLYyuASM6EoDbGLGH8ZZPSKOwys
q/qYZE0+8pyOavUorBL+saNwttMxWNOTPLuGJpPJv/OP2Et+pxj9Rv23/ESzmm4g
PMysPhmqoWW0uEhSw59Sv/dc7OkXemTpfXLMq8Giyma2XG20flvwrWvo7qFrnKI3
lRddqCowOLIDdA1C2ja1DzA9t7fE4BOnKOeJaUwomsHc8LuTxtCVqHb9FW0Q5And
s2GP7uRkeB9roYE1Z/R6SxfL8z/Eu4ZCaZSBpaOdBbxgTDRzDg0J7QPkt/Zknglw
/LECmSO+3ctM9iQeZWhGiZeqsW5yykrSoyADSuXSeL9cNK9I8H2KG172lcLvgGhg
pzzPRCwaGruD66+Kvq8sXE9JuWbHp1DZ4iEjpLqDjJasZrG7On7KAiTmCv80tMWR
LucRwP0xzR9k8v6wPkCbbY/TES/f/StG71u0W/V0Lqat+14fiMtMcBOzhpabpMGE
sVrfSUpOnuGR0ucIFMU5CIr6YMTd+K7E3Xj6dBvax53W/cEzFvR4fIjf95dGQdiT
JstZvPTGnFVHm+USL60pPkH/gB7R6ntny0udY8kH6aCX9OUuoa1ynojTqgiU4IBA
2XdZV07Ly5UgOQ718OvtP7Tmqlf9JsAqyiay2uFCoJbrZ+ImGQsnLuXG3eJxZcN8
wKUbwHNVDQ1VdEkUZz31pm/BV6TPYwjqvCGp6fVNmOo/YL8KXbRPS9MW3LIxhbcV
B2LkT1KjfyEluuEki07r6x0biFi/LNg1akX8Oqbt5vh3ScUghTGjc7MB7Z1uQhm2
GE3nk3rX1lDx+Ytek1Hl9ak5A3aAg5SoEhWEcR76XnFgXx0QN014bgumF1h1U4Yy
iJZbmRlz6nxDmWEJdRFUPU6YdQB3Y9MK59/v2bgf00ZdfQDVEglSzTeM2UXC0GMw
QW50AbhnEp0jh+q9cn4y8knq7zlD7et/j7qo4wxrMtZBcUW6meTPyq7Ubs+oj31X
m4Nd3MheRkr1mQ76RBGKvhW3KX9NofVD0oTZbDj7GCqVrzKKta6UH3TIAbZJuc3g
dJj57osYH/drC44/HmS3Dff2gUcfEKlTgM1qDSWWGP9bhKXCp/HBAtq/7b/x3npH
+buHpBsx4/aTbwGwYCtsVRJZ+gnnjuUqzdZDPUXsSfPKgO0TW0nKO7BscrSTtknf
r/3jzXL7S7ksBWhM01ssJ81F/ELwuycnYHaGdTU98xGDDpvmM28Iora6kiMY7Fd8
MHIDnLlsBKkPTNCltNGAdnRGIjNhr3gQGjaj1HprvJnKtBS+PjPq9wleww9U2wKc
s01vzXGj65ftwkeMjMHatIfTzon4E6h5K2xhow6RMnp5wFljFQAlML6F8bmescu6
iPGtbrZmFegQSsyHzQx75psmm2JsHPMRByxSmR1CWpNiQcPK18OnVFr/8EYaptGw
C0pbOEPckUuQOuK6jIERBiJ1X0AMubK5eoe0DqA7YZo90o8NRVG18mxkBbGQ7dpI
7naDV3HNO4QujqQGbrQaSbrw5oIPhbI+5Rle76CEuABR8ENaGQHNmy4TGEeO7TWN
Aoaitk2gYCgSEzn3z966Bvc0pL8zNsT+kWjYBedf+Jf8ylWi1vqUogJIlB8J9Xo+
5w6RA9b1xcYflg45hl7JGho4AGXgNXoVuUDPMZGNp1ELWDzCgJXBImwkq/keWm0+
46A7I+BPnSmuUM++TLA9sAommn61p/ryNC4s0AvkMHLOkQW1Qz114WOtMHPkDDYX
wAmTwW9mnh9ILvj/8CC6Y0z18gMV7R0StAhvYgvqjPBjchDwHemmSXUr1s47l6o8
mFXrmN37xuJT0C0pHapyyqXNipUg9Z4klDs4IlsEq/I5XbS3sl0r9nBJ8VVTjT9W
xcRn/nIdGAPf4Rba/FyUU54Wyt03ogviDQvOQYdtXqHqED6ihUjC5ViTNJESZR+f
C7OkhedV/L/ISmWvQTV0cUli56QzsxnJINh1gekfRA2vTkHfcjSQ356jwIjHCrp9
ACT4xuWZQtBFpPJDdwm0YEOYKp392FIY8i4zgBew3Ng7wBqi3krrQiJxUAFdgL7j
ryf188PcTWEEqXWyxhqerHIF37X8h4nGgzA12nri+fQ7JQJZbSCjDPOUgUEqh7Is
X1b1hzuVxhnAVEjzTjfNJZI97467T/pL9RSrvHFGgGzSj5aSapPrxQlWZM/QLzFd
F7Eiz7nFWIJvurTKMO8QZJD4MSe7DP0VZDKvYPaid2QcDVCAghsbj19KRFfZyjdn
uqhKqKfZKwstUXF1tDk2vW2LSJEpgmKWTs4OxZkOMbkfJp+EPopq+RbFJCMtBSrH
t8xVUz/TIetUVd3IJ0ijlCGmSPgGDwY20gPyzVWn1Hh2ii+LbmrTqRwVKBmUP839
DzLWjQnz2Rd8d1pfZ/GfiHKyg51pCRvBMncnB9L0LkQebvZApjboKyr+gUW4Cpll
02Rv6tt81v8GU/SYmhVMkXOyPSD4o+guUr7g5I/wYFQ+l1+4cE93eb6kpMW3WS1e
A5AwaMT7+E3XH0gbLbD1/Is45gPoYc9blX4oPwLxw5/+InkhumqUE5s0A+gbDcHY
wfmAmZqtEphDlDRjOdic+Vtj5IAseu0H0ewcHke/I4gSxY8+ie3TDFYz0Z1l3SnY
WqHF1vxFMEc+zvqxWHvvGyrlboU1KoA8IY1AZ6e4FdQNInfsoc2kEA/dqAiN1UA+
q4bcCIuEOU1C168HoHWrz9af+iXyVblNh7PghT/FKsi2K0Va+R0qKwJ/35KgH2Pn
lN0jdXRasFV0/Uk85CYJyhuJq24qD/XWhnOKOTTFOcIC7CtK0HJcU2++NxRXmPbG
g14k3+BB4gviNhUJy634xa9ZeijAFrRi98O02ipp7VGKqIeSKuKUTJMdN7bCYW5i
D/a6gzdw2tQCusczOyCoImswXjeonht53qT9dW512rZ3l6UCTpqMp9kA3XGoIbmn
gw0N+vmRX05mGqnKf0UeRTznOtt3sgk/cWk2RABIuuOOlGkE504ZyOx7WxxQxCjz
Mg8EMywu7cWJrnTXCprtPokYq6bcfmnQeWnxzliMJKFsS1uK7uMzIgGos3mLJM6r
eOF2es6cnFyyAuqt0Ho9uN+RGd2t3tdj/9FrkG9+xn810xGwUVRtTniPluXeRTmh
Ri9MKqF9LpFuZiJd7VAoQhzBhvHx+zId427Yb6zVKjqTthiwJ4PhMF01n3fueMt6
XxU0S9bNK1aBx8HusNg1ScuCHUPmjnh4aE0VZCAf+Zheb7AQcDuxmEZzk+8SYV9G
4/3erQuWULMDBaDXyJiHWxtVRyvH+MgTX57HQrBbfPr89zlN1Il6huc3iEdAIhyf
IYqZdU4Jpl8fSAK58vSOTQ3WtfOjHAhIso2zNbuLPLwDYBsSGoFGOBbkUlwfXWl+
VIQ4t62m5tho+hz6STWj6J5/JL2XIq5tBWObBNbGmXEF7uAl0YX6yauNXoVcF/sq
VBHts3DoO6eKb6z0911/jhTb8LtJVF8Qho6tPFA+2Ickh5xw8f8rYh1E1563d7qz
UMkYI4YHQt364MmCJa7+Da0KZEb8EMyXlXF7z0sOirMCAWR0g6yN4sPQ/cEVInvW
HpkWPbHDKygU/DxUl1Myk4YRZ2iV0QGPH1KT7f9x4tAzEqnDg1NV8S1FggfNQrSS
5BavkW1TXAl5KLB5uE9R0usFHwwXKrPeQOtpp49UEvyjN/UbWeK+iqVtmCnHSwY4
Pz6iMs592Beyql/ZCOGepvFclZiOkAllnv5kF9OqEwndkScULZ9w2TUF6eMS6hpw
wx9CCieW8GVTIB6Y7/Bp7ggjuPhy7m1JBjSenzQrceCsnwMgcFTUUux3/i3yR8Zf
3hJf/uR7wqaa7ttyxY54+HMp6xiu7W5oXgJz/2Hxl8DO3YwR5k2eNvvzon/BkCrw
pCffR82IL6lZqx7/Kq6maYnBSWMTbG7bREhKnUlyn/XHI9+yb4X1EXvo5tn8we4B
eQUIK3ipCzfWGKaHhgXaJdY3eHTBmVr+6tSTP0Wk1oeoxx+cOKvtb5hb+P5UjRcA
LC96OJbXEPqrsu7l8Rbr5GDU4PxKcWtLjl8hdgtz+AMzO5vziFRkoRJ2qhh6cHg/
1Biqc/LBea8d/thzcmH9PC3JCNhEN/xm/AWZkSPAob1WMcSstYTqs4oOf71bx62G
hTowA1fcCp9lfakyxATb/DyeMlgP0/AjOE2NUzup6fwuCnPYkYRPe32eTQr3uVKi
JT4krkz3QPi1CLpq2ttfzO5wU/NbiDOrr2e12Fod8f94Pg3qGL4zJ0j+mEh8v8/L
wpYegATkIsYBrHvDo66Wv0WfGrAX0jdK1OYgl9T0ZwvalWV0Jl/3u2ZnRqs9Nz32
XOUPT0TyOPy2fuFeUfykDtzFCZ1238ufM7ALRgZF4JktgltGRYIqCc4iVz0Eavum
lXSodLEI/HiG33c/ZLXGKR7FiSLMOBMey4uMBTvekq0PSmvgGFkBnL4kmhLdf/0V
bcKHShckbIGSZtgjzfz/MFQgAE3opoqZlFS4R5R4wyRbvgdvtFkYFyQiPlYTkykA
I27LtVTRK4QEJcFiX1zMVZJVAOZpIS4dQ52OtLBumPcMqW3ZEOoMHOiO93Ip9/SC
/fGjtI7UujNseVCWeMxJkL6fNdeuFKK0Ueqc38j36g+LOGf5boI0Xlo8Rre5/Le7
+gShntm/jc41jdOKJkTPdgpyY67qRt6JoTSOLBNh8sfcnBoSOfzVYVdFWJWjqBep
fyABuWAOEsJTJKG3JHzplWuOYrDiD9TJBQzpJRwK+ku6JOmQICTDXJKqIMOfcDKV
gccNnzjok1S7jmJKywOb68T+CIzQlNWW/jmCOhMNDJ07Pvbf6NcjQ0BpBqC6PBrF
ThQzsdc82OuPS72qcDxG0Nn0wuu+5Cm+YGQU3Ar3DEVDBUlCOG5jOGySNhvfiGLp
R1l5jCpsK3qqb5XPfHW2IOv/AswkIQCorVGpwVrVFghyJHVnGSUanLC9umPmsmVE
W68zMQFAurkenvhZI7XBbzOTex74A0vKLmESeiM67eJnNE4EMYGBcFwpvSD1S0ym
CypfQETOtBQx8UO2wpCOHELTkmgcHn6Kb/cGSGyULPcybAlLcrjdfa1FTjNRnEe8
mTHf6kcd1vdhkgGydDHzf0OgfQfUIKTBD2hPJ3ikT6BmrY+phBDpWfjb0NfmWVr2
cpU220yFHQS20/IoL2ks5d0MTKBlmgHuw3LFiKpiFAj9WpIE4SDj7g5pPII3n6mr
LHshfeWyzym/cdjyNJGUtrpXzPpS1MQbrjKUzRhqWnEVXyWeiDibEgZi5J1Qtmn/
lD1crDS5GEUhgwWJxkaUwHHQVfQHR09jckAMZ0lhMcTM25Hwi+Wrua5gHwOiXzFi
co/glJHcleWBtaLgPv7GOm0a6+TTDM8zGECqaIT6zk8KMAgfhgnmoSGhxIxSQD/k
NYDlHLzDsQ3s4yEHwEaIesPjOpTP7BIZulkIzoNq7ZsYj1GHEBDFXWcksB3csBIy
oh1ACA22J6bv/36aER4h9TxLg9HUdVC3MMdeZXs46CE6Zzj8Blhpp+JVR3j5VUZR
FJHdsCx2eYYxBE+mXBCEnb6+k6m6ybJZkVgyg7hzRl3r2sHu8t3avAvn5UNTcYT4
Pqzf2Q5nN1OmdTLXcBD0OoPtDKdjruAkypSD1DdT5Vx4Rf/BUsr36pfsDQCA/lyF
IFpKaWDBjj/TGYhFkDgrKnfRcpJIDntlrSVcJ8iyRxGCSugLDD7Gr8EmMnAOsIzs
eQjXUjUGBrvBitGq0hNFxefNqHHhHde56YZM21BxIHV6N85m/08aknPc+oNltP0v
Ngu/fyCfhYEaFZO/MGbJTRQeLCUp8OFYdzDZaaGHEWUYMY10BBBFlkpRa4bmIrq7
46pw5Hmw7Uomsr8Tl5Z06JDcDlC27yuIhDz0L1v6AO6MpF3KthTMxWIN/folpekg
+DjH7FRe/N9J8vKOqMZkL6a0noiBYgmJS+y1AcY25KbxkI/nI8UbOKw68DsO4xK+
UkTItcZ44dZJIfx87fWFCIxEQ5hvPcCX/MO4xRJWlE3SBlMXJI7qq64M7yoJLSzm
Bgbj1IQMfNPb3pXD68oV5T5MFeF1x7ZFaxfK2/pfgtMTvg8lDmCA2xVFFi+B9YqY
8TuVd9RkAd9H0pwS9qit77TqW7Fcln9s5sdGE7mjoldiGfWxfiz/YhD0UWWBoIGW
TA6T74C+rs85lcOyA3xPTPLBTlcF7Y7vj3rJ9gZAR0L6sTTf/98+xUDMxfje2t5j
oZCoSYRxWU7Bw3+GQya2nKU7Tj4IjiWxia5IxATNPgNSFWTcB+FKTzw2VelJ2Mmm
RvwqBx9/hCgQBaG3ykXNzKqSm5KY3Fler8s7ldIj2/eXdQrVtRK1vsmMPT+ZHtCv
BU+BKxjJx+wFwBYFSInZGpCQhux/TRmhEFoHk1EPTNz9ZU5gwGRHseBrcuZ+p0hl
MTE9g87rXhjKZr8s6yjKC5/7Yr/cWo4H8PICPJBzxCyBype8YnTUITN60ZIOFgN1
2JRAJilgZrksNlC+F8GfzrOhNkOCBZBAhxUA9OacycG3R6S3SP1twKJlbaIxeYqv
qy+h2IQ61xZCo6grsMawShDy3DKHBvOpLPt91xnxtG0LPjQttYlPnlCFZdY4pJXf
VQQZQ55ZqrYy+Bck6WwawwTP+dynTxfJGGTd0JW7Wg8UfY2AkzWhTo60FoFcsWN7
fLpkvhINsbOIFaKz/u2N4hk5Ab3kH7wdFoEU5aBwBPvL9XI6EKhSkbwiwbKT11Gi
YV/5AD9MyKwhBkeoWVcQHfMEBWxrAd+qxlShRfJGMRWFnov1T1kajzqhURy4BxIf
bCzWXwX39wG0G3aS3s4uRd6luClNOZ+nIL98ucx4hE0+bvHFvSIVA1DbDI5qREtn
4bwEQi1gftXB3hrDm/+f34bu2AWFRb0Ov3BJetlpeFnYWTUpeQRQ7qFzDk6wwL4u
LAYBMhuU4l7E/cht6hOkEQ0HigQDAy9jguUDlF7IT3spv+be3sT5HG39LEa7+6aH
SbtWIAil5L8wyENd7YoBsVdtLrKaEPRi6TcR2NwYpjqBrGIOOAsakEU400W93elx
gzQRbY/FwuBdoHc9ck0zAj3HitN/gAXTHXhGan8pQlz6oIIRYhS0zeeDZ4RXyNfO
EQTA8h3ia2s7/NWNDmX2hOv7OAyMey3GkgkwI2dYWEJwh8Yl8N64jl19MYn8G8c5
XXIQZrDknQk9YstVB2XQ6oQ+WxcaJrJ36Ed78KKE0AJLdvz9yOk6Uax5MHM0EDXS
3zZLAXKpugssWtn8f0SadmLV3IUULQNGDnY+G1/zkJ0n8S9r9veIovJTPaGUt+Ef
0DUwAQHP0ccAIS92lNpB4tFCS3YN9TBnFV1IJu6FoaoTHRso/3iWyDJEuUyQ9lQS
Wnky4H6EEolk+RecUQBwbJg9BqA8RUgExSJ0qDkh3ESFxcMkd4iagRPYVtiM/urL
PMUEmrWGwAXFCOUkvX1SF4ygLWEwPwGLPK0pfsf+BtdBVlG9weM4FYgQ6CiUshpW
DSvqAvHZppwILxt3qP9tSzumTQ8YWGZafs5LLCqNPMgm2HPwU0xDp+oU66iefyL+
UFLWuyL6GwEWykw287yOtVorim/bsgJUg0o4YZhHPrYohKGI09epz4lQxjE/XvAI
sTfGmG2/4doIsi/kKEZZPNJw0XFV+ls8jG0M+79j4hYil09b+PNauFDbMrDzlYpL
3bvmhVdDbeI9BchfRUVUd5iRIu4Mi3jzqViNlnTKp63SjmyBdhVwT+mSIfisws4d
QwltA+ONY/K42YeWTqYY5P8l/sxRmdVXUqILlxsmGpu1uJGgn+hkiOIuC7FhejeC
rM/qJ5978Kf5fMo4Ydet+s3mSLXYQy78k+nZQxW2R02puuUfR3IE7DBaLROfUN9V
Un63XkfAHL7gEVr47jhwWATmMDZ2qDOv6HMsF1FnXHpBXZJyLm0+YTc2MyyYJaG4
+lvzncBHL0sL/xZiLt39I7cDcxO2LKADsAuNPz6nBzdeBO28cN0Xf47v89OoDGeP
MnDfwnu7EOREHXnjEm58ebE8i/tn+QTAusxu2Pny0bQXLVZjWMqpxabNxU/cwa47
zvHAFDx9MEXoOnd+FGy48rHrSSza2vhVrYwHK3kP6hNbOQ4k710TADA5RXKYBCjr
AFyQy3lYcD4zbiPo2ilxBwbW9Y/BjBoka1j5M2oqF8W0iG8ScczqA59pBDhucWcj
AYIaflw9zwbGnrGi5eLBsOz/2wSYDyENUyu3a8I+ar8YXsHeFtyEEm3KPDYeID5A
RkpczBspvMVf9iXue5386l1sxtKTKj/PdSgdGNGSqw/BHzjFGnDebs7VFkpm2XAU
+RB5r2U54IepY/REbzqF1yt3wZueplkK67qghBaUmxprW8y7g9yirwgbSMZ2AL9Z
3oNgQEoFd2so5Hr66cIaLbthuPTVzn6Ydtg2MAzKpP370Ad0HtHKAvfnfNhk5JLb
CItJMBYudHiOqekYLIb78NFyS118Nucq6RqcdfExJ1bHuGe8sZnhmD7VsclRZBjw
1rle2xwYMvAiqOhM12VAGYTH7qGm2jQ3BGWfopGqUfORD2tX5VAPOubCBoIXIgEE
a+brZ8WYW2g38mi+84w93G/XbGjcwcc8CLRJLrNUQyolMXeCYsRCwBMoFdvpiP39
lfo+6AfQ4r4+zFaAtOiHqvPJ987nwWen9fpHCNa22z23RTgZELk2uXiaL0DzfIDc
4gUBXARE8YArDVITQWiwtLwrRzLdIsyGm+Wj4b5Ppec5jqeoFjZ59jAixvGTMo4s
XBXYOFVc95HgJv4TCfh4SV+7fOxXes/v/85Z8KXDdamXxufc4ToQhnmuP+buHg8r
y2PiavoR48BpXq3KPxfQ+btvyG+Xl5V6lkbFnnVSq529oEFCs3X7XwZg6D1I9tU+
lONo/wOMKWNsZPhTwX4tZtClhzgVAY1CP8nk1nOkDcMZ9Yq/5Vmok9yCipJ3tjQO
URzteyKZNpweTVU194FN1YnCDVjEOL2vzTtayjdaxxKY9Ii+qPeX8CP7xmCb6nOg
1j5DpFmDIE+o+EIYcVfqH54UkhQv4HEiwguk0t203Bm7E0txD81V0cqStsOW/o2P
devzEa35/PvPiNrjeGgkWkfkU1avwVb6EZdc4Z9V9rgJNiHFlzpGMjLtn8ZK0UHW
0e1CumbHB3jTewZkWJDZGrUCrflqxMq6KCJ5Ijz4mGbzBxNImTyaZVZ8dDXeKdIV
x4tWD+vSZA3PM8sdcxnFah4JMKbCCeiQg/ur6DLqwVqYvcs/SwWW6x9N29+X9eer
mJLU90olHNlXejyqj+nc6y3CGSJBQ9z55sqBknRkdLVB77D8x1SchSIXxMjdv0S8
CbPaipZpUDfTA7V/pkuBvlNUbKzlPUnDGz4oApocDZsSaH5ywdldyhau5cUy9wFD
ipSwochxG+xvsyHQj21L+An7mLOvfMNWBAFGPK+WY9YSm8dcJuuO2BaEfYqHW/st
9mWZMoP1WeuHSAVLcWxbaCKb4jARQSuCuaaG65WDczn1Mk/Pmh4XyOy1g45zk9vj
XzaNIJ8jtDMue1Qdi0vp1nuShCs4HKfLU/j8+4Qn6su0fkNQUSGTz86V5IJahqOb
CZ4+XesJ0pICSn8BUPqpYW67HlIOvHnC1LGkLBaHRe6dT13fHXr56t7/QcSSBXpy
rNQGd2zmz+hbs+aYKWS+RJYZgE98Twi96j9KIrUdRlG1wtdhN1f/vJsd/ksoqyjn
zxRwVhU4ENgIY1X2L1O4QyBS0JJXGixZr5aUY/T8T5hmRXz9ZE64SiYq4k6LNb9W
m9qybLoCXPEZefo8g5MepUAsv+PNSgAq1DPaWrOMdJMLmUg0C68W2ifEITfjB/mj
dmzkbEs7YqMVEgln4GWJZFCk3mIxNHC7aDHWPNiBQWhxz3OPlv2LEtR5CcjYZkz8
nJ6m6LsOBXuTcCscUMbA5lm4kTtsUaG2WxUJoAUghn1cNI29bWTQ4HYxvHxaARKd
LNyWvc2ooarcxhOgeAw8AYJt+oVsANv8JV3xDkkMqq7DN6p8UA0dYEluD528c+Is
biHzWi2woryXefDu4XGD41iEMyQDDFqRpr0OxfUbbvfdnTfMi9CfH8e040OiZpck
j+pIPBHp6fMbU8ZromJ5EzuPTUNCAJZbsL4vOj8gVXUF64o4uqwF0E/xP2VVAeia
zQ+iCPKoAwibgwzM22erRbR3Z3gHrVnLJchmETrGDU9wuKeirzR9tGLA4VvVNgdL
PKWEghMUILuo3IaXrl8GHTFKzAmusGAnG29cYJVpn7p2VMlpKDIKOrAzimg+dw6z
60EOxEaFqsvWfxo8xf/T+enBW1aQ0MugCxWDpp+HvcUEvevmzc+4nd8TM4ZvtGXT
4xu5Zx5xk+mfENeEdH91sGqp+BAZhDmI1zymwG0xrU6qJp/5ehea8PfQn29jVBwl
VhZgpSDjeDHVYqyyFu7HgAEF6HhveI5BNcWLZGt34cV88BeuAyyuN45+VzgTP1Ra
nSSO5p3kZ5z5/t+J8QqkhmRF7BDxySaltgA9h/pmFajovrSS8WBTEfbGPcUxt34y
PwT5yaEqB1ho/QG/DIBcr83bSfSMA9oT3mvQF8/gkNlh2cOGj0Sjxm5oLWj2HxH7
ikMQA350hKq2Ea9XtpDfMXxfi3p4HE6pud1vQ7Z1wRAW7s3HuNk9AYJ58JBXpKiM
OrOyolMjKVflGUHdc2dUePFIDFkN5MqpFIjhEMNFdEFUTpXpUQn8hKwQrDBjK+NC
GBAC//ztRCTTCe9LuuOikCf1IzGahQmp5/0AAVZWd2UpxeOrzU/a19QXp5/iheTu
v6vlKWXqSWO11xtXMUTNSGUqpkaCQ9l4FuG5LF3YmAgK5gMKqM64JRpGyksxaYt4
6l3op2VK+IlR9/yrn/R2P2RFCrgQrKo14db4lTlt+fcEIeeNlpAdK2bmTI2u3YSM
ZncXeAajXl4wY2J+roFcSSVsUH5DruvZjtd5nJ656MuP3oy29kqMD+7AgdCzAxp0
tEAWBUmJmHFhE99R/Hvyh9v5Pvwy2mDUojlhdJoTRu+posPQshcWKD8qBKCqMpQZ
UQ4KH+T2Ip255h60IV1HNYmb7aO7Bkf+kWIiRjY6lZHwJdwR6VjhpY4/OgXopbnP
BqeBfRv0Meum7klIKAIvRzQh9QXtbY5i2Fs6FmRJ05FFyWeHctrLoly755IFugI0
GYnEvvxDBIEoKbhn+sjhUrGmYamWdk4DLfDZKIj87Zg4O89xxzYr3Rsg9o3m0Zl6
GmUl9TIEqCGU6fCNmM2AMDt9UPBDIVpMihPM3qK4poeRO/lNd56Volr1PYk41VgL
j2DWTyJkh5AlbdFkL3HKdaeHoYO4ZrbHM4MFk2xGhCGTG58Q6Gt9jwYQx6wU+ZWr
YJc1Kf/sYAzuIxwqTyHqpBdeNMNbag5pK9peji4rvJ0Q2G8C0mzn4y0MfXmAvmnR
v4O+Fm3Zz9NDWjZ3FS/0qK9ex5J4nnQpPIqMXpmjivA80hcAUfDIbZuf5o1CogmS
Dc6zNX0Upu9srFGlkahh0/99qxfIk7CyqLuMH4DRfcVlzaijZ/WvidrsflsXHZys
xlBJ/z8bc6jWBiORkta9v7KtHczMl0B4owdn7+kse//y2hCSPtXVD2nVuIFeOfbV
wE7S9yNlcC4j8vBGvi0DP6oRhwyJOiaPAaxyJvZiAPJZRO3tj/KAkw/3jQ5YnEkd
ihqshsgNDNpBrNDtXrCMVATPASGfq4N4T0m/6g2NNMKR/XHe3tySlohHsCBLS+lE
oRBnIeeBdpxv4ESX1KeAUn9ruavMlt/lOcZN6X1S07xRRI0GWDf3mVWnaleIVp+d
g1D6ijluVCa8bCzV5oiUvglMXzGkxYPXSHe1/ksgqmQLAzNlRnFcWpuutvbt7WgK
utRe6/avDRXINylCO43ubjE17wmJ6DSlW8fRhbMNYj5CUmD5lBoEigBIPMHLntyi
ADPLFMMke6vtI0aHaRGsXBWOOEq3povRTuwMEdzTJScF8LlQCtPDlo2ZpV8JBouP
sV/0gXvDKkw013AHGfkBvDLLFOqdpgx8ezNUJPm2mtpvwcb0NiQVXLTtgyU0knt6
vdXzmTpARO+XXc2XI6ZPHOevnGyUM1VMcLDn7W1ztVk3AjMQZ88fCQtVQ/eQJXkc
G1LNDgL4Z5Jg98DcQdOHfzyj/gEXOhkb3LpS+5oPSlRSmLOMX6HAGt1jk4EC5t0L
RSnk2ij2VOo4n1tnVRffTU9LUzgAkiWFdqaAQVULFqwP7zYSb4jNbCkBI/sFQqCf
vV1+RfMh1FSDwo8T3bMtyv20+46t+5109fTa6VlACfNlzAQKbpTvTccpETa8Ronb
CM9kC5Mb1/S1ekmWh/xZSIE23TOvjmI1vNxQvA3L5/7TxmiZ7I1M5AUO47mauhgM
hvmbQmqQ8qlFrG5G6T69xFTpZrtzb9eNpCt0OqamiCv+zuP0LNkFRnBbntUkdsdB
q4FrT0w3FCYp/HQLFJtOkFOynez2rzUz04S1kNxNbJPJXrTHP4xZQx9hnjeB34TL
VIP+XoX3z4yx4uK0jsgRQ4+IfDRdxMHVT8lfZ7gItXs9E4+4GbKk9wGtZmN9iM+e
Cs17iKj+ri9cnpBt2jprwGYhBptCWzXlFxJvbr7XPTr6y08lqyD8XwE7TKhl7Qut
wM/0nvL35BitOIFosAHIxEHI65DOhPg4r3gE+NJ/unWim6yyelu3wTCn89wHRVab
tXLO3En0L/NBeiWJU0qdedxrbCGz/fZoAxzsVtBKQIdtpxxIoBbLDMfceXVNBQFZ
C5VWDJzHiFbJmwcTgrJmEhDoexgOo5g3bhStXf/mqgQnOEADAdP1fRLagNO9CZQP
BjqCMcY8uDwG2KJc8oDH4z0DelfNBLJFFhrTniphogo12fkvIeY6dn6bRMSaUk17
HZHJvhr0F63ERgU2AmeYHF7Ge+MjKD8kjLRDCrlmeESFwvGdAFNjt2+rJ1WjCHYT
DpuVCOdB4Gnm0Fz9b6lxansiStORo8B+SuJWBamPpyj8zSomeoxPCDsx5nv07daY
+KDzsHAeNlZS/QhhdM1dV0njMP1idtOS3jeAUiDdGaLRyrxXa/kKYgDVxPGBLHHH
rhm+z8JfFoJwKe1H3aoVfM8bID0/KixyfBqmQt99R752N7iYUE3y5sQ6BOI0LuTu
1UgoWNedkS+5O7M+M6Lo1O695DAmPXFS5gtNQRP5HAhN+L460pANPMDRPxFg4ZrY
q+hOqe2Rw0BWEPMyxnaxOIE4MUqF8dFbAjEuvMDAQWN5oNNUw1uhcm85PrIoq+P0
HMHeYODglzud1on+StRnLluDeSIwRUxCONgJsYruJ7qRcHXVlN3cLPYA9HSOt9ZE
oOpm5a3OqTRDs0OVbdWpqwnwuH2iktPmbHpuFcFK27/SorY0wS5W436bn0zkqGcs
XpQXzln1piaM8p7ZJYpRVitj741eKMIucutoHWkIq81EmWRANaY/aMyRkdPVHE3t
0dJZxM6crTslF24utE1sWBV1jJnWyAtSsaCdZnNEe/A9si9XCbjY2UTLEG+2/IaP
SGzLwe3aSUQv9S0X6BVMm1sPY2gwGkG1Dz6pNVX0sz1hW1ajJ9Ox/5ikcH/6WxF2
a4a9i6JIs/wrCoAzm8K3tkLfL8sfK0TFfzu3PkR9UK2KBEFPeP6rbHMMaAFNibcE
VKDkF0gxL2zccyAvWpuJAwM9llkbMlrAJIwngnwFeGDxsbrHDCYR5auMfa+2DYE2
4qWwvzghM5MENx4VeGf3PKULbKaiABH7o7S96QH+tfltvuAC32DcmvdBX+b6J9DB
2YEnJr6nkKJjatC69k0NDVulf+Q7S3OBKyPd1itZykVAqiJK7XYcADG1q0TgEqWZ
mMIh2wuM9rEInXno5dVx3t0Qfgq8FpbpSeMkQP5jwG+jo5OhocjAHcjeDlAAUwXI
Zccu6m3t9cGqWRNWKvaZLStPyj6FIgiY/lOjcil2qpXtm5dLTvD/hxWBFNFQuube
NfdgH0f/0swib3ptKvs+Dzxm4l3NXSgmX96zLCv4viJ6VfPaBvjbOWkA/f7+uySW
ni9OFS4F+8q17PDusyZcwr9ArSO3ilxa64RO6ZkckrgUJoxjm8+GpFLUxZuRNMSH
nHCfNvsFDztnC0ludIV4w75cQntLcnRDpY+7wIDY+6XyWKYZSrF6mCVJrFPUJ7IX
ci74OrBQ9NSfUtxntQ1jaV81IVenoAQGX6W45XO8UvTThlYX88LLsTyjGASVQtNC
IW224f63F+qS/wQMKbv6KCqKRkiRiuivI45Waj9xc/d5O+nJrxKjObxTzNlRs8nn
26RThHCkT2aCvWLfTTFTz8+d0dJ1nMCrYqkWwADQoPkH8b97CXtXd8UwaEZacOca
ab6a4fbgXzwgQ8SLa/aCQkQH8szktfOC2dj5x5JzqKPqJE8ctpb7znKEMqRYK1MP
d74ghZo0/tYYLITduq1cX/0Rsv2EvMtUNkZw5o00a3hZXbThy7BCXxpTict5KmbN
Wm8wrYFznw00Opy6ehi7g6/TrpNaAo656LpJey2GibExTApr6I7qKanas2aTwDiI
cq+QmlkvForaT5y5YPm+bUGhzoIw72W/vPpxG5nwB/HGPI4NP6Ehd8daYlKsCWCy
wifzNT/sSzDw5IGaRiAR88b40GrSLDi2VrcHnt+npgQQjrPx56wUWrtk7qEbHlbQ
tV36Ph3m+iiEtuwEkBBU3VyTaBXWdIl22Lzy5T+7h/4vvzFm09LX1kfI2jeoo8wo
aKqZ51LBbLoJbcgoyYMjFi0QQsbMzOa1rZ/0WZS8MK+lsVOy7PKw87gQF8VZggKr
du+ieSJU8R99zF4teapWM5NZEL5BY5xvJAEgt6+vLCUfAgwMu9UVfkl6WYQJaJqn
V9n/XOr/TuYWOOd/6HwpG4X0qlLJK8Tp3pe6ZegEQjSPSR6eDxWoEY5oqsO1i5ns
bh8R9OtlwCMI2bjkQic6N2bTGXEnBmUXc+B1zbA0FOMqFPo+sFkA/nJgw6E/OQaD
pyrELsoJUVoUmmD3+zKoSyE3cv8HDzGPZb05tvYfY2UA1fPTsIqpaqYwdNqO7ksr
dQLx4PtxnpetUsFLEuz23f3t3H/gF25F6ZCKCVLgyC6yJbeLnH2AdbGsyM4XlA3O
NN5FZOpSktD6cPNzzByEW7xg9ZW0BN7mt1P1hanZ7KmXBKI0Nt2xnHYNVt3KiqzT
a3uY4Czz0yGoGsdeDce8m3X0mkAb2jdFm9QHrxslKuisMEISe0XM45gz8IWUtHe6
aWU+iuySBnBfK+Eo0aGu9QQ7yQczHOZFJp+ZAbZHXwd1vl4g/ViE5vbla59sqDN+
UWdMrQujffgvM9rVEgtIysDcPSdmZopgb2600+GmG7JK1pj9l4ys2b2Aj1oblb3J
so0aoTaezfPOl3dbP4cNiz9qEMe9C5SIecMMpXU0DQTg+bc0KNd71mO8zTI5IvEv
lmJoQ1uJxkId8R9OdYg1ErTo6xkThjsfU35OW287wGVRehKrU2ujOtCjlSTtcrbn
dsZ+8bxPJJu0TBbZwFCnNEjm3tW4xvlxpEBBBs28GqBsEqhYP4RNzuNxkMp5oKax
g4+vWzMxynca716uGRPFVh2rbLWzrTQXxdG9DIdia3IDR5jnfqjVGCDYgs3ZMm9I
vJQq2/Dy2e5+r4DqNjvBfdqWz5NV8gkrYaQ7/O7aZ6Lhz7sQauqBZW0Fxh7C8eSW
BgEJ7NIbepMTUTvHLqiFn/0FDM0yOJ4d7SDLKsbo63DxdBSpfRTrYXwm2u3uxZCp
uz07pyRXR1vD6lmmEae0yVDHf0ZpAgt9pXFeQtmjLwEYRWl80NulQeF2Hm9sajAs
cUWic3isqUh+IOKXMhTpWEbO5ymuHn5GU02nSfY/BPP3YHZmXrayXGvEbIV+jY9P
/BsY2EcQjqiUyr6McciWxPCeFcO+0NDcGPDorbspq1kAwCXls7XkPG9iY4Ggdcb2
ZudxAWI14zBpswlmUkdLHmyRqrnLhEnm8EzmQoqMRhdxlVkt+SWXyJQdxobAQJgR
flxE5iXNsmYKurJc81p8YPx6wA3wI2ilLOfZMokCKG8PAwiryvQKv2y49g+SzFlW
0fYgGXY3GxwFAcaPz3ue9mJvri462hLATIoHbdLCRvbIzCyghGQEjnA9/osnv60M
h6Ae5AFdMtjnVl7updYwatZ9HJvqMgp8yo6dwRPxpdyBF6osYaF+Duau37c0VQI0
+yAx1V2QyZNgWF9kykdBa1vxWHAdf0Iw8wcCfYyOtmEpR7TpdLTOHuhF4ApVQHCV
igd2InNE+szoeyyTtGT8tPzjN4GWiyONrMNHZWzZLqNY0uZOIr18oQ9R1RCKshd3
p3Nu17DB7Epz/+rMds+gWIUmnXTDJogyh2SL49RsAZ8H46RR8+G238yjxy7nNmaw
W8A4s0NC7+Fm7eM9e0/EZL07o4RYsBElvsvNzQ1O5fAh5pr5Wh0aJaqoxwUnSvuW
6Qvi0Zp1yS+lA7BYXk8PFfRJ1wBKC+6UEYWupSlFaLcPonwWeq0EvrXpOQrWnZjm
Pev2xrMXxISxhdNPuZQoggScs4L5B/4SWoif+XsH69hQWL192LOSmskWp+rWf6Pj
tMmIhVP2fLjIGxnOsyKjXT1PK11KUW1PBnt1Yv/Ib2tyGLVmGBYGwZ2d6abdsOMg
yXkhrWFTyZMZHnQHAYyPRnelC65pyCzguOMAgSLZKzt2S0fTGIZtlX/xIP9aCtMK
jOdTM81F0QxdhbPRDWgFAExMlg+QgT72dA7cAi2ATdRG7+k49B2IaFC6GbaKrSB3
AJqOdmjsulgYlzz8YJ2KQr9OeRu3neGIQidNTNbFCLxJwq7MaYEx2L7WmYAS1ymk
J9a13vZBtnkUUwHYlQiNC6Lov0BaOafFiEe2yca7O88xg02of/6IUXJlpk6vkiL1
ek3MaoeCg7xO8g/FqOJ4YycVO4JqgT1NckoRV2oKQdyks+dpod9RFDkMcGJkGH46
QeIF01d44M+VzlF0pxMTm2pGubMoCyWsBm6pWHeR/wvrF30Vx7ppR1U8EUyBH6zT
XpJV6vIyJe2UVy/OxAepVPk2m0i3RLiWxmmQpxKUEunKxI49Zah3x0Edu+72DF2B
LmrRiyd3ZoPvNjhJ3UADvBxMF/Hjtuw7T5kCDIqDVPdp68UGrMy58H6JKXSjsoPx
fhu0sWSfrkBida4LIU7ZLjdTc6II8ODXObNBOD0h3bSK2mRDFx4lXZXhlmdEbOz2
QElEKgTp+aEriNzBzy1TgZ0JVHoTy8XKNkQFiuqzQKFC8TCov6bE3cQXVCsnc86T
eDQwoHMteV1jiz5xa0I9GxQpieVRGMr9+snnVIt9EReh6zVRyTzSTc0jmNziCtSv
RuIoTDoUwfPv4h/GxfQfbvGwG04BBbCnmdH3lrg010hdM3NS+e9ONUXuy8QznkUE
9U3A2VNv+uafOxtWofynIb7UU9ygKps1yYwZHffXGrxfGNJP55lXKRDQ/jCQ0W0+
EEhNO7IuGrkg3NGEzzokuhDXGJQ09+4dYvRS5qTsD9GF3cvOqXVO0BLdFeG7EXiA
DXxk9B2Z3yFeh7HiB8trJueL7C1mN4c7vnMeDtMllTS4JpKZm9nQmXow3WW2FRjg
7b/IiaVD3VBMVSqVm7bSROdU8WcvnuLCG0zVK9eDYAas2LT8oxA8xFkceWbdarRE
hIJcZQUnIl19izpgkxL8A15QGM3MeSkr3PAcp/SHaTF8v9hdPUv93GnFK4pf3g2y
OQD+v+4yqvoCABeaZtM3YmdIcBFiIBaC65C2tDd89jhIaLEVffHCLmXmPsChmZpg
vMh+kMVceiYffOXXnyYDnt/TaDUdwHxLcdwp0BKpD2YLQL8ayZzzIAs5tq6aqniB
j+BYtw1dEqBMtMb8Hg8unDnUNL4NsdxTHGlcSpmEEn5BuKjbiM0f/HVlJXB5jI/9
ZU/rwnvgKQXNHtSZNDYpHRYlcGiR6vFQHUbVjhlxFgFNeJh8EidtmQXoEt+wwFh+
lrRsMlO4jlUi+1Pd0QHZFWyf8Oxb0zSHZ8Qr3gLgB92PjQZUWbGkAcdfULi46iZq
CARqMnX1121ynOdXn442Kv2hvl2vdttaCrVL662tQwLQIcFWk8Yn0s3O+gOsFJlt
vEl9c0JAAQMbJrhgP5bw0dIAIdg6uba5atI1IeUxg0yYN+/9OwvSBgaAmayflo4f
LxhrE/BJHnhBBI28D1l48YelvGZIxNpnNg9K4rjyYUPIEUaQSCT/B6E8CVRXCfBu
UXy7jJv8Kq+WLUoo6fnPeqk0IRhwImiGZWUU0MSG3VgL43lhefgSNvG13pT8MW1v
u1DisUIDUHmF97iHY13W4Zuc+G4q+BBd8oIWY9PwCu+Pits2b1szu//NVo2xLiGk
wrqI44/UPsQoDfgYAA0rPrKeluLLsVG3p4HT6Df9/h7DoT01igcoloA6dyoR6E1U
vQ0/3uGuXtT7Ejl+ph+BXxkjiNOu0iNBDiAjcX6Jk6t/itIxo/xF+xilKOgIiwzB
+tZ0BBXWrB+yqGDPohaH3qgfW56ctRa2tAFnMWSbtaw8g37wRI3elswTEsSIv1yR
/gc/6oU80cTVOKUZcsdTrSVTdpAL58Qiuy6EvzedrUp/2CE5FkELzwMaepZlzsbr
eQtJlGdXeY9MXOn0MmI4J6fD/iDmQ9KrzohRvTuBykEAqqNYM4qa4RpQ8DnGHQE5
gFJ+yIUXxbviwegsHflVzS3Wl6l3OXLa6FMzZwhdvFAeNSxmMpIdpcAQoCoELhAp
adHCTbX/EoqrDKBOh9i/K4jtzE6W+zPppXlwE0a97uGniV5Za1SypjZH26xSUaf+
A2JsRvkNj+j21gbQ1R+dKQ5qHXrUOLRXmSqPlEoCwHNdMFdKMBcJ+DJKmnhnE8HB
FoIHQugXsf5DjaPF6QnrXQLXhLp/aOSdB3+p4pwTNnqpwZgC5GSUfU0GmJ3QyMmf
EM6X0SDwVce9m3AawPV0b5RpjVVSD91DPxSsRrOXlwpPL0BXoVqDWiZyRL8y153B
JEJ0yitLdatpfsH2dkLmnG9XrI2gTQI3K0v53d1wcoMySAC3aNJgF5HWhOxHtTF4
cqbSQX3UsZqAo1fYCoGuPt/5XGLfKvsyo226nas43cW8jaUpeaj1V3PP6Tq9n9lx
iv6ws13NPgcI17iQAGYAvOY7iSJY6vj2B6yCDDDkHbpdoxNg20IffURwQDS8G4mM
7MQ1NgewYwes/Ys8g5zOKGiHiGJVcQs2+WF16N6pv79+HDsysaHpwqztlLaxTlve
td33iLd+Sk/+hItO62fUybPwDrX9RRbIS3KFZIGHFj5Cw/OsipbGqO6mykc+Z52K
umVuJhAxJkKjYlcnne4D1EmHWIW/5tClxWVu0qfIfT2Sytte+64PiVfPTszOBjve
7O0fnspkDnevl9/tC5vmEeK0Y5ZBNcA8TzMi3pvdA3vxNQdLwuXYvJWPMSXfrJ+L
hlRvckgM5WscfnV26QLBQgorhwzMnO/yyUwwhHiouU63Q1dNAw1gxjp+ajjpteHQ
ynIij37Z1slmR4hkmdKBTUOTrS9vS5kFkA1vY5MbF/VFvM/Ds0i6yo2Hjrg+t1l2
aMhIbvQwyGx3NEjaM0pN+ZO0xoOxFcaCtlIhQuC7w5TlQqfBmUrJ0aYr5b3gZoEo
Rg9Af9ybM8Rf5vxswX7BH+NRxKrCNyPRKE+jwplUcp7FhVCBnqZ9KAG+8M3ND6mA
THwfDSkTSgdJDhcn/VWbPN1yEa9eJuxlOy1f9li4PiXGP2x7zFnzTX8uM+gpl1v1
II5K/Uyd3It0XAS1xEix7oqROVCWtCVEu6ERGvBsmZAW/jtEcYqKl8r2xBNUwNcL
NG+erNB/RQzO87UHdhEjaVO/oX1F7UcpVG0AXB4gBiPRtCNfNq1GM7bGtUBiqTSK
K7qs/iaUO0vXFGO3lgrY0KmIHcDot3SkNu7OS8eFDUkfae3WgDS+z5RGiCgRCuGv
eHlIE/O1OvcRdXpoUe3OYGUr3UZoDxqVRZjkhjykEtrWADCAdHiu+9izIWlMNguJ
GBobQJ4svK7zcOS8L3CN/LzjbfDYaCU3BMXRdN2bHKO8dV0a7WrXh3DCUoUMnaM1
fy5ASffkqradvCcx/BBVzxwG03E4cK79BYXeVRQ13hdtNjo2GPHJtFKhNKUMvxf6
uIxdk4lke1250z8CWpV+W3ySLmA0ec7FYjLvwWLh/7qhaQdCs26QvF+JUBUiqrLF
aOV1D/jjLuCqRJRBeA/fqZrS66+BH0hLU6ITsRuFYGDF9BLWE/NbH78UUl+5EcB1
FDD3epBgyZH8lWvuialDGBtYc7ZwyqEpDhzKzmcA8nRqFxiAR3KwSjNTAfB4wULo
ra5vX6gp9kM6H8l6bS5ZiwFf4MRf7ybJYbI7u8b/yUEEMQnEcWFB9IzXkKyfqbWP
25vR9YUUFHNydrDvURkebCM57DEiHTEqOkgjnMscEcKo3rkdovqDYh8oT/ZfUxJu
wp2bmq1P5GbmcW9irLsjnSMIWrq9C6XbNDXxN0APq4JjX+LEZ4z5sohf1X4cLEg4
J0OqJYbxoQQsaeSkvj4bs4z5U4BCyqdSO6eZ4uz7DXtZdzqaPWEYADWLnSfPGgwh
ftCtTGxe/gVCk7oIiQBRuEd/HxuRClJHDHrzElnos878t23rq1AVjGnzm2L/ThTX
gRvP/7MhCjRhLj+o8x+NxxzTnB5eZt39+W6eWv2pyF9NgVHZcAJ1+wHNGv9WMt7i
CKlimgyiYdPR+F7GxQJ4ylJjkX/rDoW43qfhiEYqoDMwA3egtM7A9TvJ6hF9KAAO
vEuxVduLNyunb7UK63pNU7tIAzA/4vMEmVKqX8NlDUHSFYA+pO2Ri1bb0hmy4Veu
BFeJPgj2yt+iTFK8XZ3ZLuAEPEo8BcXm6PvqRfRmECk50Zox+G/48Yhjq1Y2yRcm
H1V9VKaWF9Wc0LfcjhdTrWTkEYOXTLPQ+R5/HSoGv6DoK16meYc8iPA2ZFGM9C4P
2mSasNndkNJFJQxq8MsFA8Ewdd9M5Ke0QCYLjOCyotrJox39PH3VaE2KTt8uUKSG
ZnojqOhBXVkLy9dkc1K5BnDP6rIo+ezySheKrb+waBa2fNy1PLvocodtV88x9Wwt
xtWcN4EcFSc31p56ZunNqAuopy2dGYxtPrUHMNy3xb/qDTdXaHU8CdGJtLbIhGeV
aIkxx7WATazzv/05RZmyAygXLVKsEZi1TA+7ym9vT3VoJDbZryMqMMAcJGCgaWH1
dTmzXCyhtmZ+SaI1gwqjb5LGm/+dJFEXKN59i8/tTGe2xuwnUPuSQGtWRgWP+CaX
iLrc73ir8eOyaZV5UAU9wEbdfQv6XWvCevH+5FxJ1KDuIUieRG+Y0o6hgGC0MNGs
l6Lo4J3FADla14MG4m5io9zJvUld93fuoeKODboRpwYzKp0FIJTBQ+tJHBeruEvc
D1sMMKXfRfz+7BMffVidSvWVPzN48HAU1AdOUCAO0uHpOh8n6IjsC0CNRdSlXeI5
WvzGGEexWxJ1mzAh+P0YnRMP85esWivWVhIJLSWJGigMEGq8yxC2Lp1zMAsny247
5JLQlOXlmeAhCw6B22uZrQlmzICgID6h2mJetgdlC5h9yi6lESUfMgCMYZi616Ne
jplB/rHgE+QQ67H0KB+UnHWRzjW6fk8BtKSysuDvkIEe94aYj2+98R4IXbwHIybD
nPk3Zqh1fMc8eEw1Dv0X5YpzBwip7Pl6zStMYDDCQhgaw9jY8c3RJLlylhPuGKeB
6YXsbyHaqBT1KqzraPoH58ZpWZMQDr4yAqAo2nvREBU6MeRDokkYIGZhYwSXyYrm
8WC3qlJGtxj2sZSOuWDkqToYZY/bJdThGw61H+08vA1DImUF9+kYGl87PHAEcsB2
3Ez6aEZnX4UII2sa5wh355JpTAOJW/9VBnL59dxrJdqdwvYvZSLc83/dCEiJIgEt
MsTqEWtDYO/yK2CaWrsaVl92ytSTmsF87Fjex/R365pncKUfwxjSrjTTeIcpNewf
ZfNNJ4InT2e8NoKmb6pQy0c6GjPCKrRUMBTeAnzOfrFOGI0ibFzQwkUA2wf64fmq
8yXJ9heDM1W0dAj3bGQPEkkdiuc0xUJBKbYdGz0pm0MaYQsTuspd+m48ow170qYp
KO7WNafFIuEmtIY9avKp/2Nhvq1b6facYYsAk/yFPIo2TvPZI8Iok728ZJTobixb
pxFX9P4kH4ZHODawLm7Br2DTgllYfgV9cX7sqlMJom+evExhbALPE+RbthiO5f2y
nNcWLuwrSVihDE++iLoY7XRf1Btw5dxjPo9FZaF1q7Gc4/1nb8f28tVdHa3mOBmO
a89f6LvLKf8Dx4Y5ojAnM+yN+Eyeq2CMZpGvcJVY5B/t6WYAtCq8LwmZvo3vrcr4
aHKlM/TDNACdtFOCXFPpZVDlmp6z1Pc1twfoGBCDfVHs+txZoRQQ6PjPDYg4i1NN
S8Z07l7rbfYfpcNir8S/JmR08/hJuipyjlrlxOjgkXeFYPz7fMIOe5NME0eGJLXa
ax2h0QoY4uHr9yjkU3bW/1RNqCjOFTl8jOioYl2gIWSqUHrsUyT3bdFwtlJr5gkk
P3kfPIFuD9MP/KhqUfpojzjlPwyu8bXreMgfvXC0jddLFU/SrvPMlX/p3edQ0Rny
v776gsIObiSvGb8iPhz4bRySJTRN/0j3aMe0uKzqj0G11rEO/3j72RZWi92Mc4Cl
fDN7PxHetfUrzV2e8Mab794hQiW6yjXlCaJFERQ0ke4sLwXC5RhO3qom4ag68fXs
wEhOoYeLcK/YQj8egrKgbNg6Lt5p/sZIklR8IlP/PLTLA+ZKhHxwxIvEL7arvyBF
EtcYmIdXy7w0BV5n0wfYZYIt1vV97xqE0DLDb/uWLvwj1YHHXPcBGYNe+D5XtKWF
M8oL0yuuwys+sw8VjyOMOHjHhWrelQB5brWWF6F20k0ymE+d2gjxzmtu6vHQWoFu
0X4j5C1u876MhYGCAIqQrAW+NHP4c2KcBonznh2dn8ewIQaJREKkjXzJSK91GrfA
tPGcpV+sbHZTNzfQ8GefVV4IXz8B6ZVbMXlsDl7bMx2xQXgrU5K4SOuQmhdIhujt
tl+mQpWbwd2iKZzPUNrQ73E7ps990jHOr54KYVv8BjHVOtJi7gvCbWpWzYiBDjM8
H0kqVqG+8Ed5M/3tIsD/zjSHu/YbRm0S2hc3bXt2KhHcyRoqQp7ffCqSu8l/JTVQ
pQlXLBhGuBGrlF3FWuCSe7u3WGBLOziCUSOIVV7v1SauwFIdAFi4wwjXt2eBalwC
NWiwCaKHUyVOamL/uZHz4acccI+nJDceP8l79KNI0Mj8H+gv6NQJg1d37ZEfjEOe
oEiS1j5TsGlq9GYCAjfiYNfU7ySVqivFnhOemUBfyDlwPky/L1Sh226DGb5Vwbvs
3qmhiM8PVJbzvxf63atPXa9ORtwybOilbgH+bVZ1WciTGc47gm8YgMO+HnBofGr2
/dzMiuyPChg5H3Hvs6WXVlLVlWkzT6r/o5LHW6qGbYAcrG6aAy4wq5icD35NaDIH
vJu88RGh2uc870rVP7prqmN7yLVsf1L0bR0l98EQhDOzKpd40M4V7wOfmvQDqMjG
bRotjG4zVepahvyrdkCydz8tpRXPUjbgMNM+AhguV1133KApxoJGATEMLHewQd+y
u4QwghcKjdheK/VfOG+mCWj036pn8dX1xA3DDIwp7cwzoerxiSXK+GtrovIZRqTr
jgxiqjUPwF8IkOtOFU6ksQsZHRewlnnbOxLxMjDCjPQFjENSXYJHYa7mYeTDmPOL
heVwFZh7X1uPI339ysbQW8ZXTPGATqdxbrpbZEy8opO6uvnQB5hmfcBJzaFNaZ6c
N0RXaSrG+VEWfYb9GzDskm2Up+whjAsAswtLXMTZgE/+CKtaoPOeULKnbR3iSjpo
1Bk11YM6cnUyzXFThzc86C3PZDZB/3hfpHhUdMVuYlrVTSsqmCg+zIKpZAUrNNtf
JxwDl0duyzrP105mR3AZW8BT2gCJZahYkfIYZJOF2phCUOEwS5bV689rmyaNaRyu
y6YWDZp6zGN8U6jufWN12GjWgq8eIcU+KbO3nms7md4oVFBMZgd4FEklLAeUqCHO
O+BIyJLmv6v8F9ckr3Lf3rz6u6tyF9BNy6eudQsBh/3I8OsyaMzF9pEntO5UDhbo
FTT2VDr+L/XtKMHGI9rdzXprbewkR9E0867ShmZxTUFCwE5wnRuzkd7m28xp0rch
Gjgkmufby6jo+BOYghbDeZjMGUdOdAUabux5pomUspijb8VK808QBdtmV4tJF3U0
8cwpYz0fzOEz65+4Hb8RpcsmFpC3kxBB7RWd8Jv+Bzvn/wk+c2E+ERY7M5ajyNHG
78VkoT8VRnEt8vYNmysGBmPfqk8jUOB0s/kwVCrLJpq/n2GZpkdvyQRH+SD3KrV/
KtmcdyEerfJ2M2ORkivEG4gIyr50NpnUskxCFu7gSjXZjqOKbVIC963ftHNRf18+
PLAfnPO7IFw4F8qHlgP6PiDt2ODL0kF0574UohujVMGlxxi8Z3NQWSjzb4I7QyFF
AnyhvEGKjB+ZKNYglSx0B5Zqpliz0lk6lRHAklTukrCPt+Lma6eRLv6+WrA5bF5x
c3Lx4EgX6T3L+NlgPc1VENR7XM8R8VxoE1df25aCfgBeklgLX3T2hOPyz8KCmHCl
96KMxA6J3gmq/mJkbekNjvu4FDgetCkl2JShepwBPjwhiRzWxiEPUaSKcSX371fK
FjKYFMAVYFwJJoc8ojCfXD0b8XmoaTiLgtq8lmdfo/3uHP+h8hIJKAuvHgLcs2yK
Zxj6LisrRSOupFRUVmhukAp+FwQmTC5T4hDYuKf+3DY+il3PHR3EpbHo9YeDhE4a
Do8Pigo7qPScxSGA82RescPW1emE4HiWo7vbw0V/bdL+ZUraBaIOUbBJbZcTnYZz
wCC8DJ4uECIVwI81iMyaxBwNmAZHzig6sYNZW3HgQKKHW+Me65F+QJ9eUdU8W0F+
ogfey9T25kPCVp101jhiWecXPM8v8fP9CZKCZhmO7KddOh62a86kR8QhEAwvfSlh
6LjsJRXX9vaOBQz+SeAQUYI90lREtsTl0jY1qL6GyuA9wCcakEplO1bAglc17o01
QIOzi1740dt+Aj+5yMcgayBl+Rv7p2BIypVwv/6pQJSM1YNqh1iSi26+HUdPxkeN
Gps86PtL+uk8BJi9aKtnjwaUgSz3X2y+T4209Qc6/mXFF86P40R48lxedUO5UKQE
QBHcOjhdcIh3Jt9/lAoIuR8lizXgRpfEdfLcDmQ7QlA6fwQgbi/Zuye2iWAM94Mz
2wIUZpUPB21Cr53PPNy7id4zLhAdBKlvmQCyM2c/skR6ZyJyB52apnUmX/y/fIM7
pYwoSObp/rnr4z8AN8/5epSct/losI8upgOu+c3g5qCm3JuxVuM45SQ/SizB0w7p
rW2dtr0oyyX7fCpvLjAE/+dRQCYy8iF/Pf+AnXXDaWg/1qr+umjdpSNQZZiBHkqu
McSMsBXRqxhDNQN/ksfW9FjWHg5zU3JL4+rvj2ZYZjRhF6urXuqBn7rr0qIAYAxy
6HJ45u0Vlo19ar0qhk+gS6TtNv17YDtTzPFwMyiWLlJaEB8QnIJYWu7GSzwzHjaQ
u7bRE8wV8oCSgUTvr4jGzZ1bZlRUKxQ3nJATKmjePIRrlYxtHtrU2rCo1zS005b7
qA1gtfuud0vQZAy6IJhydzz/5nXI+6kkD9iAKGyfglLOFjFxtTooqxX1MrwePJdt
iUQTDG2DmtwzJigINNWlJwpoD9hi9yffLzhsF+DDBhXlWmK+GDuIbJFVuRJv4QGf
0auDHkt5b59Q61jvtjQnWzi/dglusTuBcOZZutzVjvdReu5LfBW4UJe4wSk2suwb
yZDbfpXsdqOnMgH1TlekWZF/e++aTxyliruz8URsToCVWJ08BkLokpeBjGhWKjfZ
Yw859dNGC4paD5Yu55vJ34IAAHkt0XL1qG7Rj571G5fMes4ZSegCqIW+17TyQnTF
9nV+/WcqmR/3WRDhl4u8DCJ1q5+AKr3zGilb/wRYMFkmqsD8GSc8gjwSGPRwncmL
+WrLRBNUnnYsK7RYKj8W+nXn6oGQiwzTHfMfEMD+pmVPLOi2t7EkDBDvg+LS6FCI
uRJZbw7DFOAj3W6Px+UFzdh6SxZyORSavWrMR2fISpMYsyEoc8FY/3pDXI0j7Seo
VkLcjXHQZYA6lI2ErS6dvshvlBJgqHoOJUz3dBgBIcZ2hWYek2Yvrpui0VIuTbBy
GeJX6Al6l7uDDU0uoVzfnDnv4ZysRbnK+BIorHkRIdfnupyGJTUqFXI9AX/BxQUi
O68za7UwSWeR40FePxdXnnmTvrj0tjh5NOJvzuSSTjgbP0nBekHSND1Zm+bbiv55
iDFqT120z+ND8ATH7y5QqMFdaiQvKSUorzrRv2xIDNGNnSFrGa/oaofeMeG729YQ
il2kFVyzd0sk6FSvjDdwpngyhIjj+Wh9zzqj677uNYrxDVdL9M5wl/UuyZ6TDysT
7weM8RYLKxT8dtin5XtxfC9/7w07RmGLTJpvRWWqh98TikWjxz1YMiERPUALhryM
vCxJPdef5dqu781xhPbYGvmTnrZA+Yln8zLcWdtT+GafErFE3qvTLSss1IMh+Pp5
n7AVjB9guywXVeKIQkADtE/8Kyt/CptjEhwXRDIL4y3yM9UYe0U+yL96wTz4IbOC
+36v+vgoJs3ZA0HE3IF1wMThAG8+M/dvjvjIeiDxTJsTPd56AQ768FcQBHt8AAcD
ymWAvKufo5S6Kg42Kq2vZkg8/DwaCkRvAwAzI9M6ymVlOQGCp/KybWcOEbRaSOnR
edTsqUet2XhoJLFFzYRkweDAxMDn8fZR2eSHLPX2+fzUNH7/MiHzhgfFhP0l4570
uyhRfiq3PfXpGAljlEhvkJHRQthdZBcN2mhwgcvMrbnObRjC9/AuXkFvKMggbK58
k6EoAPKHl4Xtg41TiJNfdwcyKj5RcLjltZH7qJsCRTD7EPiAjfAY6zOyTuWhqAfR
AuBfowCp2EnG9KqC+SheuTSzSZrOjtqEg1Wix8nn9TJ4krrxmtDb/poV7uRd+vZR
ppl7agblNmFwVDMj1R6XAopiuOSYAdDCSdEGsuoX5OhDls+34rjqwOnmVMigXbo4
8A1vmJZ/Wnb1hnaexAvMeXaY5gmWbb88y7s7VOayNzBRzXvJMCK8/ANuoWxo6YKn
wt4V9IUgGeNyR9FmE4CPQDtR3RaphO0xv3WX44vGp6VltlzETjOzowzn+5kezzZU
HFqyrqI7YPWjhlgvPXsRYLXVKu5D3VaJid0U8+IG7jt7thVvVgXhwDoR0KSEi4ax
ehocDztF4Cg0g/NArxpSNnYUG61i5UQ0UzFHaDes+91T1M/G2BxBTKCLTW8p/as7
PYNUrkK29cNZQ+wbyF9/oRLdFX57G2S7j7YFNe0Qsr/0niNCCgsO/4u/6KFRokM7
kxWa6gN85vKNRg4ridHLoFDfsewtOOc49ISdMWwOHBBtfDQrMu8OZvvkxv7L9J7g
sQk9B0nhBxpT2a/nU9+Yg1YiOKnSumh8icUHMmpbK8M7hJPed7o21nBCrE/2H4S2
SwzkoHm3UoQEobH89IcWew0c8RyaUf9iwP+pJrX9ikdQbWtdd5oQHbocSFVbXsbp
ozhBaXlOc7FGcRMVGX8Cx4BkpX2Tl+VdoOkQA5icMW/6WwFN8kQKNK/DPBMPGYRG
QHtJPr9ktC2P1DqVsebHVBh9wLCwgVYhuMayhvlrzxo173QqIQa3uOed4COdLcX+
sRsUKXOtrn7yy0GeKgl25vAd39wE5IjcsqQ6YD1aBF04aig+O1ceZEzrlBmUXbG5
CZtLqx7mEt16bmrlcWcdazRj/6E1nCHtxe3ez5ckPG1XsLN7eat5c9GmyiFSt6xh
l7Nlh4hXLdSf5czcxwF32OHvZ/bTSYd3G5Sog4ZA+Rujhf71eGkLyjoxK1eNBWe0
JK3ZUYf0bj21ZXdCZUs97/y/atF4F3Bbi/B6U6LTZ7wNfSbnm5Ru6Fw3CzXBl9pL
o2TogQzW6NyaSDqH5suzh7VsBRx8srjr/Q5LJr6Jjo2OMSFrk9CJ3TTvcpgH6ZAA
wVMezROo8UhMVEwkjd7oysh2ggpobpizRMrBPTK+Bx821aBK1YNf9iZ2YXVM5Kmi
FviaB0REjxzqyHi6juLJqjHgzqsxAvU0QbPNvoRT8IckIbH1NibwwgYRm4QJr7A+
BXcJWeNVewTr6iNyFJ2wgwDNdZoe5Dbd8NRFKudBECwyGhoy/lu78bfwqhB73+B+
zb7mvZBg9l2b4slwBfFpuZndV0ZkrQ2pkpKzie5JxroS9Sw2lkbyR9j0xMhFWVX4
qD2N59mr3j+lwoWW8R3X3nUiCJU/TcnVKH5LqFdxJzJpOazMdiMDD1m9Ja2/xG51
H/PytT/6+SeZSu28rBXDEHNKJkKbVv5JHV2/gkPiheB2y2dIg3f2XiCMaKMvS5a/
dwm8FNMEo49qUCfJlfiUgWQUbl47FqcG3zVgNWgDOpP8Kg6IC0y9201My+9Y8G7E
oKGfa7xZrIjhFi3xT/slnZ372Zp6N1AOXPnXOjbgMNMwCHQOK++V+GDleb1P5BrL
TDdye+YLtZfGmMvtHi1sJBTPWKh7fgIQ9LTaaCKuji2hI+VdMr6bhcGNbStPdKCc
RwyexZpUsHu395uyClH8ueHGdkTCACM0B4buN2yD9X/FUe0fPK7GdJPV4T+XT/aJ
ING8E0TkoxMZzOaaEGQ7ayNlP9RgflFNDeUx3bwAcUKkKGvyQgKzQGwoYwmEnOra
L1Wq9Z1nK6n4T5D5O40khcQk0UE/Q5SWzsvws5sDnA1lg641GJvYVLf7wU8yPeIe
5WQzgJoPVC/4gs+rBnkWdH5YpWq0WIDjjNJ25+XcTQPtmnHVbznYAH2P7zxUNSxy
ebWpyMtlkKEgk4y38wsBqe7dNKTAE14fFkFA82xkEif5T5nvAb1nPSJDGKH6s2AK
9Y2nUXY16hUJr9d05ZTqv8vEQDJO8whK5YvfOqu1sbvx9adItfFaWgRYbs8ooI1P
dODlszpvVQvfQWePr+jG/lJY4edcDVb6YkCxge0MqEFnl12o8I/6LQSeB37LCEeO
vtB2AM3oMJIUX0zVp3zvui+cNn010a0qY5WM8vC0Nb6NkQnAOi0v+1qiJRpRaOf7
RbsbkQrghExkFP5fhqiank0p/gep9dnO3yBgsid6PJpFnfpz2Psss4lMQSRFKnYt
6EssgKTNU5azppPAfK3qNMgf7HbrsW1tCC6hFfOnwl285+Gjbyd7hCm0atLF/Qte
ZRwDTmtXOlRlWGO57PT6/WBbaE3L2sMM9ci19ocxhd5U2Zc1UTyCob4rUgcVvlST
UC9wZFNACYlqZfWataSE/OeSkVEozr7mLMr8Q4j1eqOH7KZ+Y3XgM7NNG7dLc3tf
MmgaH9tnwxhEaAJLE076aKnCeO5qj60ChF5K6BG2BLa5/4KnbdURJpBeKqw8h9WM
5WX+fPTEIBKurt9TnD86BHP7l81e9b1harju8xRKk5DIoJf9UP1hEib68JjMSlcU
B8pJTgkWiAHGNOagbtjcCLTaVSqVK9HdJRX/N/u4N2Aht2hovezzbYVQ1iF/DHyl
K4QCYP6OT29+Xlb7P6X2ETIkfX1AIAyEN4axIbJh+/iSUeQzKklGnmJmjxzNpOcQ
UVAvAT0AAq3aA2ldVJJ2Fj5kkpVENlSchy/wncUu+6IOeUszahgkyf65VfZVOToI
MUbOUJKFStqOGfuaYEQzrWRtrMyTsY3G7NS6FoAliOazv1sbmBILRxssbq6BOflb
1WeTPaIy9u4Vx52uWp/+OdO89Gl020Rn8+DPZm+3ito2aEc83Y2fmj+s7yWRBBgD
vO+W9aae99AKY4U93ySH1Djif3qplt9JdOTRrsoBPtx+ZxBdhcNv6HH0xPwsdmFj
UbZdflKt66OTGL3cCo4frAW4zngBriMcOyqGjKkXBo+sHb1MjDYhrxBL1tJu0wiZ
5BFcBikWkluqCo2MROnXRcasigb0333LX4+K+tH5jlRN91FWkmkwQ2fQqUyXwZc4
KgiPJmXShgsiPOh9Sh9drIHY93fi0e8bM2zDEcCC/lWCMoscRgHqUVGSylGQisTl
HojGmdlgFkm7myRLeYJvCsb/+OXu6+pqvIavN9KKjfCS7lhX91PHCd7ia68z8dl9
o9NsEBz7fBIOxjbKXLoG+NYhfkGlDmQucc66ul63XlMIwWZcfuV1bTpTBgMwAYDw
LaC6GTvplalLSc9KW6OVRouPTRKx1yU11bZ2KdTBoQG9ew1unaQi23sIR9L/yhG9
wQ+PFNpp59ge08H7AioGdALG1O+rRBDuYGrAM5FU0Lg8WjfCP4zmYwXsO0bKPOnQ
1NbdFKnBaaN9IqFDS2OUxU7exoAimXS8Rnyz8/RDb9syCstoxynHCa6mXiGbY0An
0BO4CN+VpnD9aur++ejJJEx27Zhzhf2VuemieOjr4WW/s3M0SAiIPV9woyvNzkx7
pWs5ZQoz4KnL5auqijEstMO/LEyTReRwmgj180pFHBNV1gucNFIcGxM76jZyTrDE
Leb/JNgv9ljx9L17k6uHAR5eQyo9ILQYk21rKbaMmYTPOpWQyXV6vV8NACZNCnuB
A/d+KXXmPX4szsxoVWsVA+189++YsoNnqAHZwj2FNaIqRTnHCk7KsdaUXVV050LT
qaRhZ52qBdZAqGCyoTM0TzSdrsu+KssjPnjy9ojLshrWKZ4EdIYJc3UbcuHoC1s1
wy9X5r+9HCrDtQNMcC7XVSXmafBfNbK2ZrU6Z8cB/tx6YKNWq3LEm7vMQ/RVSx2E
WT9i/krdZWOreHzbUPY3Rcylyi+Ur5H5jTYyUZ1GGbuILV4FPecR/0My7Ub55ESl
Ln9aCpG+ZGGimehsuhfFecW1ND5gYsgSSfEiWEXhyho1Y1T3iqXiASyopA2yAScx
9WcxFvK+SB96pf/eczeFrldQRsH0ygRyjEH1MkPeaR5M/rfjZHILpjTEvxjacu4P
YWKGPhPWISXhC5U5XAyfu7QCpGBOzGqyKhX/U0m0hSmbN9aOgiJlkAo+nwoPuwzj
zqvMG+RAUiASWrAjng68k2HfaU6vJKnA3dS1CDMPGcEZjTZNw81XL9gk63VGxNWw
5r+OaIfEQPLFbMvn7Mi9lTvSxdBRxypPj1XAU5qVUrx63KIxBlmPXgu9R1TbolWb
WjizS44LEBGEZLvIIvPE7fwEkSp71DDubprW8qxRAtSJ9WJh5B6o1bHGOmj0YLvv
suzTAyBwrTr694AcO4bQUKq7KR5jvONUkJuaJwqznDUWJSUMHgFBWHerl5RSh1Kn
TsKYhVrsQ6fAw72kxhaDepY7nIMLmTsh1txGnGk31Jfaqoki9jaTqRGxqiqVTZzd
cEAbaRElMI5txHNKFEN3O0bj75FYPMG8Ok3patCm4+Bmzm5bsye4XvhCGbah76eR
RZjNJzNuq4LwWZIQjTUyllV2oVoZpVc1xY+k5uSqtppYjSV938wCUq0ssAYAdnwl
tnWIEsZ+n862NNVsU4u1E5+eHaFYLOVJembPtXhFYhSSOsy78L3lo9Iz7ViO7g46
pbxRIk3WJHDYU0fxVijMl+uc2mS09F9npxx7Ge6OiN3DxqHM9NYGAlqNQBV+1tLI
cIjTAn6780sWdqs/xJFR0WZ3lgqx1TAvl1Y03Z2GBbVSMKud59YUNhWr8VFYjD7A
/6Fv8z9vbmT6OFrukGh3zKGHtmXhhyb3aRlz6dLnUBR2AyjZyLS6jbLq08EHUBWd
7vDE8cJ1s15qrIDLHh5q9WNjHOV8ZmzGMoNP2aB2knQCaSwS/JVzQ/O8eQEGDu5Y
TCoX5XT2+TxLngfCoUcPscZrtGoy9lQY960bTS/Y69hKq6OLVlxgWpbVqJ5o4Yrr
tAs1yvAPMiiym54SRfA5kI/FDJZ1NkftX68EmMGqTlAcVRl0GCMdiupcuVsL56y9
/VH5wnTVZYSr7xB2pbAZC+03pVT8FJVxp/rwkAM+2U1v/YjSFRC60uiihoMkUFKv
nlp90b3NGgzaxs1bjfZO4CUxVm4e46xOD97vic56yQ5h4hIV5ToI5ePt+BVNWZgh
mlDZmN7HRwpdwrL/4RnB4ksUlG2FhhOvpt5dn8nfc5cSPcwMw1NVqfoISa+tnGgY
PD1LLQetkhVNtaWGZUY4XH8PSpqG0R16s0JF7APXFmxkiolNwqeEPTpMZ4vWx4Dp
9Lvq8gxJ0veReFkTFlo5pk7uRWxlozMgBD/HSxtsiGjSMd/YRd/psHlcYiON47eb
9zgtHZYV41WpHuIUGMYfcrtyvfxyT31WHn7L6shlCDGat4qj4t7ph0dPKtO6tbgI
X4tAuK8xkvuhbUHP2cPlj2oMncyxW2vrAW2GhD6jW5B2HFDqxpJlKD0Rm85PJ7oc
51squZeNXZDqHk89Z+n6elqhsjB8x7h8fu9PjKPTtRzvwDcvmvlTLe9mq5QLEqpv
1/xcnj9xPArgmE7ZNGnHlmogYFubuEPMv28VowD4jzdVlIZoAAao6h2mLiLwhoYL
nklKS95Velt2rI1UziuvjJDs4JztY0SeYIXiewNVPecjYjnNAllmaziIV2sbNFWF
hilpfCa8PLqt3axPQaVFXmQJxpLpgHtPWZOTaHxUGLN5QtwN0JyJLNNFarxTxRhM
Xax97uBQvs1zETCFGa/P4nlL1vYXy3/ZGZeLVvFdlYN7Zcyxbj5gjL2DGpAt1KnQ
lJUChEIHXap3OiGMJ6YYjwjgquTertbDE7LesMS0j1nlpmEGnUmCHqLw32MgW+KQ
8jyQI6krHNKPSOzAAozG1IBoZq+TDOKUxkJXLZdgoXGFXM0mMzo7yvBF8QW6YdF8
QfAeODD1p+pbMqHXo/AZBLG9U4wDKXJ5CihYstMPOrb7KWZwz+OwUiu1z054b1Hd
90mxLoqHWqfb6aXyyviKbBlloa29/7VP9W+EiUwXdQd6L2KqnP3hT+mjSANFrkIZ
zC/AJbTPrgIPDTRyrDuct4WMBGPNJ2XK29Jdo8utu+Jvdsj1Ux9534oA2+Mg818Y
YgjFf4shyi37OtpAWgZ3I9E7IYuMSZrYcCLgaPm9WFH35Tk2I3s1LYpNC7H/lfSW
+QKqdeuXlaiCin915BCUnfFPxO0HsO5rQLpZtwZo8DrNYMPFYn8UntbIdHFzvx4/
7aKhAYk7A8VOtzVX9LNIbUcfX6Nr6FNebLN2NcWQNYomuIE3DWSXs0+Q7Q62MiZT
Eg5U9cdalJ2uyXPlPVPVLtKUN8//CBK6XgFJYd4wQycvfP+3wiXubyZE2Jw+QotP
yY1hHl22MMN/zTEUUYLf2L8EiP0bNhKaf608i6AxOQ/xv7tIwQrY8COkfyPQHZdo
7Nc/KM3JyYxlyRzd5Lvt3AuNdWlMzQW3O6hQQT9oT1WIPspm24Dc+OY0BIyu2d9Z
Tcrc/NirsfAt9rmHZ/X1dI3VZqqXqonqkSWYbL6qm6RrZdbtC/uP/UaakA7cH3XR
LLLsqGPk1sgWOW38ogKwV952KTTgZsvl3JlzxKTBJXDyHUPSdby+qVAxW0kLOe5e
IkVllPZjWvO4Gfli3/GBe4NsITeRT7RJX0qeYSjJq+XA3MaULXckxdDNBrcHaOkR
NhhhzBA43uMf+aSSdahac3gK3Wu92luTo9XIfXPuC8KkTNdx8DRIMvQORcwGxVgm
BLG+8+Zr8bCWnSFrTNpv0lmgYUQEVyQ1Dn8bIZWQ+l7A56IxusKZ9SWkA0sTCLHS
9ipXFrRneQXQr4afn9kNWcHlbebaFxAYibrRHBAQ65+yMS4XvvGV/1liv+EKb09y
ed2nNtZX++cFmwz/joAdKn3rIdSSe2NhSrhRUWvcDTufybZnTox+fKtiwZA7+dJL
4lJiB5B00WcSwEtrNM/xlv2j1/mQoiLIifC56NTrPzJ008gQvUnZulI3AS7SGk3Q
e3lZSwQoqlsqPfxvl/S4uDBBF+NQCWU90C7f59J4QN/gQdCgIZqrVlmtyW9BpGKh
FPx59udvmWdelaGaNA6skFxLtxpKDn0m1+NJBrtzbwUNu4KVpF80JTeaHml6Pf+J
eydm+dJsk/8ikepWLowja8Q4E5G1Ut1oYoFb2kbKeYdWVHlsvgZpA/UMmQoEIt85
qKQxAH+OKlQ7zmXG+KHc6fH5uIoWWp+a+WtGTERBjRTBOG+YW8rqJNm6UeuFt2FK
8k+jYEE9yMdJPCcEfWwjWPWyeGXwPsTSSvY+HWxc6Rv13xAi8Qz7ObSEYR7gaZFN
FPOgrD4a1EGARMAWeqFkOAElWZJ9z+5Tg7+FpD2t1cT1xHXXcuKvcXey4aWjTI9W
wmSdK2PVm9prYAkX3HvGN0Y1p9piStRi4liJrYVFGlUwpXKjPEFtIA5lPgdxVQ/5
KTtb7N9yBDrlywWJy2K2/xM+1bl7M/nxIc/++beLB7wFe/6vOCY+IwIG7w9yn/61
gwPNFUOALgstueUd/g85INTsFTCpoRtNM2yHTkdM8/dOeWMyVyvOROgLXPgTFGcO
TEcFcU6dF1iTHKV6TTn/4XhSrMW2ijWImoyEvyodQFZqrVxApUfMoCOq7+4hypYf
h0x6kidx4UrX7rGcZLiICTNQ7eGV51Szump30AhL7GCFA7R6riKacp/qBqJzjiWU
brpIS/nd7hpjSVHYXz543CKejFORJ4qeLS2nyU8UfRzVK++LJ3HjEm1LvBjbjTok
wlsBPWwsUOB1y5xZ6xlh5lnU+DQIxlDB6w/NtuhQa3T9kcZQkEU6wQCG8+oT6gBS
LBqmchR7gXI/3dv58YJBCXxCawf6EoLUQVHvmvNS0t86oc/SoNb3MkY+xynKRLi/
2pTxmbbvdjblehPn9lh3V0kLrZERANkag+XdrAx2thR98mjmYMyBXLXwRWXgbCMl
fWu3RugA8F886SadLATGhBFYJTBvFlXRMZseLWXdVLgV3shg2bf6S9pdOwMbUITJ
5CS5V8Dtf3nmD2HW3WikywpYuLEdKulDnmeJe+rrvS5n/qKKm+C8blhFQH8Q0KHs
EXGx+vaTJW56+Myv/a44RuIf1jrQGbHVDUZNyAL8VObkKnw76eF14fu2ntjfvydi
FTU1eanS6UdPTuYg9VOtl/uPrkC0e2eOhzm2Mq8OmEgxSEtJ5yqKzguBKDUBQ8mH
rZhx5/Dn6ZlHN4e1DBCsbMd5VsCCUAR4c+XcEQuxR8R7l+5/CsMncOTw4wcPA6Uh
BUL/3yLPkKP8spbWtYN1QphhWZxz767CEd/okbRe+qJbj7RGLtmdtjdE0XHjNvP3
21X0ae/c3t5AQvC82dKEgMkbwuAgnQTHr0AldUgC72iquV2wZOTVftO17HaXosdl
Ly6Q5CIS0wua96iJZTSVNCsZiFQQgPcvrvvTmfzamGnHM0FzfW1aCPWJb8IMgaIT
XMVf3bC0QQgBPOqbdmQs/pqLFb+ysgXKCW+LCUNRvLlgS9iodTMUdyIk1eR1ykWx
YNSfHnPNdn3iuuj1aNEHfERb9t5+hqjbxnDjFmkRPr7lmyhCV2ql/2jz2QIqnO99
c8tyHkioiywxjuQT4pMf2gOKV3BU+09qqjn70OaLqEYtcVZXPwO1jutmt8M8nWwA
8+IOHSMXHHYLA89xLMQUlLPsl+VuBgBtPYoybgD2oQhPY6YrvB5O/XDkGBA5SO1f
JTAVykrAYh2xE+OJMvsPxiYi3SwFEfJLxl9tx1mXjj3lFXLOTWWDos+/mmJ5+bOi
O/QhylEMNldQHQXzle1M/rPMTZiayZf2MoZxEDHWwnuGTYBjs/OB990OvOQQzVR0
/+8LRKUVrDWldHBecIn6B6pXXznLx+24zr/FBUUxScnDOiqqCJKdOMYO0+0TXFfb
+sWW0ZIpJwuTvUiBmkwp5581OOStGgg6TbXkfcLugk+hL2uHqc2umAx3kbiJ45pT
5YnCymCegh6t3jGvUca6epPKWr/pOhb8ADSTIZpBt7RnAhN52wZJJmGGmfIINb/c
Jdz3YWXVCGkSb/YLxDZW8yy0CMI6qUN0R6ORsNDtJ2ER4qGp9vhmb0wZuBljRbzw
T1w58oTkyLXlxkgFjSVRFB3/3H4K6iqCjc7MCsU3iky7xH6c0RqR0JBWLlaJHssA
DH6x7Np+c7DfrzqHUEXlNjnX9M6XnYGWTYCkSX80rfB3wGBkKZcH1XLjeznprGX7
UKH0mxKIiRHkW0IBHmRuLFbKh6ASIrddDzFsPR0yxtuUJHi/8v0WtXr2sIgWtZl4
H92hQRbt9f9pMTBiFP1qxEx1URs1SZCurBt1J76D3744DqKy2cnOobEwlYCgQiGj
nvAz9zwGaUDJZud2v01xI7bHEArZWtB6qMk2pYEVOazXstPmHeh/i4NPLY1M5M2j
dRR9BBTXsEZXYuEdyQ/b6Yv5MswxuE+UGQR0RVVMqW0DS4/buDUekLhXzB/TOEU7
2FRAxUt4e52GD0u34mEqMFo6dRnZ4bCgA0iL2REbC9ax+DrdKXhB52ZQJjbSGDdL
7MCfhhY+wq2RRKD4TtRgK3jixJJubl1fuKzH8MCVZNR8JiQ0xwoIH59k2hGQuHF+
R2kKoXblWPh+wf4cHlyP1dLUhahflhznBrMvtchdFHX4myCJAeVLu23SqYCYXSww
KNJpY7G6ZznW056CTsUIsVMLeAfZreXRLZJdlofu40Udovpj0YHCEIlVLPmfbwhB
mDnylSWRcZediSS6nB//kVdfRu38Kga0ow7yNNq1jfGHhCmNYY3R43e/8bltjmLZ
aPxez8KwznNMIVG4QldZ3nNW+in3qgc8usJQKh5S/mS1NJOPuQVlSWAlBB3fRi26
chOAHI2x4G2+dFyXNV97o5V779twKPltXghy7uhnvvdKtzmLFkPnO7h46Q8oaHVV
27s6nATn0E0/SyfB9n2AtEqlHvP+IkQ1NtOAFTT9mjCJsgzErkkSKP+6NlAMC3H3
NXdG7j8DsBcTClqghGx6q4UC/+ke6BQn4rC4iJAX9YFNaV19mj63D/JBPboTTXMC
OMjDgOgugBQAOhSSOIoVlwgZIGSNviC2pvIvdJZM/aX+C1PwYzLjnHbIVQI+Mnh3
DTTy8lIgyFhIFR5uAuetSq9Z/vXK5e+ObfvQEGqnTdlWxeJMD8mL2wKN0NiWUwqK
MM8sdwcfkSVdULdsvPK5XCNSsvUIbN4p2rHvz6Oc503G5EkescqWAljq0UBxJvws
ZK3smv0uQBfdHmVUrFjViTkb/5a31GAgBwXjnFDV+rwt984kGxVb0OqbDAStFRPp
mUDTozHnFXGLQh1VVWyrZJ6iUiKR/gj6NeXGwoWD5F3GPfwi51e23girHsi6EUCE
OoDShBX48UWLqTncWXAHHHsb8Q4NF4jDIVupXUsaCPfgPXqO3oGEfR15aYv/nzmY
25NrCFbyqOREYCTFzt4DfAQmoX2IqmSSRLenIKjKXEc+Trkud0poVn7uukO/8wLc
IYJCIJhvTYLte0jOUB2rk7UmvRPo25KZ4K1RBfjtiqrflO22bnjEaN/PTUG4/KFF
t1ZDhAxqbS3i6bXFpWV3rgzDNcAFvhsiMs+tDahdkSUgElc8HJo5HbSZbKbpVcKB
JLaRWRNJ27rEozJaT0LdlVd/Y8VAI4lN1o/K6eEIyOhBkpcAI+pH56SKxyj3qjie
MS/bKwRlysHI7uO+6QH2mvGIzGkBQyXeE3LWTknmfQNAfAdRHZaAashUTMm3E9+c
ITmhO/Njd51ZUI3ok6ncEaGNdXAgKUkDcFnwYi9Cscns8srvS3ZJu3u4Dv53bryF
HfEeqPtLQcMV5KIi+gNzRFeKPRXVAq3J+7oVvWl3E/LT/gea/OF5oXAantXBUSAZ
usZpndSfp1K1RjPR4sb9FF0pGKL6Fscxw9PwdaF2sQndMBQmGqi8TUtiQpqiRHbT
WXUvo0BHq16W6jrPVTi7q2mX3bWq0p5ii6fYbClHCqDCpU6CW4rZ0eCQ/GltRrf5
YsNERkQq818F69hsqc0VupGfGx+sdJet5gAXgSzBqlSOxBtUTlyd8UJP67npxgXH
pWSvJciiKlsKR0DgjzLNegDbETwziAKDOv8IrQSiK6XJW3kb1vWT99/22LnK0Mwb
lVGbvc/o+Fismv8PNrmYyRYH+2e+EpCVOH9d46dDNqV8bp0oZLOniT2o9myrqliV
sFO8bnkCKixS2LQfgTBm5VDEpVO9GhMhOj27lJIfSgNDVyHPWSJjOO9PYn8oGpI2
7c6001IWJPwZYGyEpVZcoCG8HMGxJpJWwi2bK67QIJlirZp8+FgkP5UfHT+ICejn
SFp8evfB8ibzaCXSgLdlVQe5Dg/Or4nFpr++Ab38UeV/GqGyYSYjrZxQPmtEpSqw
qMNA/V+IEjIxxdAHCjqGWaTQFrYDy8B+okAR8kCHVpyncAZugYd3Fzp/bjOr7P+3
gsCMPaEw2AxURTDYRGMvK8GiUeywHQhBwLrw4hn7sUVqsnnxNddQDBGL0rYtf8Pl
sGrL/6MiVIg105DiJyjU8f82AIraRxAzdaVia1S9P9Yl7WnJFQdMjf73X3HU404G
rsAsqKDGQHUfTJVIdlbLJALecg7UDfU5xQPji2ZEsNZQYJUX4TSUGmH9v7MKhwtL
JKSI9pm8U+rroG6jGUbPlVaZJV8o/wN8Vbj+jS714PEcLh3OEWi0U94XbsTY0q8s
iicMq1EwaQOZVHTh4sgwQ+oLRj4sGMBoxyNGiwzaQH1mUtiHcXWBtqw7yz+0ioMv
zg8WyWtaBt26mpgv38ks3uezAhObt+bXfMmejXypZNt8iyGplXGwQhznUNsbfGDZ
eer77CnPvV50R4nILSvwHDK0iTYGd9bOWjdU6Wm8qkv1JsdmQ+zNZChBmyjTGQpm
z0qYqIGmlPIG1N6RXRf6CKqNB7hRlhW5U4ILYdKf/KsdPd5wGVXmuD4vx9wFYUM1
s56MlM940soOMeg/kmHlLcLnv6qpkUJ2c3wv4zQvh52Xfjg7QvRRurpV5nvUmWmH
5lkbMloav7W6736PLT7qSJDthc9JQv1HWWaw8DDp4XsQfeb75qyxWQTCReDzIFXz
fRYd+ALIxbtlOa5cJsGHCBUdRycYMFoo8QV87HW6dZPJV3ANnug2odmlogKOKYR5
zYlxZD6R/FK1pZwrlz86zx6dPevewDOAxsoblhAu87cSWladtFexRkmjmGr8cxYu
vn5JfbBZkXn3W8VYnKNw6uJHOztdXCSo1qA4jLnROUE51xxJI20I5RMz86uVUEBD
vZV/QGz2Y70lZS578X4BeCCApfN6uf+qLcGZ+tZvO/GFqXxyLt2AWCzFT1ncn9sc
HwQY0zYbFfPhPo7js8A2Q2cl4e6qTdjDpEyfKXlX4zhvsHxdtuxy6f76FfOYu8p0
/TA6Y3pBXA9c9clNvCnyrnXGKEorvNbnr3PtVNleVcCmrpigHqEL5xq+/TJ6+y16
qgjYBPuxYGKLzv89KSpGzTEqzidThebJfhwmDeEoggI9ly2/Lh64ZP3L9Q8zVYJg
oFbhjjh1UH2HRlgR4+j33E6nVlYLryU8DzjC1Oy7SdQo+brsL/tz2h2WUzuGp7n/
Bmq987Zd5Glfq5QLlekH817dOWtjHLssHQOcWaq5/GaCb3uT7r27WCpb5oac7kef
MEbqQVu9N1dt95MCe9V7h16X/glKb6MQjny3MMqeyog6S2Gen5i4zN+v7K/6uNkw
FQB37CQw08wOxtsz2R+8wI/jc/A/7HkRfusQSB0e/X3feEh2IPmdDPrkKFApS0L/
Cq/U+KV6Vnj2dyoWanFRAD8OsHxNK9A+WnVu5974cwaU7gWHjDlWqb1ZgbmSpQtB
Er5j2q56bVQYZ0az9+6PPth9Sen/7opzyCekk1BJl5coAQw/LjS5/99JQviDqe+4
w7tZ9+rlqif1DTu884fbaMVh2GT3P2xyteM0itEk/B5dYe85YnuD+2VpxTR21ZUC
RBaJJo/FkkznIDG+iPJVLda3Xs/UEKIyqk5Ja5Mkqfi1mLiiGUpNykx8fJXuQxyX
Thr7ig1Vc01dJrqQTt9UCTuHWqboQF8yfVPSnph6J7qZFcHTbi3N6bwZeNhxbhIX
jx0durzjSyPHTTc/sjhZVkJHkbgqFdWB8CPNR7wMQnLVVdMyWDLQO/3Vi1FmBuhd
5Y6ywH+VZeCAK8zLCGz8L38ter8ApvCGc1Q0ovAEXSehqPPzecZc7heW5B0kmw5i
YOOOpgBG9epgSrvoFEHn/B3bqDEro7XcwCqDWxgM/59jBDbZaNRysYMYtZSjUEJz
OKFVgKrGyqU7W2KyqkRuFeBA+f437p/AebVWQ8LMZb791esK+WZEciLmW+IYiU/Y
Q3EIl+wEAuOaRjwT1hedUzopgrkR8iUuQHLxoqqR0SmFT4Rd4Z6N0l+MNxSe004Q
VRAf/PLzEJcMowi1I/FkplRo43wVh48nQmyTNnQeGnAwzEBNsllxBPFaDdjlUtBa
mMSc23DQVpcsiSx+2VqCj/f7N7Yy/hDDmD60Ils58PHdN4/3G/Rwg/p2XxRPiV8q
vSGSvx9HTh6lTfjkYcRMhd4Tb1UJL8EBM5VvYMqclF7GwE0JYcSZsd0v820hboJw
fUkIQ8Ov4DFLTpYZHlEPuLwHA/CaxknE5pt0PHBNFubqyms83QOYlc0VqVBQjxim
pjlSaXch2UsXROPScaZ9YDecO/H0xoA3XYszk7Yiiv9cAp/YRfLQ05ByxTjflZtB
hipb6fTTOHMruhXm8wj7LKMCbD/cHFwR1CHhsgOfGVDJJ7/S1p5nwgcTpXAIuQ/o
4SHPnZD387t5HJE5ytme7wEjTNtmjCtmLDonE9ZCpby8YScH8INwq/yWiVjObIUM
6tUVSB5q6usTEIZdQW0yz28qWqCjXIiMv/7V5ZHpl89Jy1Ie/WjHKvIED0SntHD0
SBovkhcHQ+pZm3hC12iv54uPJA7DgxYGEuqNY31h7TuY9EVq8670qxs0+Wqhk9/F
mf0+OYLN5RQDjp9C3xcoIGVg9BC6SKLlXd9E7zsiK4kP196OvQdASMIat1IaBNix
R7EjHkD8TOnlG/fd0nI6HpVQuXjY7Y0XaRG2G2AjhJwDOMMq3DvrYnoKG0SmANih
t/s1MHfAAEs7UdEv13RJGVsVAo1dT7L4GA1Za9IwOSTnKanATlVcjudoVSMmGjAJ
Z/t4RvqisX57mcc5/62MdEeN47BEnYxQ27781rpFFiXBWtmlr44Zl9+jno7dxTUA
I1MiGDBI/XaF8g5ylTPv/rjoygn4fDAXIcb2boPuPo13uG2ngV+/JdP3c8SKA4iR
UVIN6KfZgXIlb7cy9/ovQ+nxoZskEtyQQgMeK+zOvQPS/De3ofdT2da49nNAo1OB
I58FSU0WGG6ID3bqYeypsxKZbQkHI3qiAhlWCAeucl+TOBqvdKDaxNY8PGE9NtaR
3mjhO9AyqWpKcPrd3zrYkuKU1Ni9gE2IZocQp+UgvWLMXrblrorWMXBblowGrGmL
W2yMUh/oHM23o45UHokKZJWKAc3UAo2+m3aUKQh1RtYaJ2J2PnYf0Ty15qpWxrGM
l5sCm6fj4osXgDNwEXGIJhPOnp3l5iNOdkUR2UiyvBsyCDMx0KerOPXjlUMHBP6w
nshWAmnsHvcD/LcRF9JO6qVLtVryknlmXlvTBe1ooqMGpPuCqFDNH83yg1328RMU
xE5NaJhQtUeiSARxCHlsNFx/BK8XOBogvw2bjyWOAhcSab3PVjRFoKmS+6/Eu3hu
Eahyd4gafDO96stn3tv8XHvML8zs2WyYdWXrkMe8gLqX9eu6q22efsLzo1M3pkKV
tCcEom1yF3XnFFZilKpLvZhiBJcQZkTpXu3QVf1Kv9hv0/upMp8p1jHWyeZovwXd
C9Y12iWG0f9/taLj4ZAem0jN2j0RcWo4g4yNTWpH2nnWKpNrzz+3/sKTFi87S8VM
zlClkghUPbhXau+iEmKzYWvWsVZq9EWmdTg9Y9D5AF0qFp1EGSfeIGVkYr9hle78
fY8LfU9rSlBGw2gC4VxkxLfws7uzbxXK8BQMAZ4LUFa1N2q6An0IP0mryujCMIs4
NT/PLm7afeBM5gHe+xP+NX5dwplgNVQW71uWk/mQJm8i04kjjAhH+LKG21+t06pT
4KnKGHVJlvsO5mXrjW7N9YEpsY6ZXfu7nOXX4ija01hjteSxwoEK3Sk5CTRyDUe4
xEYpEHme3agIWnUhg6LPmlfhd3aWdSKKnhXFEssDnFF0D79y10XjT9Zzgq4QH/Rv
fb+2k1hSWOnlRWtk9FTjBo83nSb3jhvmn12/G7TocQND6Sg8ztcWW1uNLK2dm98F
4NKbi6ZlOcfC59lKYUPITomqCBHziSnBt6GTmGmzDE7zPtA+dhf9CwT4294rM2lH
RcGmFHd0QDYX54CDSNYur5x+CBQQvfVpZF0oKS2NIV2UvaDwGUyx6pjZ+rA+6/kF
0N1uWAEQyX+6VNeVVSPMRn5MhOOLjJL+6YtGVwXIV4RcwtwLQ09Du6sZflLvIB3Q
uwWYfIDDsG5I1hy7uJckKNbrdy8ZpQlVrOMvhbChB0oQbtN+4h+lYTzM9psPTAwe
rQFKIZ1IwgjalgTEVPsZSbj/qORaJeDDwD1MnMgIUeBSxkSw35URC/GfXVJTrVDS
zBGuM0Ndglva01WtmiUvlXGsvtqbd6/ce5ZW9pu8ycsPI/UhOex71LI3mcFr1+R9
tufImg6JbmqGU162kW3LvftlWKgxlCEowhTe9TO45nx7WvkeMvWofLl+6ip8mU1U
iiNHXNXsNHAJOhEIHwKaP059sjc0/REGTf0viHr+/RU4GcsTHgGyMrjiWg5jHzTO
DlZ1DpsY0P5wZL/Syu2sHLwV6xFhiCS+SDBnOrO44GL3mmk0QDlo0mEv9CLNv7Hd
BAxW7M7YHuehIBbED2uf1abGP+NTtzzboOSzKoo5q+2Jl7HlOZi2ANmW/bMpmrhp
3Si/CnAoNElzJuV452eaDbzE1N+EH+BX0UnzYtdD4mnWqkD9plH25TCAAGb/xgW9
1rXXKOYgWp5xFm00BvqGGtSt87VhtIzLzJ0uJyoL0njuWAZofaZxCy13SS3L1YfO
VbU7nWwfImf1YBsFCFVuEMDcPL7oh2ZMkY5EEQWSQd1EH4jD6x1KEhOC43mC08QW
TU3fZqOsXS/U6a48xUhcCUPbjuyAW68CFAAfOG888tRWzmNZZfSBR1xxOkF+uVUx
VcVhNNLFtCvOyxPZLdJT+uzSQ4A6xQ4WdfO5fdQ4mygL8gUxF90upFbd/fAPooo1
QGpRG1xK0Bk9oVacKmcj2+oKCC3iS+z9NGC6bSBCKpZmnXom4Omn+VtHD1vm9Yoy
EJtMbFKoqyoHvNNgPjyFDlOHru0Y8EunnfIADmmT8WFHgM1fns0XJOviIM92Mu62
NsGqrnNiRxr5LpsIyV96sFJZYrT0MqMecvIObQK1pjSpGqZO5NWwaTaVA1E9jNI8
9qrfHYRD+dC8riiYIKHGWCcx2ntAnvmO894D+BZtJJOk/xpZlTyKgwlxPQjWfzyn
EIA+Wd+5+6Q3jGdszaleWaiHkZv29iqxHA/lQ8sei+8p5bcVcTtShqLtDEuZfTRW
BcNg+KhFeH8G4q1pYa4uMDc0ogATHZHrA2biH4IC5tR+byGAJ0hmdcY8urAFEpIF
ZLpOWeu/gyY9wLY29lJsO1s8BgGfYGgkbaAiM6gvTtKD1Z0wGThnyQQijHNHXk4B
xhDJ8OlbSkIZFP2GG0/HIjAVYYqi0Thuy0pjy1iNBWsdE/N8g0eQxzgGBJogciQo
IqYj8I86pIVeWHlKCfZrg0ioFJsnHwq1xAppBBND4YThdnaq3O7Bdo3c3bLN4/oV
MLpq9diXOmaj51VcPb0gD83jeJhnfCd/UUVvWX/2T3567IBA4Anj2rl4SMVAIA76
LSJsTSWjc+2qrAhlRi3rF6JKIjf4TIbn0jbgFIKbv41d3fqDzhhj5Cu0PLf1X5VG
L7h1nVWQLkxIdNIvm05mC8WBlJXv8jyEtZNf87yOmVIMuNVAryfpDPPevVBMpeRx
WXggTwjAD86s5vLN6ppl4kWX2zIMIICQ/8r63N0o5MhODxstXKbxUbQ67IFw+WxQ
sa/ngHdom72/8IqOUzM7L07wBpPZz89zHU7+xhUH+jZYvxj0Mop+tX9aiR0ViJ0/
BvuoCloOe3nKQdeGYOakMP9GyYgoVCn+b70IM4Tp+XF2CWq/6on4AGKWCf/nqyfK
11Lk3m5EbIxQdHEKwSQbMjvu9wh65UqCKsCs8fxqB9p4s/QbdX3H+Ev3JCrG/WFd
jPj9jGFCBH5mVMgYXTDXqWfZggDGry2kc+M4w1V2fNIbd7U/TvtMfsT4RB/givfi
kiq7T7/0BzAf2JDrkPMaOy1ucsj/8DIJV29Q7UhszAzGll4OVCMcUNlYzG50q2x+
c9FnyGxe/UW9cgJaY32f+z4RzFvU7PctUPZue05GbQewpEfz4k6vqXuk18HPLw/m
elaZqDwHEuOSixji7om7ANrZkU41FsZzuB0etVRUexdYDAAtYblsCIcMRKEV+vFa
XQcdJ+Fz+Yw3oPcBwTur2PrtW3qi6QYjnOS27ToOil2E6LcCrP7iWiOWFFI6rV6H
dVQd5n4W2bfO052D9rJguisad6egQS7gZWOLvOicvEHCvbH46C9vr26uw7dN1jzd
TTCyuAxLzlx21fDQR2OR1NARI5M7Fkak0lAQJQL3J7zHwL7WiRENHvP1PVG2ZcM8
5ORDxzx/W0x5ETrUzPAdGhWxLDCigt/70FL0CM9EHP9/wfiHi+4k2A6yV5mcnrGp
8W+5m3zetXKG2TiWZazE3YmgmecPVKnaAJ7Y4nmwIyfjBWWQsGLUYv/Ng1w+Rune
9Y0ycuyAYW7yuWbOawtIhWDFkKW585sD/VTjyv4kQISxrS00R6qw8jNLFT5c7ihR
YS0+SG3FHa/W8wXPAOE0KJSfkWAINbkJrfDfxnlnA3Ar/hstpH60hb/o9bU8E8k+
2vO4RdYWxIlAO+TjarzO6Ru0nb5E6/S4naYMmfJKZ/PYNcQQhIc3vXfAE80KDKNe
h0/hjhOuum/M1sYHU8qw83Y4NjPEbNH7ThX0KU/3dozDZkfuCLXqcT1uCQK+Jhij
qm6xRql4E62BGZBXCSlDfsQ+RnaTDK7Vb2G4B3KoYaU9DwF2tH9sH2PofwSCMDkR
VUuwp9RLBdc5zkAng33TjkW7Kzcsrkutebm4mHHjk0OWhRjqMX34YfUIv6l7Nwtg
TX7PoznzWJRfjFM/7406Tek/d07hcHTSV7UCKAxUXrWl2N1sk4Kes7wskH9wQlbd
I2zSYxYXriljJKvl9oNxd0VZD0xHh6siEMRJs5HESFDT95dc+zX3MNu72n043Zs9
huco3bwHpzBJ/Xdl3qqY1WVH6+KSVR3SwOuyCvXlubUckKU29p6eaTkSnJOHZSHs
EO5xbFG+DB6ZkJ0rfZrX86p1cO8elZzOYIxG95sBEXc3iHd6vs2f7Dlox2wwsXe2
QfsujD5pXjNZefehwZ2QIguqBSIYf5VzANBYNvQiNEF54WQQ19Sif2sxH1SmMZL2
rqv5CX1inmJ1F2zT8TtSSyeiPO9Ibsd7uHpITqM58xNO09mT4TI66HCo1epfLXX9
amnM++cztDNdn14Z/B0+bvGL5ciP/yQJyZrCgNntA0b3WD0zNCPkSGEmFomuTsez
u3Q4FnWmJ4lPqY3pREPLgumnYTsmd2W5uY0rvZEM5Jx6hLjeqF0W0KyiFRHnsYln
p5SVrJyV4TXjG7kVOscJx0ofqVkMBuSb/IWBInexo3agzTW3UliiykJmTzBVsCaR
8EvFc2elx2+Xs3qSlW4selqOKiEHuR7GGTEugNBY2Pgic9tV0bwUYnHKXzI6oGqF
0wkyiDAZr4P/ObxSdSAUiup+9cDdjaGwjhTxfJiVoCde1KJ2trPuo3Ozmw5hw2Q3
I3rwtvxsloRj6b9NcpoNNPI5Ju1JH7Fs6cX3LjPEEpv6R7Wcj2NNuzAhBmNPNjoo
cA/pBwdAznGaLQzVMJDvP2Kq78Y9VSwqBd2OCHsOsPrktQUUJ7pcF4XVbXKJWkoi
Vc5Oit3sW+ypKA+bSdRlcpWucd3cskbqQoGNablDILonVAFZMUGAfWZ39ZeTb21x
4fxT/p37oHpxN8mpAJ5iQstGHxLbQ7Lo4SWRV4RV4KlPk8nQG9SqlpRNWWRQ5gF9
I0jj9kKvmPNcUQq70BxEpWuuqUJRToxAHy6+cmhZWuZGWHFt/Jzbjrlcdc9HODNg
PDPxGQMQwNabWEclFhocNokhn9uQ+L24xdif0pZ+y5EyE94I2bleKktLtsWN6sLf
F+PikPFyRShPLqOczr6wkDUjiOFPfIT/CpZe+/sVIqe1XlZAgoOT1iduRVBUWgrq
TIpxj5/F236+g4/K1TT5ywMBJEDdxrhUhV0+oIhNL0Fx9F2rO0CkZfrrhU93jRNN
LnlMau3Ruk5ZuQryGEQXKGC8a7QvATWUebzhOx/BTDCgoJ1Hb6MYCbJmn0+yGqKp
059FI6luQiCu+gCbSaFbg1xouWkdRP0LfzY+mLbtvmRkrY5eRI6nXW4FBaswMePf
4oXtJOTqvtl2aj3gXIuvQK4r3dagJfV3Mp2plmKzuEz6Uu50vrbZnyJO8jeDDg0R
67rc8C5UwMklNw6Hs/xcVdKH+TrmyL3Bwk5p3WTiTL4B2lBY3NntQzjd4aw1EUBX
/PXSRoXC6bqgr8JF+6pCRRSw0/vNEu+upN2oO5yBaphvc7F9uWXh++Lrlq8OFoG1
hxsO9MagyT/u74UcPJovyzsjU9Vs7Jfzsg/eHup+z4BMe8vVfdMGk8FqLnErd7EE
4+4Pe5SjollriFIHeePsHZC23OHyX6KzCAr5jrKKtOwUptzF1gTiwXX4SZQ9f9ao
myXhVEI6GaQ7okBagNfMT+gge2I6JKt7enLVmEYbJJP1Bf8NmD6hO+WMVtTjZae7
g92CtRIDvAblnDrcNlmVqV3VX7oQpUhKlO+nXsWde0VfqHxeppIAAqzN9Va1AvUZ
51zYhJjc9/PDTdh6O0j8uajNz46/TT38tfRDFbqprudtAHt1KjZAA4BMh9OI+v8T
f/N8AbVNS4MsALAC8D6N9cJtdBGecjp3AVz2hQsmbLETmfkmLtsd1JPuHK8skptY
DNvAbofXhQy6z8wGNv0daqNMkCdbpzL3mILYzmWzYFu8PnR6+uz5ZWY5Y/WHhbO1
DNps+AbTihy1DxujK6hYgGpxm1wmqJWyvC9n82khOwR7xAa6S6uVuQR3jP49WxU7
18zeJ75ZFkHI2g9LPDrlcS9iTlTAeMAp0zRiOgceJ4Jr0RICeR5fQbDp4XONLLe1
W1/OImc2MJjpDGvaMBlub3eMkIpgDwTnxo5AVmatgUmlTtRXWVr0VMFmDFpbS5xR
h6cVKadWr1pGkngZbQgtavo7syh7dpQBgmXnQhYXiba1X/e6GIC5l7znRJMZQNgl
/zuJmCKWwOl6X2OQwSTWBz/HNc0T1+5cmk0m1kPQm+MLUfU0QbnX+DHKZzVlEx4n
gEdqcBymCb4irGVRdGxVU1vlN+u6D4nzTHqz0o+0LhYZc1rG+90KlvDI1b9WUGlK
wVovXhroWskNqwN9vtWoa7N9EZ9R51PXSxdzyGH6UjQnphPrToof0rLK+qndmc/g
F4zLglFMop3F5PmakjrSDx8WKVzhN8OZhUol8i5CvdbmJnPXZ6K4GWd2Mdgx/u8o
LQkFsDjWM/OZgCwfvSaacnatxvpzr884NP1zc2PixcVY7I5REmP4tTEiLbovN6si
A2vAgsU/umI6zSbMdII29n/lIt0Z4MUdbyRKKW49txv7govXBtTEge/e6IP0kb/J
g9FdnAgSv0sHpAJuxVB7XNXnhWoZl0gdw8KUvaO8geK/IhI8JLtRc6QhjqL2ZGZL
SMd1ucBRl6uqjVUCjwyZ3b2uEf8DWeIKVJrGZwcmuxVx5VcgIIk/DX/+jeEMNCPn
ejKWZTfAlnjWsO8juJqxXOioHZ9cMpXoRaEUvChc3YZKbbFJOIVbO+Y6rqEO0Nxj
rCoNBF+V9T8Kc1p/ggolYyRZgSGb0y8zIudwAXqdXIs2YdWz2gm5jNcJmrsVCRZj
SlV+frHIkk7Bnlb46Eec8y0qdKIbwZwwd0uie5wtWblqmis5aAt4xSl4vKz1wb8G
lyjNK12Ule0oca6R7V75707G/P1yvoKZx+Nh8cyg8u/CiG2gp9yHXwr7UJOoknsW
d71vn0crIpGvUgaYfRen+D6E4ZOpZ+UqVb3rUcPl/POdIJAPFKyey36ff9mZVH4Y
RDjSWiNjKYv/FlqJ132BfXh62paXMHHzJ09TLJ3XRxQih0jZx8Z2BBTEmVaGso5P
c8eYZIu1C9zEGt7o0auMHtkqA5gThPATNc3Ek3MwtpmaTIsrviEaUbxeiUx0NNAY
2I/6pgB4OBNFYWD1BwG4E6bmWrB2TTM1qrPMvIBhwdCsRBuPVJtIAvg0oXc2mXdS
Yr5xGRdErEYtmhA5quetMvKRgBDymhjgw3/LrEiOv7wm92LMwirZ2B+zEJiukjvM
gHPpQFKrsdHdVKdplMcC8GITVfG33wAPuz7qDENeJ7QX3rxFqrcn69N2f5imrjz5
JUP/Axauu/RcHRLPHVESDjt7ITH5Ixj9ek4UwpzCJHMVaere+zZI5uHHKy+NSnp0
0YgLU/BhfCpjvxvYHQZLufwUgucHV7mdpIUjNoaOvX88XFqt98HhG44p9sJZkMcz
yn/tVZvfsA72jLBYoRR56F/HMZNWJioNwWHlML9NI41fdn+c5bROtuvrXrB3Hhpm
fpqCS992G0VcZ9aXwixOSNrWZJYJcY5hCbyDia75T9jbWNJdeSKPFFrIBcYaNE2L
BAx5hRMINWdNlndS+C0opepTG0iqOPmRIw4f8WnvMgaXSwumCkM+WP+4iftpB3kG
8Z6+nLBOXIMLh/CKaZS7q7kgCHR/EyPqecY/FbRrJFzMFeu4Df7riohJz7EZC+CM
XGLTZneOkdfaZ5m5OJd2ER5JS78yMrT1HSMMEVCymfaf/OMTNqGatjW09OFPWjg7
5jf4f3j9JurxekwmGAEgSNEvKq0a7s9qCWe70rZb5/aa/z1PDJNNPhzXYkhY0RbH
T471OZK1gHS31LMCQ/sT4wXJaTC5CoMz0zGZP3yTS8n7J+6KTDmGhUDD3oO6dCGs
gUKpcGiCSOYxANYBLDz2gHdpO2G9Bwwa1qdNtS97BHlopxTlyq4AxnJViNgkHVAc
EuyqUdHxgw/xYWVIUe6roLyslEf0XjevO3PZ7c2iEEhGdU55EqNJwGsX0nQt0WCu
Iim6FFaI4Bsll2YAM86OqpSmqHngrr8AAaIxyNWXTqscZm6lH5MthteJIU6osD3W
ZhR3tHcmueo6jgh0bCn1zjklxMtgAfl1wEaq+U+Ny9nF+gJvhRnTeRRnCzDcrg7d
4LNGFk0qQrCq8lKEchSXpIaKofIY7vdyQWnsr8cmUlPntIY6LbsW/pivWNaHKwgo
eSTBwKDMQfQTczBWESYmrTQnacufOy0IZzsW+H9OicYBzEAK9p7g8BXstu4SlTig
/5WjBodzEgbGa1d4wtpDi0s0SlFkBO/YmhK4xo9Ro9eLGin52AAMdywyLTgGxGdg
DBOQVKmdAcv4vpIAJD2Op5fJj9qAvXqKr8fQ/3Ljs9tGvN1mWu8+YuSl0KyQRyIv
F/7AexKozGtpA88FCddtM1WgtEa6H4lYwPm2flmw9CCRtSIBVdrQImEoP5+mHdTL
qCzMXsnUtltAiQygsDnMrvvuy6OvGapbtww1YyS6Vs795GDTntpq0KACHGhJ7V3U
2GRD3LMPgdR8b2HR3AljNyF8OcSbO2ri0pzexe5Sdrl2K1E5IrcHzWGb96LX852Z
+/w65Fh+rFCsts8SS1H8eAbwoFDAi3J/ssKru+AZmmrx0YMPAqtgBmFWtnEXXES4
RwCL1Xv+WOSzWBtMI7SJu4S3cIxTG2JoMtwo4AA5efSiecNuVF82b1IGnxnSndRr
k40gsB83gPjYqr+N6EWnX7Kaw81xs8CCpvy4R1yMa+6HSpXYIS4b9PZgnHkLqnc2
9s26JiJvqyAAqq0gJipz+7nUO0FozUqlVgVXMqw7vzR1PXqD5iVYXzud0wg9HyaV
E7o84opMOr0WI/Q2L4iMgbkhYcKlhfBn0Wfp3jqu2kj+NFp0upwcO8bnhEl5hekL
z5V96SCKSCI8Oz7wTxyUcQcNBr9Plqwk5CAB4Vt1Khf5Xyzni7ebHgliUavPu706
0lc30xNnpV+KAcboEvQHqwca4u9QRdKRIITi5UhhjCagmq1ElC/+ZxOORs9hnmHr
5siZ2/Lg488Do6JzFYJuaiRaiY7wzdn1YQWKzSP/CPD16kjIx7/IjucQMEISRscA
RTm/FjwAW3q4s4QGH8eOWXJAmVLqXbaPhZOBD3xdizkp/VGW5HVp3hgLte7HaVz7
fZTEF3UQapoCq4nU0GTMjdgFgH6jGR7EuyWctoJQQNc/MOkKLz8miwVQSop7ss+G
oZ10NMo5H7YlZF+fqhkV3v9tZUmDTJ/f5jWEoDBxIrHMQOm2tHdKhd6wqg5ELR0z
/8Od+N7Yy4SIAdAqptR76VmtCIfIapWj6n81ngiR6VByg3ndrbDMUAicztTyMiNl
GGHBjkKSahp8G0J2SUM/J9Z0Zu21/HZkJthi5S3DrqWBfShprJv0sBzqOWx4tQEK
DnOh9j3kwXXbIbdP9RRoKNOZfmQtvO9v/t1O12t6qsJ4AEyu41PKNqj3JUb3+x6t
HJ7RLiNuGiBLGGz4B8orNcK/GVTstqlxKiu4zNtxZBmJA9HIq3XzPUd/mIrFwfyy
UaaDg8Su721M83z92EemsCWTfeGixg33OA7yvTwGnxIFFc9uuVdYibpglCqMpQNN
Mc1JzHkk07pu41KSr1k2HBTAiFBoiv37W8jU/Jb0A8GnaflImW1xzq0/F3YmR5Ue
IDP+JvtnK3+NWea97zf9UJ4MhAPv8jATjS+YABvjVUKGimFdkEicrq5XX1B9Hgzu
BFx//KDGtYrVfwMbTFgyvDW4u+wTERSyyr73X4E4L/gk2olJv9i1rxPYWRRhxeWa
mtq64CChb2qwShor+fchdYPqWeKZPgZuGT+i2Xa3Dt3pVHq48/Kk+34q62IC7jpn
AA3epJ82TRsHTc/UIxPOsIx5EJz4wdM8fL8rOKShIlz6tJLnMrk+lkOUnP9PUWTY
zNquxm7uUt1OkAfl0Yq4yCQ6SaPsKCWqdYrqSBaydjELVWZIR70aBP615K2YAGgk
AMHQfU99B33oTAvAAUulojIWXoS4dUzKCGJZJjOmtlMh9PyDwcn9UTiaP+ag36Jw
2lfIlDLFWLWuqFmPYvBKtN0/UugZOq99Qqmhlha78MZc/T+LCYjqShr6jP9o7WpQ
LC6jgs8WtltWLUgMwh5toiV4AlGjuGsmyotg4DObmK9wQeHx56KAS5+x5yIXIR5B
/wWyWyPq0z+YfYeeyKO7XRLpW+/RgqqSvJortX2pgeWV6XbRnDCvmfrUbRWJYA3I
CO2ZgOocMEB8VG7S+1/RrWwVICe54XGE87BJe5k+hTcDkqkqtBLV2bVehwx31Td0
Qhzpe13wtByJFV1AlJMxEVct/dcTMvrHWoxB42LwRB3pULAa1ToA8nogtDPXM31a
VzwpsvipJPlyNFPi79IExBeX+GlmDUdQjIDvEj1tqJdu220W1L25OWpfLLoccGvP
yTFwgZPHvuKGgcIzJWWMsFjPiUB2y61ZBDvr/1iI++75KEBTKTP7oD0CP2gr4W2C
EgS7yP3rT8XKYIHZlluBG2NjlVQwt/QWKsKhsMIDy1/Odl4n6f1xwyCMM+RZaBSK
n7juYnwu7xIq9LHJvUAgWNOviL461axjC5d9YD729Na/l8EpqZa77/k8EYQOLHtq
2vHL0l0RPs1udVaCAFNG8PE+PlaPswMjcAkoMOqttqD34A3SLDAblhih8hw9ITBx
Ger7VwGJTkgVRrq0TVR36th4/Zy6zub/agc/y6gIqGts0htjgtr9Zbu1+DFgxeMB
NcozhqIq9OF8jucdz4LDwFBjCi3H3GbtiMmPjtHP+ay4BbNeqP0+g9bMqSYwrqO8
zZvozxTQEiZSz5tSSKG8K9b8WGEuRsjzrXJIxUSeN+/XDCQLBv+3QpmiULFXourC
aozsYrB8V2DdTgVoJheqr2vGwQEYgkCDHu4qtgXpxCHpBZX1bE22SL7w64DlnVE3
RZL+yV8nFLSMC/0IvS4GO6XW2OX9t2ok7vgDeo0iiNs+DV5Q+zJEdX8Mish6oqjI
/SCfc8vAAgfqYmAUT9Rmm9thrEzcrdELtLyQ8Xm7JsXFrAqQ593VBXJigmDr99jd
GIWQlCm8qQgNHbFeA7xBU0+y2iIrGiNkLT3lv82cVpuuX3JyU71EpKOvKmtI0+aI
q8VFmrv3lEwh/qcfFpC6nMpfksMkRJ2PlQ9IijWBzq1fh8OcINeX50AOqTZRmW/M
3YJkDS/QEr777g30Oh6Jm9rYZdUHtO2baOGW4p7dsHjSDY2VgDIHzNljzrDsn1sc
CLUfa4orc7tmsIDqjNg5r2Fzq91JdU/obvboG8E0RPJGiZCXjbespX7sPGG9jYtY
n1Z9VPhnF66Kx0VREdcw5mYoyM9IeDCNBKpEBePdJ1AtsA95pQC0FfblledNHrem
SChOIExZ+rDl8AKnB1OngAFtRQZpsPsr9TTWnKERlpbnVTv2QYS2rLFB0nwy4979
wGmNW+KwLzw4WOsGoMgbX8Fa0u19ilxcgCyW1V9SyOeME6cJw7Kku8h5Dl8obXiN
t+gn+l80JUUyBeTTlvUpMSLm5VIKVUIBAH5FDA1m/R6i5oGqGpTyF/9tgAMPwbfE
AQxqvBrYyNDVY5Sm+/J724ybohjFSSYP/tpG6DTsWP1X1kefuxVvhjWqGnlU+f0o
BLOKO+jJGlE4wi/D5+U8p19LL3e1gLujcrt6jYZzxsKBhSjmQJmZeU65/BFtbA7q
BkAI2cv9jj1XN6Y3WIeqpYhLjwLeBu9V/FgPE5pJEesa8Vqv6yDUtTFrzKjVNbKw
PuwjAuzmy1GMrxsDaIQGQayxelAZjoq9YZVzg9PxZjGDFlB/jPZbhSPkI8O3fZdO
ba5C3RJITzdyRGHisxM+lYtalk3PZBArlGIL72T8OXI4nQQQjRz441OtVLisI5rB
7Nq6ZigREQPmw2YazGt0u6nPQD2R8i6IRxsMiGAr8oLtCceeL4olnifCKc1R86Qw
FAFpybgwwnQWQJHVJhH2eW2hmkxzdnp1CHugVE0YqHLKvyEtvHPZRFdX1NZZUgwk
e8cpNfy752pF1zIBTiJ4WeHCUxUbU10OK8bUIpjNIkN8Oog0yvYoxB7IPF8ZUiOq
JFILyDnfWKHK0stAExyMqyzRQo88fpdilFzU/Gz41WSRcQVS9SkSobr8I4fJSo5Q
IbSTGqdLHpNxJABAf+Bgl1aviH7EpttZxqv9Y0SwoiGGdwbN/xTmy1W0RO7ZqhdA
dcvMTUtYxoIFzEN0NfkYi8sZ3LZpGB9drBjAufR29MW+tbwxOJS8elPVFIluBrhh
hQ2ziKilWkF3TdoJ2/WUGNCL7BZX+q3XP0nlcNxybuUBdeRf9s0Eh2t4OHe8y/w3
SAGPNRUgmG1oH7MpONUhXbcpsPNHptn+3QmFQh/DBvsFZSv+9hhxdWDWKrbH7zSe
BMZL5tQ5KQaPg4YlLHWgBSVJeITwqs9iQ9XdAIp3AsI8IlkFT4G+vIgJ98tkmcmX
j6adnbSPBPd3Vy4Ted5/425bTL92aOj7I5izbKSsgpNDlbeF66hZw/qkamGr7O/O
RayoB9LwobLxTYJKYJRbpWydspm8w3aeqvEo0Z1/kdtYqZ848B8RcXsXJAif8/tD
2hliy79hIA07Zef9SMb4ydpfr0D8L9xkWyQevB57kMy0Vw9JoqkIDREPS/n/1DL9
63XkF593Dq+yPJprGGr6Kef6Qnjz2RxBk3jRueFlae9BaZ/UzaGhRb6ezxs0eNnq
a0OVfBiEO+NJZj+POl3U/cuNrAOld+9Wr7+DmtUfSGQ/TQ+3QbIM44GQTiMBV/9z
Nb21CP3qVShVT4iBpNyv42CCWwp170+fKi1HEVuZnxvmz/0ngvAytMtMoHdQHO9W
itfwcAWGMGdWZkRVE1teFi5YmdnV5DoJAx2nN0kPT9AFI9r/dVPZ3dhhcvTQlprf
m9hmG5EJl1EdqEELCrXxsRO5HZ48V5gDtYMwxyVxm8RXplHszFuKDFMMS6O6mP5P
vRuxHdEvljoCxzwJIaLKPvUbPKIB8XM1tM94xfDnFKJ+OaS0n3KUB3XDbDdp8Qzt
ygLqnzF+cIp3Zp+BrKVZIXQtozrG23H+VDrGl+RrLMs4jUAglwk7F4rnh3XjVI35
1zv4fWWrLlIkrI74pMNOp/iLOC9BUuJU3HgK+OWgcRsyB0yZYi+lMVXcP7lsTX0L
yeXvwYHGtWIDN3gE1nTaKbxywhIlHxzFBDlCgW/o3sc+doYTFiYWjIfyowtPGWbe
Jh3Yh1tq78T/fxcSxMxb6UA6lrqqdbAIolQbzGTTbqRfUZjUjpMfpoQWYbEAi0cr
eJrCzSgxHULL3qsVok2vD56AV4Up04MgJRUcogifuf3myayr2CvGimISJ0+r4dn/
nZiB788LNkugsOAKVlTT3F2YyujGhz/pjqWEHKLd5QsatwekWUTiL7yaVqCMs2us
jqF1DPCwrCWs486NRXSgacVHw2xpsactNo+9SchbkgwSEmsykNXWezk1RxoP/sJI
vbNzRXQ2436vNchJgVbPack8S896A41qy2Z+G7IMYG5Lfk9YmIYUBx2R2oEOjSjz
8cMXNW1uSN61kY+CG71hiepN1rkPcG47Lmfi9BNN63LQjeyNusCFzu5GG5WIpqdt
eoS6m9ftlyYhN0oFV6yVj21PvIQDjgtT/EzhWgLSnev60yTQv7MpkDvTuiBKoDLr
vC/xCk5UNJoaxwz7hClJqcsrKtQTS2JdFaj1adgdugijE0mzgZLzZCWgsLHLXoMu
Tp3snCKaItgasDkNIoZtvtHOqvRKK4kAEaI5eW0JSTCH4lRg/EtX5/D8u/kmS7EJ
jbb3qV4ctlqZLBVf3o4YA1tFqdnADV0P4mYYC9fzkLkL6Ji5YHVZFd81LhDuafme
FizZcL4CMEHnN/DTk1UVjLGUB3J5TZ503wZsjGbXiUQE0p7BPW2kIDkQ8/5RrUdn
XOnTbhzNYX1GWkzDf86txSAKJAi7ax8EFA3GDYRgKtyGDQU2duDLJH5hWI0589o3
mJQmk4B+GMsoEWqvYdWNBtdf8YkgegtMLOERbQdna5RPZjk1qE5k9JaZH/6qrmHJ
QhT4CISczePRB1rrPYrO8tgNY3YaomNlbxvAyV+VXKDE2Zr+43REtXQJN3sLmAVu
nDJRbaioOGpBVGh4PXuIevE8CJIrVPc97P4aKNb08gW6678a6BNHVsJDljyWOcaW
gAYBObY2VGHB/YqnPtlvuOXKxbDGQcUKMr4aszwJTxvYOW2WzaPAN4gIC6CgwCeY
y18iFpALhcS9gwR74huXYxD5YdSgAlmkvQPE1FlPnjWQKpqa0vlEz87WYDW9Flj5
M7gbO0+uaVdThnh5oN29ywDstQQdnpIZyuTi0fQBM3a33j5ewGIzVYQeH6cHymj3
8QJY0glAr1XMzcLwrYESVfAiXFK700PDWDCyTX5fEg/gbaZcqq5w2WzJlJnIWSSt
k8pfhRw9ykKtnPRW3ycfL8apCkvpEbDN9sJ+OtSCxE09dH6KusXRwujh1tNXmt9V
1uRjWr9fAhKWLHJZNhtfteyG2KsTqEZapuw1v/U9YLlaZQ9qSTIgTfaOiTEfBFrg
VaaiWEeYsx6hRMccMRydeV8QK+73Ii4CSlC6aF3R4WsQBoCULF12KGgg+/wxQqJ5
Vb0vw9pLizw5MwyLpOc8FP0LjU9Tf+/CkdCUrb93HrLO+4t48Fqi8W4CMxhtqLEq
79JJb4l+mDpCtmrVRZ4TQAdv7OACvgRd2C2zJMgA/Cel8Qm+tC5j689sjXL1bbQ2
inqUl1Fyp5PMFupZlwgMlYxXqYiLM+Y1+wA+ERPxo7fivVyMFZj9r9q9wJKCuNxX
QMzN5NmBCiqFyQNBfKsuHxIo5IbYwe3dMy6WhJ6JPpaADkmVUtEXMrgijbhuOO1v
1GhxnjDGziNeEtIV0ajKdqVA4E8Vt3pr/lT3aMnztLxk8+w3Qo/SbzhAdpifrPp8
hfgn8HULTY2oUmxgylLzPF2G5jC0kAE2BbpyhXWe4qFi40+FgVWZqvE+E//z2ljx
PXWbPUrtcX36aWNx0YIEPttkxOno4/zFcpG1gG6IdXFnkGGU8aLSH2sPO/h5PQ9S
64CayfzhvmlIZudNIq5HAvZB14hRe4HbmyGwVNwJVZwnDRAywlKnzejvsSzhHWdw
VRXeI2OFh/R/1lV61LUQ4LTW9o3/Nfre+JlxS7Cxw0o/tVcL4ZfiuEhvFiGaNldf
jlG022qpDRdGKgXK/DzGfuh6y/gDi8ZmvueT2KxLJ9YyB0q/RXYyzPBIh/tbkh91
E7x8OrQ/zZ61nIefcaBepybxNDQjzQfuD7mGRavtLqJkdDLiDzmSSFocKE4jprWB
8iZyWNR/a9lmMuyyMIKS89kt13nRvQp4DU801CchmKyjisou6L65xnfOLp6YvQ7V
6rH8GG0hQ2Lsdx960a/DmLMEFsgV32d11ZUg5IBApuwP8CULXTcl9LSUEt4nxvqp
awMNntDN1eGgUrr96+7oO59/feUGYF/L8z+bczr3BU0lno/OcGRwFLMh+AA3NuRr
u6uw8e+kBQuVeFmkVWI48BWtuMtjAC9GPwvgKXXdo/kjIvcQ8GQSOTzb7Tx/0j3U
hOfauY13eh+BOyYFGVAIM3paIkKw53WfBq9ourPyljbCjrsPHTDRxms/+XjaxoRu
W/NynxDWX9U7GNoYshZrhCwOFQ1Rcis6eBTpV9tCLiKkViy0AIrgURpRavEXj6+E
VewfQ0FJWRr1WyXOhplOtIxrl24EO/ZryiZxag+VwbrfWVFMF3lAVkqB9npxF4E1
0jL/GZsSCYDtuD9X5TF65uIAcFDrNuGmRiJoSdnUKXzsM2I8Hr2/oe9oZQl+07DO
1a26OI2eE1/VilzecrRuA/PdNQUEsH/RchEW88A4cahpKYf3G63Oih6+a2T1Mj4b
Hiy3m1WCEu+lkbZmzZU/a01XDy2SXxstyqunQ9FBva3A5IDjiwZtP2EFHRr/+O3i
uaxTpe6wzdDUQHrWbg1pWf7YsoZu9TZYJeipKwJucpBpfAuQ6fZqIX9xF8IMkJiN
CAux8mCJWO1ISLhxcA0S2ESOHp9naEiGiWBrEZCRlsGzT7twBmWz5mu9KFQ6tQY5
Tyu5DoeQI5vbeEEcyqjXGGA3wCFaoB2h7Np8raQ2OW0kS4sIVigYm/MBikz9OkQn
01b4SF1VlK04+GifeZyuYYQO3uWu/3gsJV/ytd7wq7QQCvEPYZI8A70US0hdIRUs
b2JEPLxofcDGZCLuuxJIH0QZZUA3PVLa5fmpQd0+5Jw5PceoGybVfEdwxt1qgQVI
ZbvQgIKtbRW0L2QAbRjfEyuKqd48VU8IQKUjCY8BMCj2NK7n7eHIiEuGMOxsjNXL
hgXXxZBmv42CcYr0+oUMf012g78J1ZI0qMVbyIkSF7c/Xgp67bX1NbGVui7oO+Mp
3HDWlB8OvfEwbTTlkX0vuDoH/mtsBT82t5Uygyzr0YgQKNJR0KbBD2stLT771y+3
F/GGt9Gse9rQBQ0H2plkDJHFw4cRUapzOlWKmteSefX7rdFgZUbLjTf5HWcdPS9k
NNF3jxbcXwTR8SAkbgo7ZJ9V8YScM7SaJbN5lT6Xmfb0oebAU3CsZUqnmF8WRyw9
QkqypqRujJwxM+XvfPS3Y/F5laWSHSnTa7g6mMaajoFh7nK3bsr9mCeqKA9GZl/f
CURyuappB9VRRDOjiVu9ixvFaDlGA0tohXT2rVFxspl7zpwjSXN8tNE7AjSCaycs
4Q32XvlgwR19FDkX91UIM8ILhIyk8tKheoC97OdjM//be5BOgJm/kxgNy5o6zo3i
tSMecm+/25qQym4TxvS3NRWCnLw1JtKImt5olGnhtBE0IB4CfXsrQQ/U8JulunWW
bPgpo/IKDTuvV2t9SG7U5peVH+mpFo19vYB1Rl8nigm1tmyhBmVspqD4mc+rkQPH
bR4F5FWksYipVCAL4/PSLzRG1ZXPq0HE0TCgie5RM+d2Oe0YtbxPL16t4ZxV0oun
cuAjdnIBlWaNqDywAnl51w6fqjK69qO1+13ugHzisKjj2x2HB5g9wmRrzhwOPsLj
4C18tWt7ynIEhHHvVPU1Y6oc49e+sk/zsJRIpKEPQ7WHw7kC2JLqG1pTS+DYScDO
2scnr5XAkIaji9QzksuXEHygI+Ds78bY3SCVl2UeIWJtPJrv7fKkuR1w/c6x+S9i
QKqjeq42lpTpYTPOLhmg6KQ8/OsNjEMgYoImflDQT0jFK09NmmOMcFjKs+7MoFCr
J3K52L/gS4+RgGj7MnTCu9N7oXgKvZAtkfEES2dumD5nBxlX7M75uDm0GeIaM8sa
WjVlmUIYXIfBi7htkbZL2NQdusLQ+Zm1VIvPlSCggmxnFqpx/jcm90f4zzqSwUFo
QLYeSjKvpdg77XHsi5o50Eex/g1sj/mhqIehdq/gTIaLo1KoIVmnoXv/2a/HgKaD
gOdSs+n8v+xYhVwi/cVoI9tgt/SsvnY4NJNZa0Il+frpsSapJCMdg7Ebr+1RNl8Z
yUibenSz3JzEuKe50Nny/omP0I0ZnnapX0dRlQJ0a4WwbE3t9JcZGVyLhINohUKI
ra8xR/jGS6IpPOzHxuiRHY7fIXu0z3gWtIXkOKNVbWckEufZ21WNSTukKjDLuIVv
Ss/hgmgv9ec0QtajHUncqa641UJyT/p8HmqAC786XbRLE63wwQCfcYzMHXwACvDR
J2DP1tUYxwd0ZSzkBDNhmh7ruUhTFzTLZ1Je9Hg9vV6XMMt9S/L/FTKZtRx+EZ9u
61LPXHrh3Zzd7pwzQcvKq3s2iThuaO53vmpPnKN1zsbYjuZHXLfE67hVuMVpqkqv
+v4FLOSy10eXaTFfktoXHqQSD4NE7culV/503p+ppAtGk45g0fWPiUwXuf0iO8b9
JVc9oAud3Rt1OPr5dNT7EfVjW7jYuJNxd5zgn0hVYIrKyrMQ0RBTjBpcgYq0S1T4
qUFZbwrMQAgnj3JEJHhvqKExmPQR1e02WkfLF5Y/bQ3t+njDfvssvcEKr8al50Jl
1vxvByrckj3wLy3c0Q5EqGMwQYVAGAXyM+SnrCrGFbY5kZRNixFoWKg1IjHqmbjm
b6J9CwpaX/Tz5CQCp03AzMBkPl8TqQ17nqRqX/c+zJdlI/b+IzaKHIlWqAdwIfBE
cxxs08Cp/x4hNcwG+lqueKgWXlD3UH+syzyirNqoqMA7134czZmmN8ZnUM5ikIcT
N4bAckKp+TFnekUhYKbGT3WCLA+7P2YyrLFVcgiVHRYpjkKY85TZiRoOXajRO1L0
Ex9zOfzIbI8t40txZAzfVJa+tpZlEJ8l9IKRrN8LZLMAcipfOBAan97ZkXzQvtk/
xePTEmDBNCGaE8NcsIBZG8Ifa1GRBzK1juNSlGZuSiroKtsd34sE0hiqgyN1pxHL
kv5/tOzMkpqPAeB9I06oTn3JwxnQPUo/0LqjqmEJ9XRU9way4pc8wsuKOCSKBSEo
gd+G3BVgLKex/5JH+E5vcjcWZH48+3W42a0D+jf96/8A+bSJtmFPJ3B0/7n9PqOP
+zmusyXaSwC42iQoE/OGug7QTgwNgD55C6IRw9E3NoDtMTJ7obLbkXsBM2+ts8cW
06bmn89oJem8MqekIjWNO/VEjh1R8fk7WNa5r2HJ5XIGAlAfdhgDyX69aRLB3XOG
VTNWgxCIXJ5l4FRqiyNy5SZ8Jx8oxX+hd0+6txFbGP3qz47rT44B0+zKsDo/w5RK
VQilZ38LuyycdzCrd9m+l6y/eA6/91L1rgQX/nPNY8Uf/tiF38Icqc6OkMzLOoPl
9ytKLsy0z0Fjx8nDgMK4S9Kl7fwsafDS+2k+Ew+t196tlvy5GWEu4cYhRAEt6wl5
K7kKd0Ox1rSmLt7NY7CKviuvnEC27UTvqdYhKw5DUyjvBuqI4PLYSaZEXXDYdxBs
VgCXp0NmNVp1Xkb19QRI8iMQch5egUSaMuFORbDjVaXfn2iT5C8Dq/iKAP3j0leR
vPMoPisdY2wARl8viGdxTXAfAPQyu4xnx/2HvfavgFekN9E/xeqt1V5McnrzMJng
WeskODBZJiObJV0I25NatD6rpNrcO0vr5XuDPZOwxAZLbkO02TIXrdPmSs1uDHaZ
dfipRcDXaSqOSQh5j3OFatMDBHq2Flw6p02LnfckvSyDE9IsozGgdB3nEdPonqL/
1u7bES1y6350c+FVsEUvU09j5jm97dCtFmurOUbmzNsEDhYhZChm931L7Aa7vmq/
Jr5bUmkg1aR2QoNkqVM60Y6X13uVE/RHbKCp0AwSeUDoG37Uv7AoJy50x4mNzoXn
O1qVKrh2ZFJ7ZXeG2Y0RgT6Ko6ZFbAX7OGZCto0ZJf+VyQXqSvyvd08IMognoUqn
4cAAUUeZkwEZhcFnbGfOFrnRUu2+lbkdJK1EREdNGRjBIujGWaHNf4qzTUNIFACE
RDSy5mpk/yGFom7FY+UF3OVanzRlDM0qIkqKxfHwo0n/kUkrEqpLe59ITTHxSjld
UFtnY5IrrR1xxZM4X30r8jVD+1BO2Ls9UCBtxy6HiBH2hVYqZk0QJ/i1+d/4tjZM
oML20AwccXq22Qr9RmFrumKHUbLG3yK3bBHeg2GRGB8Ozrfjid/h84IZeZV+Dvzn
CxSokslxWGHX3V8NLSowJbBrvXlNkhC5dT+5xc0DQUrEJFG2IeWFTJNPj+90n9WL
I6BHbsDezQ8z+z4No+CU/km9BuVtF9IbiHh5dbVWuUHxlwzqzAaeWCE8Qqni88XI
m65lCP2DJYHxqWLfz5xii/6d42pySdcQ4s+4DhcF3iOCkGUUfaAb5s2nAuk8p0u0
KrKcc9dyTrM+yoU2tJauS0KH7DhhaVQhR12/IHs35MRhOBNpDvlniWQBaiNBkQ3D
Yng5yWU04B3OdcH+nG2tmX3PKnrWukbjUySs5OcYp/EKNMrKUt3hgQ/hU4PZ7t1s
f4OJSn9NNfJ5vic5eLuX8w6Qnxf1U+xWdCd6qF/EiuBYjkb5bkGFI7+5aEsdgdKD
tdhVvTVzI48lhzqgAtvdrAN6hT0jAS5iW3Xoc//S/WmqH2tvS+OBLM92G2mAiFKn
6Khdyz024xmh/5ujEjmeQQfheIj85K+BABoSdbYHS/xUXhK/Iu1u2Ve+aFj1Gu8P
HPvs8Xh7mMo75meaY5QM5KoaGEzotGKXr8lDHUubhFecsP8OsrAZmK7mXS0kIOXS
O6Zu7nBHkd/nxOnwUgIZtegXH9kVlWvO4mudE4/XG56LkjBRZ4deQZ+ZOtJMQLSw
Z7Upj8x1lTrtPm4xasOyVRL7/S5YZYQp6N/WEoxpxAEnrHYbm8bhfHNQtqys816L
fOmZ6y/HyvNHxVzrtzS/acTom2fv7sDlMR93H0afeSHuqyVUxVvNCPkWTY3MN92R
hnlp9FOmHXRYbuhHfNx0ZguNZMAbCuCichP4UMayZT3RAt9623BDajQ97QpleYFP
5fYltd+vENB4qNEpQeUkiH4tehzWMNJ7KRj+eTkYnqdP81xlQTM12md/Y8F91qva
BajEC1Fep+Am3NlxA672j0VaHfjrMnU8W6Ik1AI8M6o1to/PvURXzjYM1fxU9SHu
2EGSaU7ax4r8lfJQkFlpnCCpByGsOhOjH9aGrUHFQ06LbTmiIDDbNrWV2HvHLFQU
2lI/OXWEzZ6LiCEk7Bb36I7ipzcXRG3IIxKrQquNVFGFifNAQG7J4jCgGTIjf5OE
0obM9ae0XKJ29IMfZNV1BB6os744dcIO9a8wovgFKp4ZqcF4H7wZtjWtQ4yXlsKu
wXMibGnGKro4FZZhbLlhTL5z+Cl8uau+yA7dOBTs+wjOWjVwBlvjSJfCTNfMJXQ3
22jVUpE3PdQeNHBlORHcIlw1cuM1xxt/he3dpb1vppSI5HZLnNPNE9tKC4H9Jazr
XINu6e6BIiKSwZ06z95ik3942FMsmz4zsIRGtCxAu+kvBEn/TdGQIiQnvXtN6pML
j1u+K6xOQu5gpnhBuF1AocQFVM2uZy24z5wWnGAVvgUDjCopbssv14Z9VYEstueg
+qquP2I8yDiBQ4vXl3PFUuuM22IVQ0Fq7xy7yCnviQQLnht7aWRSZt4kHhbjYL6s
1tq6xKrb3jKvMxGkUxS19lCS9ktdshJlbihcryiY0lw9inD8LsXPMGk8mW5pI3xc
RBGzAqdtHtrP99dgF5M3jL99oleKRZOz2TtCO6L1nUrIVEUTK10TbHMm55dvrAdN
QUi9fX+gtF0WopkZzPINSIG6GA/QPSj6r184EC8eD8Mj+Hrn5LmfnK6l8j3CIBzv
cN8NEjtsR6MRWaX/FvEBfCKc4cxU7jex3Sgje2flMQXmglOXLRUssjh7zlv8dMZD
SzCExIGJcq2KqzWITDvqjVx3Rj+GZg7AENmBVnOFZmRU1q/ah3nXdf5QODQUjw3V
8sfuna4GhD9KKUzIDdx53Yjg1pLh06s3w2e/jrJ7shIKnaCSp5HAh7tBlwyjTV/r
yF35Eq3MMK+bTphjoDu0X3YyH/nz0/rsfcCg6wIhJFgFKK+w66BSkIKVvEfKYQd1
pO6DQkzWXw5zUHH2XBWoQEbASFAe5hZ4lAwpJTFsr79FRktASL9PQwhkYGT+5UU0
PqsLBTZxy1CdMaZDuecxwDuHgZFfvh8nENRgYGt8lYH8tJEGUtA8b/w7QW3hWDOm
45JVs+EnhKhwQOU9uACLXBUG3aFqcRa+qZmVV6vc7irT3T1hBRn7Sqg2zLSMyhFW
TzBXrRbWvfY8j2NjybqM1QVg52LA0fhLz6DX/ZtKhi9mg8plYFa6kpnJir9dEQOz
Zbc8brj3/2i4NmkOc6ACDzKhDxLT/sE2PuG2vdF9QH9z2ZNDhcyFgdCADY2yfirX
6wDDxo8ZMt/tpK+EF8F3gp6/1Voz63EjljNtG9rLiz+R/Kiiu5JGhIXJbsZ0Y4UI
6gqb3EwSOHB+1kHyX+LMHGntUcZp20+OYLTX4otN7zKMtTzRJqevkd1ITjrtNunO
lYX616HdkthYN2Qm2tpDtPgyxFV/MM7CcLTzqTtREKtskzE+1yEbpOryYZRGaGOh
2XULX++0RdLQH3FzgFG/Roa0BTrgxoDb3/9V2SdNEDQOkl51hbH4BrETUvQAh8cd
h+4IV1PSpqq5S8QJLmFZlNwsRvUJKRxeqUHN39H1le68HDUfjUloxK2qQuo4sJ49
kmj4LwPKLE75+k+LVAWSRtqZl4yzN1s9/qWrFO+V+RXFZkPRXkAoZnsWVi15713c
IAmSIv8mSML8G3WQvwbWHXsRz/XF7GuUFqlw5HFyMeGLSNSDC9Vh0SNwWmvW35Jl
ayF2z3MSJF9LZd6g+5gOXVAnhnZghMmNkai26r4f2OAYHZNNTc7krSyk8R18kMyb
YHYGlwGsd7u474CL4dJJ+I/SMuHZkA9BBC5mUh/SNvXl3ch6b3aeBuy79TYxeSE4
UJ+4/huatxxCvhzVmbnFKu8YhuQy8pYFUPs15NxuD8VUlRT43o68o0UmNT2R785M
IZjFHaevHoy9ay2Ahipk8fuaLQboPargIm/8ov/syNo8xRbz5i1+Xa85HJVAP/6G
ZaZ+g5az+z8a9tHNAsapnG6kdo/tlfPG0lsqAR4cW1D5oMpl69pPr9zhi3RPgbuF
LXvmgHyyWzgtL1qsAqwp5IkY7pJDGtiwqOVrhaJXArCoSvM+4UyfMRv4pOKKHmo2
UBtJtUwVW4uexWLMyS+WuxtUeD0a9r+2tuJDVIPfZnW3RTXy/+wi5yrTZhnveOmj
Sj8ad2ADp9oNwLkAYxfghAZuRozDvSIZlTmwULZ5LS/tTsSE44rnKDIBjB6M2Ypu
THmfCeIdjU+c2Yfw/QYUmBZ6z6oDMX0AIW8C7gnqsjkkEjNKF5vcGmfpMrOnlYu/
U/FTc3QMwPTtWqfuQrHrGsV+ytvMq0+IHFCGZITu5xJjmtKYkRfCpJqNtHNU6Pkf
SYPqYe9QUSniUq0SDTePXPkY0T2rSq6Y4OGJsYtDOXyXy36sTuBi/M50Bws9quNw
N3uGURNjRfuf6/96zLqu8eJBUb5uStq0MSiaY0Y5T1r9Sqsx6T2d5pGlZ6wZael/
XdeFWyNOKc+MNSXZLucLm4I110cXPvGfP+6MitMv1SEJi/0BLvMh34KtJn0wLvC+
igaF66foXLEdbdGYIAEiQeX0+ivFfcpOUr1Y4qYrAZNSOsT/og+Ekks/34pbKoyK
Jc6fjp5uRO8YEV7mWbmoN1YD3r5FwMIRjBEFDYX6v6LhhI+6lOH+Qo4PYegyKU+1
U8Vfd5m8K8d7Gu3x18I8VKF3wAstaoVNmAJfWtdZaQc4I73fQbXfT5yf9rmDJKzH
1oz9Fl5jM5RrjQAID5YegGdlAxrmblvf00e//hV+PEwlpHvOg55b/uMM/bD0APai
pBB/kfZXc3CsYSYB7UNdW0kbD2EpegHKQR5va5nMhqP3y3uZjFIMWXv/wPwWd2aq
rx2PuZjLxqBR4zwcopnmKpLvQiFY1YDhtsdQwPSvPSFS8Pa6bVG21GkW0MIDXkLS
3leHheeGoiq4fAmTo5JAe8BPUPZ/9hKGLmQ6lbGFrvAgQF859pEd/OPhNgfSV4MO
kLgBivUE+wNOSwXEJv+zyRuJSLuEOU7C3vG3p9WrBAFH4Oe5ovXEPcuhiZNQNpnx
8n/p22/07khZ+jWUIKg54mDxOjc2LigCQR7VlSp40nUJb0Avy4wGyZ5tzhPA5IJp
R2TblVlk6prkoY0f2mV12ZP5XEvGvy4Bq1qUcZI1VNOIePETl5e3GshoISJLsL4S
pV72/QXH0zA8FVajNtadgUrq+cHMz+MmoEZuSCPWB+kj9wNoG7ylCNVsHm8OWH5Z
Z9qH7LBU5Pm6tjilcYzRfzzq4apMIdrTU59lmxV+Ixcpg7rVFo+tRJ/WAWqDSK0h
CgOuWTMA+jsc6AyBfZHpRfCcfZAPJLA9CpE+9/jd1s84zQvvj+Pe87TpxzzbRIhd
B0OWoFxv+99hd5vQKA+AVTBsz4ck4faEEKQt80Dc4qCkkng3T10eiuSIu9j2cWo1
2unDeEwpACJFe2IXymJKbiVW+jrklmjP3EzL0odBSJYO1UDnu5S9Cvn39beuGJMY
rm8Xyj5Dkd6PcilXJK5YBUVuBd9LIcKa9S8ZA9ZFH5YkG/hKIp+91yX3NYmTsIiG
7OnOCDM8OoYeObrYbnblycw3knu7oZiOoRIIJRbV4ZqV4MxaUOGVCM9yRAN6aHcv
FrG0FrDUbCVf5hKxMSF03sfDnbp6lG39nPbTlj/+U3Rx2vwgZLLWf7Avd7BH/hBk
yMtIOl2HdWSy27PPe+Q2m2XsueF+axYlqtyA7TzF4z8nnExEzYYKfc8jXqLiYgeO
An0xOJEJ6+lh+tIGIjl49q9HCQueldH9+8tNfuPljye9/SDI8FA52+zwJ+8ciOU2
6KpERVfjPoMqZlchFVS1EcoRDujAFCeXCNoc3RCsxvDwfGHLfpEWpDTz7HTd/Nb2
cJieCiA6oBdcqLtAGqsNyvSn6AoJALmUUAVoHqRR1IiQhurZWQEc9sDuCqhbynVv
8/U0k3pHiJHzgwAcce/d95JKxNimDcyyWImVzI89QEU3McWtuNBBOYKAMfOANiFb
6L8shzCvoWbodbNZ83ONm+N5nGh1fJJ9mbMlciPIwj+ZNKzAyDGZjv5llPyWfHCg
QnwYd7XsAS7dNZfT/cq4galRyTyPrxxKTKt/dY4D+AZsyY71DEm32BRX3uVLxuOh
NjsjkefBvoBC3zT7yjEb/cJZw8jZVn5HJUM4sjYL8jbkyXjjF5/2uW0o/3Yvu4wu
6CtwgzSss7dmY1Bl1aT1hIDFz1w2aEv82JE1yMTOgtMumFMGwAIK8lUGXRYkWZnk
87pw8cZKYnAbnYAdocdu7e+Yw68CJR5MU1X64Uek+YaSMikZEkLXu6gClM7vnn1F
rs0bh7ZpL/fK7WTOMUCvyWicVFLN+rLL+kzVMZHaEEtYRDvHW+0WUpH0ke8jE6YZ
WnXcEpRlsvGb7uKDGzlVPjznQkyb+3fdJTqYA8IucdcizgRJFokWQgnrodKcMBQ+
5VipQ1i/BHMkcGCESPuU6isRAQvB5sMflUjShFcutxlbU+Sfo8jVFu+qByRwtLHR
+zvjYjO/CmqzTzt1QdqhRNzZ0xqUgvjEHHeIe25/vlzeD521yFF9fM6vjDIF+kpM
vbrvcOBA6I9M0w1oQONTBj6OVZKIDg+IIHpjs1DFM3QdzTKuV8hyjoG66w3T6pgz
zhvjSWBBdy0FP+EwUj+wYB//XmXQxr43FIwUYMQC+NrhUfYiJjkDqDadwOW0ORMg
R8U6cJ8kgsvRBWEee7bqA2IKbl2EGyWbQsz+BVTjVDWSyyewREsqHIq+9DqMdtpS
zsD/4NUAYcz/b63cBpVwupMyuZmGt/ODZAlJO6qYJKtHv7lB28SY07yM1iMelKzV
AENgDpZ25fEJp/oDmlLt0HrK0H2/0eFB5cC/sED+MrvHL8+5MuTCfLBjp17gd5hF
+V72iKQPnLrhDjGF0vBxBT2ijD1QrL6X3l17Pz+f5ZwMdow7ROQ+muineOdU9YJj
61MsDdVOrkAEB+DZcUmKpWCt1/m2BqrqDhbILZsCYjg0OKEE9yq5FOoqWzywHgSE
LXjyWCE1Km+pJwe82oxHqOkt5HwV9gDkp7A8bY1a6Z06rZ0wVPVjqQE4MDC+WvWO
95qoJEhNbwxF+vahY6Fb0OuhKv4rFnvTu0V0gAK85GNwFIwrxLTEPxbBovdhQ0qk
SBwJFknDCHe7A5fIYEjrFE4U61gkAkMv/mbang2ivGyhDZx5exQbLZqBC5Fc0t6W
HvOVdCjPRpu0da27yuOpuaOdl6209ylceVosMol4DNP4wRqx5A8AyD6g9kRxKIXa
hoU37twjnWY/3WTRTqXd/yrnYURi/NLX+sj03kpMZLCKn97uvB2vy6iJ+6RaLRG4
+lf3Fs/59OFq/3+YcooptIBzIjAOLLrBCBnq9xhUeSgYJ0euSGVkq/Ry2iP3SN+R
/e9jKubcBykQ2lTGDH7VmzgVVcngLSZpNECql85ufZhWzETasdHcAJ0tiGoA7u34
6O96GR/8iHtnRrBbI3+iV0zCSP7C7ecsQqbVwpEI88Ff2kI0BiZ3qfrfphGKc/U3
8YMo6Is+dNP3lKeRHREDUBA39duMIFn/wC9XpPFYhBg6C63sR/kt9D8IzXZb+dLl
6hqUfCYYsjXEjkXARVOy725URXiWYkwCq0drS4z9WXLpTciD0KpK7iH773ECgpga
L4ZHctpG66Pd4kwranhH7dahdm6bxn3COTOK1zyq/Zc+pZtEK1wJHv3GEU3PcVrx
c7agBeHky9RpYPwkRS0ejAY4mgdKujfABv5DhjRme6jdj9JFWvc2NDKQ4gqMgY3p
AOuMmnwVJlbGW+ryxcotl/3jdWZ0e3RJdqifHa+gGTnga90ieggYkd2hH8iye1ok
ANhsN6/EB3U6a5xKKaiTgZsEWfAIgGiB3Aa/gyoWzsbM39EXjGD+7P9GSytVg+Zr
/BEsCuV7azbYJ6agHO1yRTQ7ZQjr3WIVSYCb8XiYpHMYwE+vM6SxheQSAs6gQGvY
7IEZVYkDE65QMkgcE/I9pBfAX4I++GmQGPVpyp0LyGYnHf761YZHQ3Gqh7eLJhFY
hlLweM1Z2b5C2pKazwL8pVMXLTBdkHdOuQxotSFZ1MPc2ANjie78e8Dtysh3vFcN
7TC7rPnqny7KA5qmFJRwm3hpnpTgNQEw0RLm9TS0MPCaIKiini/qjbtxoIZMVriB
wP4amuKzvNQ2KfLV1hwlXDlkkUupDcbptMGN7aWT6WHUWQwsQXxUc1hPEkSMmbwh
+CVq2Rye45LCgdJ+Lurx5r10haJFpDAg2JOeQxD3UMWhCmD+bgL9U9PcbpGSbgWd
KwL+Pl0OxTOu8RZyYYQiAMb0LLtN0vuH2B3RcAvsNFk=
`pragma protect end_protected
