// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YZAP3nNeDWVVkMffTUFhi37Lu0zuk9i4CzUOhZrCJq1LcrnP+m8Xp88WDY+y4wMr
amVOVfnVZOd+DOw9Nsy5FcnoxXGgtnIM4GNrxWZ5wIaWbrUi0zCwv7hb7k2rTZ4h
lVYQfmoKfyGRweWyU7mPTKj3OUSWj4r/bhN67V3yx+o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22784)
/MlCtpkl+O9H3MUgIFaEGeuiNh5pH5D8IH8raiVTRY06HE7KN3KVgEn2vrMlrqOU
EFR3IKkYO/qzzVt6OtSQJF61lZ+CRpu9fmoi9CY7ZBkt9u3wJSIDjDxiT1ZDJnA6
GTmYdicu/yE4ek9sHBNa7jGZtLPJ7NlI5bxRJDpIeBDOAmgKipDJqaScOw95UIgx
wR6qwfSmozeVq/ijLSSuNR18GqtmoH7YI2x+CWMaWR/BZkrVUvAA4NZSQIuEPsPw
4mEqPty3tMCos11f6hgb+sh4KeRbbA+1Ev4KqnCu/oiQfyPqMu+jYPtoT0YurNZw
4XtUzFOAsGcnUIo9cGuVwm0oXW+ApdVfHMDK0uUrBhx4NN+RMFCgSB/91/Uze/hr
UHW6R1C66PNXkyrjm4KoKmuLfo1+QOBXGk0JUSPD8L/VDh6mfx6LqFdHm1ban1uT
RXGXHc/BmHScLIMYxpZblxUpuPe+2vTXiljOhwPWaeqd2Hdy7F6IHvuJzGal/4Ko
y77mcA7s1x5DfuK1NPIQ93KFHoP2vMUi7Ys+dw/Ggzz0/Ws1rf8zGe3ElkZOLjLo
ZTGxS1IXkNxe6GJmGKFIj8kZWF87Cr5Pg5KUzMrWYtbHtNaO2QJr87693KD19rYo
ruP9agQWydeS1jQ5JbxPl9ZXwt6W2jrkv0OJRON2stzXVHA+/dBhX//foKxInF3d
0Wdj/QDm57+dl1ItJQbn/8Oiwhuu7io6VydK8Ye2QP/Xvz9DiYBtm2KZQay9Nknb
Xxo9SQ7KnLAhJi09oe19RQdwCJupj4hPnkOsd70fQZHMJ1RzKW5OzVUIrMZdnuDc
rOEc2s3yPxSYW4IV8fuLlkw7AkwTJkIEyf7dwZT45MD4tIKy17RRdPGHZ/iP/zCU
Kmf7+swBe5JBPYq81ASHihZxHaJxOosrW8nQ85LgVrdYeSG5mLm7qLas+zezmRzP
b+UVIiN1xsPh1jt4NCJMToy96JbUTQR3YZhAVejnq/mCzMgBe5zIvg7W4SrGkGXw
692qxLorh/lHytr8e1qiW1uW02Uha069hYKmAV3xuNYWD+AKvgAeHkJJyIkqZyVI
SlEFE7a3i6lRnBcxpBLs96NZ4dR38DUxedBqBaBnfmYYTv8IgaEgVgzPRPsoVT63
WyXwyfEsJDcUnHY/6MRdHoVG1cvaySJD4iWEiegHpEotoYaQZkFqXvCkGOBelO69
A3+HIZe+cPkXcM4c1ljRj1DI29uDIgL42xolkvmZBoYvdbpNai3NgIZJvcb3/2wE
ihgKtaTb/EClvj5hi3ARKF9k00tDBE3PvRWbIJqD51sg5FBPt0iD4g3f3gS4mYuR
TqNCJuQ4p5+o7HixWcLgp7N3+S5Zc0bRUYHyn5j8mDF20P7dpeI0ffGh0NUh9a+5
kxaaYUW3TMWeh9AOAsG8klsXVYlqiRJWdAQ5C1r/JwywWSRiutKQdNRAyxuQCWRl
0IWa80Eowz5odCziMs4JciFa3XC29c1VuCE6smln4fIOFOUJsxGzS+JSkCvgp65a
/ATKPzkrT00xwFhEZhiili+Ur+jus3xbGyY85TlnwaZYDAn9B8Pivwp2Vw3dPizF
K2lz12fQVsCm5vWipBOhjuZrZ1QQX0Pq2ODTGBR6nPHeWw9NynLF36ZUvtDVBIJQ
y9HZLBYG+W77J+3dzSjADX7DfztU0t3Rl3YzY0zkOrHB5z8VCVB32VNu9CnfWOH1
B/FgpsBkmvvbftwtmnDZ/oOtHDNCM/EJ3t3UNk0ZKBr+zJfwgjfPTSXGqilnbGEB
lXVAspUjNUtMazfhfISymVePJr1D44/Vf7gxztoIzJjd9bBaLQJa2QrKPx4gtPeF
j4OTsgMM6bHTpn6H3xlEjJJV+TP0oP5aTPBx8GEGqgwMjGgqaz26yOoD4Dl909rA
Hqy97u86ulSTrHyEcdZRFPXK5XoJksc4CI7ZDPNHsyKxTrkb+t8x3brlpnyTBlXA
QLT2FQeuLH3SZvpxTRosK5JFJLXL5USJbPTksyTUSygAzOe4BPqYg7/MgykpM8vo
TV74cHJc86jhe3riZ10rb/6YrHza6ydAbHcgC9k73ktWqdf3szgNFaEjID5wPee/
owP3POa69jqNWrmQxf2lYAmLKS3KqQUXG3BTlgeHbH/W6olpqsIpwYOW6UqRTkwM
Yl+NOeR9NIsKTNjSf97xkGfLYgSXMKliII5Ocs7obUwsCssUN82/jYbKC2h+Gfwu
jT8j66AbXLjigObvZsYuDe8wE1gMOPvQbojZV2Jj/ji064fofq60XYG9JHoWWSVg
6VZ743JmIpCDEelCQ7VCmwEfo2cMDA+ZosHEGO4drQqnPqj3YJwEI28KuEJqWe6I
LYjvQrXeOxIKt/+0UoCPenXW6QwpMFOh6UNcWeTtlpolrJL+VXciRyDXUglYvquG
/1g59DSyusuZUpDI8+R5i0K6XB1+4Q1Q1d962/i1roMisI8UkVtUQ9Q4QXWLbUyC
yUbaBzFX7XfM8i7HDcz6hONW5cVWDA/3U9kQIsBkN25XsgbAribkkeA+2Q97KzZ6
ulVS3HIfpOUqa88GKdpPVpje1CCsifQV6OOUq+YMYzWqbhfwnphF++N+maD8Upvn
jW/F7/6xw8X6V2hPtLefY3EFe0tBnqHgMBgVUgm2yEOlZxJGp3s14LSW9iD8OQKc
zGeSs3/EsP/quR4Vw1X2D13ad5xH3E2rpIHE57qvUbvjied20rotIU9oaknT1Aaw
44d61ZRtva0ogEtWz5cfhgnXd0uvanCozA9UP1+BWNm8B4ou0HxhCBlgRRhVaCqt
AtorBRyMjhu7Me0BWFsEFy8Gxjd7v2NCYLtl2FBs/cXZSGhheJnLA1EmPoUT5koy
UXtHU4zHtovjlUPgtz8/qR8gZFj7ZX/cltm6OlnU0iaqAJheuf6aecpyz0su1Utq
R85EQRmRdG5q9WLDAtCfOSZoe0nRmti8msRH/r8Y2IyAJk1vZhqMcCTI1Cm5wlbI
a7UCrmLmKZnU33kL4uYMi3yzC+5ONufQllD29bmkgsiBoXemr8/G9jXatndJexeL
jhk1dEdlCYHHmxsUBzFtL1WlfXIJgpDbIdX5/+p3A+Wh4c2SsfwWLQiUTwjPIS2H
uilPGSQXbU/mNEeYxkxNeoALCrJSZmGGklcU1NvXw0koc360ykT7C8yIxLz3YR4/
LtGqE+m+MTvEkjTpQUz67/QORaWkvIyA9LrrG7O75d1UVBwcxcIxxS6/RC+2WCI0
Y7gYxjkxeVdHiU27nDHsIzg5hLIfdcauxbMZp4lOnGDPQ8zo8fVXyBfBdhgVJQ1p
TgUaEujFr33rnIangUsq1/62aSQESPv+2hArDJUiFArAVFlxbI7iGbhSu9pxVD/Z
siPRHnEhB1EN3Q+j7xK7xP5OFQTCJiOx7+MXC9WdMnX6yqq/yWG8PKkGCmyW4Bm5
z7L9kgESjNJkIpFu+F9ZVeI0LLz8G9CxWn1W65pyBOXbHgXEDt7Hq04OxBRg0vKR
WzlgAzU5Yi0hDxQXKcSU2izeefR10N33norEPZFAvrP/2mYV/b+edBJlmhqNkVEC
okpC0Kcjr1LDJReFro0uC7ZwzYEUI9q8sPoAJQC4y8cKb8tiDFuxH79XRdwH8if3
DiIxq0A/Nt/zpXd/G+2Pab4TIzDiKID7dArDyXSyHziAK1cCvJTvwh/1ZAbMhrbV
G3gy+JvZPjstIwe9ZNf0dIpozdLhhJPg7CxrJaCNhFJjNqCn75hz1oBu8bl0bJli
qDCzcEmpFvFMly+AovN0IhS6bx2udeDb8JSRdWH6X5Co2d+iis9ke57Pp3y+0KPC
Re74wKgmNKbtuflBo9eOj6pMDi6Lzs+Yx7e4WCl95N1T2/TQRiz4My/sTWZhJPCy
8b58xzqu8B0rn+Q9Qvsl7t8GdiJj6ivzFRlCVGNtgIUiuwgFh9D0q6hI3EuaX35f
EbGHfQUPc1R3SnlnV1ULJwUiGKgWjngZxgt6oDlPN5Y2YJqbKIbH7GRo4jQexCby
kgBdaSEuNMiqnr/PIDB4hHpfehsq+CdgKsXJKNmnj4P18RhfYTWGJxF4CZKPu/bR
BMRK25jLuilS2Y8dVWTUhsHJK6ECT5acehIO7yKIvY+UrCmzoZ5OUibcuy3d+hsh
u+saXSb66omGBrV47EeisNiiXB9tC/chXLSQdfQwcB/gsE0Sq7OHb+3zcjNSFr9p
Qr3GINNtZB3f1eS6CdHHfXmejqFa8dpseFxrEixunHXpyex7eGqAlTpcWP6R4xMC
ERNvYddNAvm699HCtkbl0dd9Ob6fAGNb1lGzPjnFrVYAbfNlLcaKJwAO0YRQMo/+
BL43iWdtrH1GlZWdfCADbMgkDk5CoRT6AHuiiYnOPZmYvOv7yWLFnxwM5wt+E50T
D4+HGew2z/iWzjASAnBnNnhQLUKecV46FzYhX9MzkWuei06YC1Uh0ddwbiwW5MYw
XwFrtgFJ5Xxn98nBm0U+R1me/SOotRg0nENBROv0OdxOsUqH9l1y0Uij6i97HzNS
Vl1132MFecGDdtyItyEI6F46IzZb8PRIZIPFeGkIaEyb+wUFkrmB3Gp2vb2otbQD
/4FcdZdkA8X4LTPGqTQr7AIWzDPcV70cf2Yu8SsrE5KDNtsYPJK4F7T70cXL0stK
5YpdVWZ+cS7YMjKVW6IRpGbbb93nyefGyeb+6ziYp6IuiXbMRtEzZJ1UyP8X1zRq
7nogNEfdstXxzp2cl19XBtTE8mLNHL5p/+F4MzpaOPySWkg+qPPDIiljtsBt2DJI
WcbJNVMTG44Fdjfv3lyGKyPjHUiydnYK6NCppoZ0VLdY4D1Ergu9V5rUHlBkiq0G
Vrdazg92ZpAfPdKoSupSwc38YJPnEAAlwz81u6REMEfRXwR+GuLhghtWz3yVF7mw
flswNQAQe0L58uWGLgiSXcBefZ/3p6UyIS4ci/u9cBKpgr7TUoXRYTkGjZjRM/bg
6AmQ1AY7QMrpN4Yz0dE752zOSVaYpZEacWmdpuCtKk4pZF6R/IhX+TNhwzEcipFY
B5WjI+vWwvkXl962Wf4WB+U4crohit0vXyqokQ1HM/Fq0Z5lEFTyzNqCTh/WuTZC
5NczkoBoaV6tO1JamCKzMspIzwTtbjNIUgBGlHMhfmZlVVabFayjfPRFcq8SjTaZ
q2ttScJiRdjqutWMZA5gJv8GO5oNT9r+KUrM2ia6my0kQ9LXnimwHPWYTbWw3YBu
7iMZH/ssz8jsAVVkHTNfRZwYCetRtVDGpY09uXX53JC5Y9k/9KgmEY/se6RFKo4e
EqPHpu1oWFHhjWi0s68VAYrJxmukDLJy+G7uCX2AjxMgJTSVDy2xa1c91qy3Kb+k
EjbITmc1SOXDxjFaVpX1fhAj3cEOTbrzwdq+10BnllT5RsJS+oxpEU1zxqi4bOkE
QpPLtaLUKzNlVZRhXzLDNpyvPYPm2JwM1Lrs+1ldhxeFTvQKZotCxPCSXJWN/5Vt
n+Jzq9VQbohKyq2jgPH4HvthegEhMO9aVYpyN3DbywUb5hTeAxrLnkd9fc5s1OUm
hFc+s9TdZbzp+f+IwmXDLFLFnw0YjwKSNxIHsMUfUoqyF6a59wA/xeeSpcTHrMgK
k0pYsC172YgpOIh4WsmnIdMcbs0Z2QSOHLqufHvLVmMRqdqq0Od0znK+iOfhpYm+
80n2sJrw33IbzMQHx8TvnO1CIGYsoWKEst+eFOYHuflTRBKyDnZtJbiwppmKUjgq
fElHK+AtxHXaaf7D8qUZIujlc9qgAzDN8Lgs/7gRmWOkIHuRG+FzAWRVpW+ktrcD
HGZ/ZPrZQJpfVl1TZBs7hNOzUZ9UR0eA8mBXPebNEke2HEfuDuYG1eBppJb7kHzz
xQlXsELWWtxcb0NuOfQFEvCH0yGTNk4DKkwdm30UFFXaw/hgcc2mNYEUpRDuV5S7
8AejEwxT3ZlLUGWs9bf8YTA9adUiiJBedydyvH0Usu5jUUcM39ABr+Tm9H78sYBX
U6m0gDAgJCUcIkrjJPNfUfjC6xRtK4PVoqY2oBGGJUihKdIklkS7oZ+rps9M34LW
VVA3PRb+VjDDnZNLW1a9ECiXoxPhSzAH1JZnTvPYRnGJUM8JjyV392rCQ5OdIW52
+6qKNNt6hwqrb0QjmvppZr4kmwzEbjnYdcZdX2Fa3WosQQyKvg4lKdPaUpMIYu9b
bIkXOQMAb5BCw3LkxJ8OKJ6cKaaKgfiIZqoJheetqzxgwjqKvhQ7FENtwVOzHxXy
jZpYmobOIa+aQOL/Uq4SKsSyud+vZaAE7ifb31Jea5FXn2s828LQNrmg84sRInZN
sqV7WtTE8/kG9Xsu5dgRHy7L5y6vDUaUw2IpspzFjaBz/sibZJEoAazM7SVB5+xZ
BE+TvX8cwV8lwUkIsPe6fa6/Kp1lOifha/6gfE26h//wzajQeTW/OcLmuwqJBrG0
PUyffEc15a/9xvycfO/rEyYg4O4VCXsQZYEJBM0q1hQ9DZJwGo2hKX0xAhsdVAkO
iJZG9oDdeM+9/duj+gjVCOT54Xlep0gP5qkIDYIXcEkmIxA/5S9UQIrgLQ3yAWmZ
U5cO7QyiNE6Gc9TnZbPEmm+K8t6mkPf9H33fqcG7YUpa7kztSoxUmTfXJSjjveqq
sBZyqWZuF6QKJpk4vpjERVz+l2Zp80aLD+FS8f0HV12qWDA42n7XA1WhiCCkH/JB
uyXXB7Du6EjbXEsQOJ75nNRXbmUm9FWvX5NwYntTB7D3uHayti7Lb8a3U+XnYEC+
RMCRXNa3/kD707ooscUaQ6gWb5OEFrhKiLLOusTZBmaxsxWfS7aVt1VOcZ8QNZ26
dkaytIJu8VGMpvEowfEtSmuxe/IcY7V4LutGK8UHvwo8FVpa3O8X6ex8ZyrGROuO
TiVjfgtH52JCKrHkP4cEmh2oQE2Sx+XcyTkpjQssvQhOoJRd5CnPfPK1q6Sl8ppf
oVs7/JM3Tm+sHtGiHJV7Y3y4ZB4IMSLj2wBXCbFA9Uwunn9WfWu9NrtcJcYiLpJq
2mhCCIDpI2wrQFqmSv+sftlr2sZAVfaqobhJfq+8A0bfy8UEXdUfK+tGtK3TG/nR
Zx1iNRWj/o7FzeGFLUMxJ1+tOetc3qsDUtVY+2zvaLAUzSTyZWwvSH8IW4AuUvrU
j73rXKBX7ho5+N37k4U5crxNAU0ScTP9WFqd9OgJxlpk9QI4LhTTERizMR+gedoe
hu/vIDx5uJ0Q2z5niKHM8EjkwiorV6KmKvyXWJ26pVBcZdMPNfjf+WsWjFiwemRF
vFmoCnISiDpkUtmnYnZJMFHJ75ZEbmsFgeKwSJgXt+Ir1kMVUe+9XOFRNG1meq6K
cc36s+JAnxgLSGs3b/bhDcJ1qQpBfRvQcoiOjdDrIHk/Q40HiNitpYVwP23vGsVy
lTwRtqkzv2jLdfr+u8/CbpdVI1AXOCK1s/SIXy0ZFV3Q0OVgTts+QBFheXdc/pxX
zHPFHW9rXTkceY81fq7im6NHc4AjrOJ5dI5wq86/s7VbUlOWbuvCQPcWqZofyLxA
MWzEzhgYVYJ/ejwbERhZst4nrUke7fkWI2QNO/i3KFgVBvvp7pUWFcLB7UriZBKL
JIRrBCLDP1up01FK+MxTaeecSMvTjr2Att70oK1DyQ3l02D4vnF++QCtSA8td0iX
Kf3XBOA6Bn+k2JdVhuteWbyPXK5kereJQLPe8ldVTL1mZdPSJxS1fELLyxU5+fQu
iJEdO7bPtd/bRq/wvKt9r0kxdWPPFUAXnP/kfEqdo7RGKMdgS/ivFzjc0kuhei6z
NcHw0Fu4mrsFVEYS28Eq5wdBOZ0MG38hSDnzXr6LUxbqEaW8zBPSjpdsxCL+GDhG
G3F7YaVhSvMgvm+BPRHNgJvgOeLlPbQxn2muYCt4qgggHObYnLBJqmTi58H+M4rr
oM7/Q8sDWF+Qupc175TOs9zO7pZwZz2xcwq3nm2BGXm8l3ws6Oqf2T4JlYCjvgBy
Wo6o82/KHf4/uzb7v/vWwGhmCm8zM92V9YRXK3QhGz9Lig4NI1ujNlfT4eHlh6Yq
QxiWPIFP+KsdrXv0GxbvYSiKNYkkEe9I6yVY8tVWza7FBxcNl9sinBhuBTSUCa1G
wBrLPkZ7SQNg8FBVll1ZOpqp4387s8wPgDBi7n6g0dJRlY5blOD/oRyvBlgr/M/x
nDMRTeMYxZa7xCoyoxgDXQpSWXV94Jn3aPdzSdhcBxI0oIj/qdS8NwTDi2i5FCBz
1HZEZaD8Bgy6da0ehq2LbdcmFFutNeEYePzDz2WFFkZhhu+j2b3yvFAjohvIjtGI
GVicZlBs6cW0Om2NiqFCFn7Ww7FBQ+1iAlXYH4fIF3B1j9wIFYoDjTaf3WcqlFmG
vyoBS/tRT4hDY7KBBbY5ajd0s+r6gRhFSMcI6g1YqilLaBppNs5Smv25FBsXx1nu
baniIJMMOPVbiQhxApdnA2ygfJiqxo3nU7/9hVrxa34P636Gq2OyodCsvYbmrOmu
RDaqp60Gg1ROJ0JaRQeEstHSTpL1p6FQz1QnplC1ir38xBfLMrFW52JVZWWl5Bp4
EjoPDXIBhgrWNbT/yvahh/5UQS4E+x5TIw/iD3PE6lvcfw2pkC0DUGe1X331fInX
q2ru0jll7HWSmdTuMnTbZokDUMqdxJ0tGEXJVeA1X/3awDoZhChrMfEy3qYRUxEY
o4B8ogUSdYvrysEZ86xTGyyr25S2eggPYxEAXRyI/LHXBZJppAxfdY0kfQ1Za+Jq
vw6opZEHsoojpqqIJKkCXAkWVBBoQOCms6C/biSOGK28bHhtCTXXvacLvFY/dpG3
na2+lCd9QfcaKC02TQFWu5kRQGaM5myY+L9QIyo3+Pbqj3lMSrQbI0qOi0vB5/UJ
5A4rjMwjbenm5GqA99ORnFtTyRsHvoy71jGavcvKKD3kwjBRfqALTxjv2WLOo/9C
8jTA7QtCyo5oo8HjX73VX8TJsexesjyNBqElhyQnHeoct00KXwQM/ToG/WshW9nh
8nW6BAK4z0qsQnbMXi/6fwXDFhKMni2Hb9OSVLJOSNOVl/HNs5wPv8aFf9XsvHel
znUHVa7jncHk7rQWvZ0TQ2VEFZ7mXxyL5NgD0aeBysNKMZBTbXZsvr+uEFbJcRpI
Ws7glEYnbZUxhDaSono9cOdhpKrf95xscwV8BzKxFbAqcMubTPsqLqApt1lfNyFC
+dVmunIlm6ga4QJRu2xU0ikk7i9Y+NtzzP1u1EWXp/U8Pcobyylu4v0AN2LXIsww
7REsI9lIVUM7A19aqiP7bHVZc4a3PU9VfGaV2QvWmW141WcHvr4AO/RC8MCxam5W
999ShYj7i79kQl74iPmgkKsUExbvnBRAqja4jCoaIzBrr362QDsKbQETAHo7gV89
bNXUYh2R6+Ug21TMemoSKmLx1DNtri1MU6wCSlfLWRqy0LfgtxowqvNlAAnFes9z
aU9FuaMK+/yurV3QjVwaRlpHU0d6nb/Vrrn9BrRvUXZklUSDeE7MJ4OV1HkCzqDT
7IduuEa1FUtSa9mLXxNLkjouIkBfJ2cFPnjkZ2NGcHWUEeJMctLnjW5U6PofmfET
e5Ea2bq18SQ4y7XhPyb8710X38hVQq/ax0yY6gj01hT7kle9SpzG551VOKGkrWIo
vBIGgFzGFqH+PmW7PWVo/GfhgTq3TZFM2IMYE9DYcE3EM5ZKNe9fb3S784MEa5Rt
gNokuh81xWrgj6LUqo0/nNSBFTp1Piy0NVF1dl7IcY5x/p6eybZ+SeEDwxiV4iiD
LsFqQNYbrdCkZxUu8N0X9NBGrZpjc3/YrDzm4y3O+hSvC5/8UE78RyPNq4tMh/Bi
xfY1wJMJL1VVh/qUbQWFIlA7M/gSNsF/QVQVTX/F+mK9Tthi/HKHk8QjdOtPYfGN
vZqzgmAVEBWvIbvyIoDlYp0pUaHwNFTXN2DEEi2Z20HVADYkD34G5T2UC4Md5CF1
AZCWicC/nHURuD/Ailz80vu1l1JzMcjE+SgyFgNqqsb9PeCyGVKDG1JnJRBRyQzA
pidBmiX/twyrceXRVtyF1faf6VROtZHDl4+eJM/MacD5UTQQHUjxQSxZmU/1wInF
KCYfpEgct7NAJNStOPLWjvoncQWtVj/kZUjreAInU69WVTJsFAS8PeKtkgdNhmWl
u1FQpF7FDjvGvu8laNgjsJBXH0i00AZh3R2TUQeylqsR8J9tV+lQPrDrtnjlBrVW
KMQ0bwGHFZlb0mwrItYTsfFzhga9bLnIDhydPnN9eRLS1ivA/9lpT3a/WXgqCTNZ
H2g5jcF0kHgEjxRcI9NtFYbk9zjd3+C6yixG/gLWNRrJsSfQmmbhUS4siS5jokxq
x83ZUXNWL/o3pqLbv61ehqxwegiPPthSCXoR+t2szESJHyZwRRPL6zJ6E2xcQoN+
gxa0x6bz5dskhuW5dXKWrJdSM/bhP928qStJ0wSLisL/YH2kBWh6TBiprZ/v2/Fj
2ngTat1SSnuO6D3MEgLphlUvA6ie7Bzubu355QELdOCXGnCMJuRFxnIcJ+qyGD52
fSE0dSYAQVURhH8nBj2bOTBz9dJc8ardEqYiJ8Pa6mijpY1b+QRiEnX8Mh+enf4k
0dptU9GFwUXr6bZzw+KWb6dzMNQ88ls1jVtKXZMfB/A+iwsInZxFvxdBXYVZGIkl
BVK2e4kpyaoPGkRRYTa6rZyO14cErE+pjPfrkNNPBBcjSh+UfPCVJqE0uXNrQL+V
nZcuWb24XGoKyy8ZI5lL4jxe3JSigGjc9kGwa/5Wt5F6sPJ5gvZmOvqN/V3VNitA
d/FDsKI7hJPGtUEpC6R6wkbZpB98WZ7dFKvvGsxtTTgl8Sk7YxpqMRJdycL70wyY
xNVLa7t+DpuXyY2wnkMnYMTXxrJcj+w37uJI3bInDh1g9Z4U8C3BsuyNdX5m2YJI
s9VnpmJvquPIw4fl5OiY5TiZxCOWiQcZVeX5Ib89npDMmckO1DzxGMmpVu+n5gQu
+8IqKh3anOO7BNiAa9o7pDJY1PEPtReIvV88PeARXeg433V+DPs63xivhKf0U/Zf
2iogX/OzLqPaSy9+cTpaJrmzC/ggN3LfLm4xXRYrPu2ndEMiCYJ+m/dxpeIR/3+M
HSWdTkkiGq8RHoXsCa3WmnAwh8VpdfxvX0ZYh9qQyBQoxk6VyuNGFpe1xRMLO6Wa
/qyTJKzeJRL/FRn/QDfmVp64hUPpr1vDM5z8ibLCyNVTjAPuWyBsTGCuHO/Lz+3J
lFGBHr0H17uN1OoH3TifaSBVlBLL0+zvGKbBpCtA1BaOcaaTqUNf7iPFXYciKSep
U56ofXwaG7EYsepcmg35kpHXCZQ7hy7iY6XWoBDN8TDUTsv6QgB9VNLubZKXTp2/
qezpeTb6Dh9hdsoq4r1NkdYA/z82K3CHo/v724yMboc+wCluuQ7HTzH3V2BJwgeh
m0wYAEu+f+ymYcI/zltC/LRTHZCPcC5CKGv+n/2Y5ZoErTLb22xavD5cz1H7Xv3H
UdudyNAtLvdUecC/L+z/JNr/90OiUk1wqg3IOalu9+6fidby2uu34GB2fDS4Gf81
2oi0G4v/CSt/NIl+Na2hOwM/se4LqYYsG4OSTRe4syCJNQ7TmWsgBCTDJY5UPvK1
7T4Tsq0sMD3Q+HNmL8bEstZBYAJHEamhyj2XbtRo6phj1qPSwMzLjHcY+I6306YG
O/hRnn2jnAQaHBcwu7PiQSftuyqx570yPGocEmnLVd4XT+pyRgtPNL+grN2108Cy
NmbDphPINZZjDs9XzCtc2PPtr+tZXe91GUJfNbLqUWLBfNyKZbeigZ4amDQohz/F
TjZYpPwBSCaCbaXeoRQUk14X2RunHDPDNdCGXMOnCzaTHgqpAwZp4f9vVf33IU/e
rIwn0A9UyeiWQOUSNds5TOUbx/Qc7Q7NjJ1tYTerPihydLkLG6r9l7uvBevMjiXl
mMZCPdyuhiT821/7LFfuk8BVbqh49Q7MLJ4JAeJBrSHvZpcPOnsuDzT0R1RPFywI
KY14ucl8odWhKuG4ua8AWgRb0pEa8OLeDPkaK1CWxTO56IxHd5ESpEH2irfNWv+M
+OfVCTRf8tdNPNWjRcmWarKm9gsa7dASuzl2F5ONJpLReD9sbXucXW5PwKSParcd
wcGSp6rS5UIFmMAyppTX/WxHaL3Gp93xIBjc3OWfHcKa26Ukir4icLlIZga+Nd4j
Hl58X24yu2T+Q9vON40TIr56Mv55/36faZ2j0RV8hgV19AAsrEUrkqvetpwKkUT/
Aw3cW7ZUGtvqc3DaIpjkh5Oz3hqGWwLnYZnd6ehXEfAsPKkAxoawg/RK1c1YYQYe
85Qazzwpu9PbQZhlin5NuHhuaHkZjwYD44l0QX4YJDIUJ1Wu0HHFzBBuOWOQE3Jm
mV6V2CZ3S7FPDAkx3psVFUkYL1oJKYjCHoSkh4rbw78pxtzTsxNTfOoHCKtzo8ch
nD1y9zEjK3NWwBYyKqItz+0FPmykw1i9UAgdNC/YF8XHGKGGGgdzVDT2QMJ2ZNLl
B/S76q7dAnALzX+KVoSkRjZws9xcBn41Ds/Cb5VWqfg4CYPUCrTLO6vgmTXJ5eBQ
Pit78YpgVFQZs5z7gRPpMDpY2JxgWuy4gRZTrZH/xIvuo4AwZT5gynbvl5/ILig2
NxsBqBQe+IuO6l9q35dyoRwP8FguKcYly5Kh/dBXZKD+B4ieF6sbPD9j2xds4jCu
BSwXe6sJKhsVuV5Sm3JFjlGmvZMSthNn79u+1NQ/LN88igWj+xVX+E32FrxUl2fI
6q/Pz6gD8nw0TuuUwNAQXXJSKa/Ol1XG2eed/AoAXgoA1n65LOs9YU/Eq/KN5hUV
B5k58K/olWLgKchYvrEmUKWRVoLDdWstAXvnE38A9YTgfjNniHsfdDHbHIWDRbV6
e11FdPnQDMx5Xx8gawPsbOgg4C/R6sYwDbpfvbQpGCKAwJ7MkxBCoSRyu8UDD3SH
Nj3WmBwP+wIug4Y3OrWdAx4LWSV/bT4ULGFCkkD0rrOlh+Ta3gDUngmRRA/KMFQq
6bC6bAF/NEx6LInySDso9I7FfKu90vvmUFhYWnVyRHp5/s/tP35UKaLZ5aSuB13G
Ucu4i0zddyPIEwzlE3Rfxv5f/LbAJfY49mukqftA3TF9J2XSkTZzB3XyskQrgTiU
3IEh4/BD+cg8PN3hEQ4lKxBzfM+FWr3S8oKQBiElR+LFawcOW3VPLZ22Xx5lYipM
sTDXnCn9esdJw8aGaFy7I54YrFunI9TMSaX8Fz0F4WlAeAWoRBZmnVwL418c1alr
QqokfKT426EGOJL3JlSVqibTpMHSEO7fWqHOOF7fzNzmeQZAtVm378uqKPCQ7Sji
JH/q8Gq60YVp8e0Qjk8adhSaVCpOat8QutadphY3IjYEQTDrLZ804z94LgbueacK
z29sQtTYRP4QArnwxYBKtJniejp1b31z5/L/opzM8mavKBXUI2Y9AeBqCPVSA9zq
lzm0IqoMqMn0f316aWQZH+49CzUam/5nLwJyu55A53vdWOJ1Xq13En+6y6KuZEdR
2T5Q5P5UVekNpMBi5pQJXLiCVL4oEVBAYnMwCM/AYZtXEld5ff2XmH2lei2hnU1l
192du2G6K/EaNAvObeMts24jZbLSzmLINbAcV9tvu2rueAbjUXxerju1mm+T4j0E
u9IN5lnXBWpUkB1ejfUytEhwZ9n40KfISuNtW5XAuUFrENFXWZ6CVAtPK4WsjaKA
xXrf20v9AGmnXV3Yf7U7MW34rxdXErCmDlcelyKCHWi/Fy6Ws6iffFeKJjRkJG1o
KjK7ReDqlzFyjOg9bThrNhGFmFk9Vw6fH+P0AdJCuALdvEcnj4HD04oiHuzHU0Vt
4sjY/8Ug+pMoAGBjjwxUgGPSaUhaZ+TqRrmclaJ5Rb0BTIMaMdJu9u8/XzFfvM9U
YPO+bGo6ppVGR6aCvKB9e3NdpqGIO4EcoK7d7F7dITZF2XaoPAzJz9f0SobZrJym
xi0ZSgn7xcHLdHaY7j+obOHkTPVSVY4/otaA+lGYpRxbgJNa/IFzUhBUV3cBU200
brHZQFgqsiPP3ZKn/2OMlWzJfBeisMZaeFCEdoMK4N8++URX7iWfwIGe7S2wvEzx
rKWpplIyfh8fk3rCouTGLRjS4gQ58riH0Fk0a6sczlNtyc8kFaJnGytW1ahEjjBU
Yw6mXK3yaurOPpLbcJ6BFh092XrjGoR3unQAkwq76pp0Iv1Syk04w3MfaKMSFNm2
5fvVGIc6BK1st1sYyDPkJuJcXykFu8sTyRyVYz9rEo3bHOdu2xZM3xTHE26v+woI
hh5sQU94HyAYXOXb17o64Ubn48qhn34GOXqBgjvdoQfGQ4NZ90XSadAKrbRfkTaf
htrBbjsyqQKxB0XB1g1yRJf9Q2ZNneLsl7tcsX6fkgfRqsk+fEfIvcsL7azMJl+8
9xEsecEtjO18VwVKMD5WqPouCy4R0Rtli81PM1OmwOQ14mY5iRgqQxePWDS0metp
s9/0FOsZjurbfzrsNk4Oaqa9dX5WgrTD0TF1F5VmFMt0wp9wutHBqSnToyTty/qU
rQ5V7M4P4cLgXaKzg9wCu9vv5C7St1WA9ra2sbzB1c+WqK72gxRwGyLp4HM6wfHI
M+CWe/YkCyTDyjKW8oChDokqYFRSgU3fcqvJMDO/5LAfnXxshWHpa0uuyJFGx77Q
fZOgbUSrK7tFpWKeeEhi1eg0muBMc53FQwDAiG2CLv7Y6BsCZCUtrN7VoKrvPS1J
pc91zy6fZd/wthJVWAv9lfDUdDiEgBly+nsdewWtL0OtSDNcSh+9BCeZSUaQlOI7
PqoryVRqZgNVNDFLjapzZqn/89+Cd91AFydVYVOQjt4MJXTbjqEvsz9R1wf1ly1G
CWt7HofixmAsNuArU9lG67WUY8CK7lRYGK3vCa9rXnxC7QIARE4s8IlCkm8eRECR
1NiZpYqGSASzC2eDV9amkFWmHIcp0rByaR+2MMSjAE9zcNxtq8Guc/sNoLC9rJfr
t0Y/kXVWdDHuO2J2UcL9YP0J8MVBYHH9yDzyjvFc8yx3bX6jF+rFkH/vzppPIrNp
7LcuyRzunkogPWkyoQJ6SE3oQaKJU6WNNJO9HWMrlYC4VC34+rH5wxRxZp7uOAGd
k5/irJerX9upxVYTMJjlhpcjvWmMDIWfuG+Myhrd8lRxsF1b4uyWbzYR0rK4Ny/9
630aqiLnSfE+KxftLTQuPjPpjZtquhKw1ot48DWZNx5QNVyTSAZD9wm0QTFKs3u6
uulJAuV9Wa5b9j/HYkiNGnI1s+57Lz0r2Q15RrO4XpuWc8WR//B4V9Jh6zwvqcyF
qZ/So9Xp1I5oEpC+wmxr6ELzXRVWF3o8CEHRni1tVjNHdHyMk5Dn0yNfep7FCb18
nmgd2PHPZI42IMahJUHzO5xcQhkxMI8jBAsUNhj+pcoBr3cCAqBi/8l4IHE3Ig+v
yod5fuCzQCxSG4gxy5geKIWkpMV7EwA99jughNf0BosjotEuVxaK6RbNtQWA4C0p
iO3HIInielwT/eQrk/w774+cbpRKbxXzhaJTaqQsqIRcDuhziYjDSP3DUlfhb0Tq
OII15SbIwixkch99nq0pArlYjnDrasrUHtuHn1p9H6kBTzaRRDxHrBjEzyu+zV5H
NndwlCc0bfj7SsC2xlQ/orB49V4hRGxHRzLRUynmIfvdEXwayELc7aa1I4hui3UX
ReorNUT1tDjN62Q9ihMw33nMGYrUsvsd3uOMlYA0ehG9NCHhl0JnLTHSO4f++pna
p4bZjzXyE5B0nN33PjLjOH45kCLGS4zBY5CTD6ImdtFkTE6WLJ4hXeYAUifNdDTF
CVj/hQhx715jJp8K+Fm3rvAJZwGcCBTVYOcJ4cDOx9KHhbx0PZffv3JjhsVh3SBe
km5TAEAmu28/RvKinRrbGV5BGUJmrbskflYUSaSRAF51HX1/SWOmm4y2dzESQToH
ZdOwEOLPsY65/f89YRg8voOhlY064aRuwS054O+IBMQG5DV6VRSeW01/v48H/C2H
QT8D943pcDgzNLteCJlr9U2OyE7whmJIsb+dWYyqqNQgiwsAHAt9SBCTdsEvHmLW
15wIAWRWmVouE+0MeyRqyZrsQJBNUDGn2k0aJIq2rbHTC/erAR4cqeeIyFP6xeUi
OveNQJdlYDvzFXov/MC/lNI268cpHvIxqCl4wF87uzuL6Gz1WlHHVokr6EeEqDhb
1a0deotSsrSOvBDNCKykDGPqFYfO7yedNrM+uDXYgIxmj5SaieHYqBBE7y6PQiRl
WYpQhVLCNm7TfvDbaJy56LPQi+qUvG9x1zUpWedz6iirqjFEKvxVMqs/71BPNhBQ
IAcg5XVKvsOj7RJ2CdpMGbOOp5aP1T07A1lcMTR30O87NQKqr7BS2zOZ69jSMIby
Ihyy92mmzrV40kkD6EPDXTpCTqV2o3WQOsbFIWYcCMnsT0LjUw5YPuch2Dwgx42w
ox0rvRBfTJBKhqUS1Z0xUEKYLA3oUQsGZci7VomOSbS5y6iNgcwbJlKlXBfW3ltY
b0tyd0QXwmG/uAB8tkJ0htfQPT4XC24Z6XqxEdmeNY99l17KF6AFqnEioE7xbzd7
9HV3yio6kl/WvEuSpo7h6oEn2prnWD/0kwadB79vZCLCRg9FIbrSPq1w4JaGq3C7
NMR1UGU5DNJQ7MJXZmhGbpWxRtpmgdXjeG1uL06F8mWAkfG1a813nTnEIkV2CUa3
1qjSS5m+zU7TQJlzGH0bCWSqTBRXufyY++8VxtmF9d+ZmlLJxTqrlXSTKSb9oMMC
UwPHfz/51pMDGbZf8WcVaLSYIW8iLoqZPaIAEWruhg1vNCv8+nscXwQCHDDaizl7
c4aGEdJcRbKGm0TbPy88iLU75ooIsLpFGTg1wra9BYR6hF1m2Msz5/am0OSwBsqa
O2yJuo9PDELtySAux7GRc57qvHIdMH2p8fJFwzVowRYMPS6dcWYmQGS/WEpgPpj5
VNAwIdgh8YRnkt8GUpwTDx0Ha8qGkhuKSXyk1gyTyjSI6FxQ5Ap4oVoLs/CKY7tJ
URlnNNKdI5CavlBOACH3WPeDykxMKBNI7rvmqbxJcyGi3YVu5UrJPNpuK+Kdnisg
t8G7bVZ6k35nvOenHasr++est5kPlfo/eWnrJZMK7pDd8h3Alt+22nhutCQmDDeM
qBpmHVoqqmEDERb3tD4axLidFTNUVE/9QFjEvULE31clwqjP88ZY+TOpVkhNoku6
v9C+eKSWg3OzVyauAbfOcJiKYZOtXluUxnVUFGPbaR7XcMB60uMnDe/jbekOMB0B
qz8RkMoRW1dy3WbnpiVlbbqTt20MilGlWc+F9MPYyjZLde1W8GpkGud6b+4qumNi
YmDkrssboU8uBsNIo4+lbEdI2Zfkmv53pEZckdaSF0kJxbatt7+6TIySH+WrSplX
6BIZyZWTMwbaZkBfsa/LRq9KiNwyYe84ok+2crhN3ETaxFzRthAk35CIaC+r0TSa
pAYFvE/uVUN6HnxeeS7hTcxGOkjaajkncjLD3gfpaOQdfDrZTBfTVw17fNPdNpie
mGwZL1MniVh+6q7UllJiKrpeWQzdMbqEUChNMJYpn8a+cM4Q9QZlFzzAAXJ9Jbvh
O5xblQJRPbvorpypxe60DBn3hiSS9M0UONOBx1PAqSwDl80+Z+YAxrkO64dOvW+H
PG/Dm12h6+fov/5MmswfXt9URE8Z5iXOtiVcYcicFGS6A/VNfo8RlqIhrW5o3wUf
792op1OEYzQWu6lRrHV1NpuYgAfuyXyqKT7f084OKYsIGSHbKSdLJi96JM3+EbIO
op/s3ytZeuVO81F44tNrj2ofUDU0AIUDPjYQVhFgSxaT/hEKnJ2M5pWdWUxt+1Ux
HeO19Qa3wFV+4Hyi7Ka9DmRPdb0BdIp9iCwYhUW2FffvuWL/08fAgDPuAjn/01y5
fkpnKAu6+KleCGHMV6QePwuLgx+T3ivpPMpD4XT6YF7haHTrYKZGkwPeDAojtvTx
ghM/JChfzx1rwzO2zC9vfVNx1IitzbCwrNYUc0prdf7m9bYe5T8sp0Icbc6j3YHF
hVqivrUC1Ryby3ZrVaJjc3cgtYYwj/mk9451zSLl5BYX50AOINM3/XFXNQppPt5r
Sc7qO7KnYK9bAVngETuIiHtJuf0cFzvQazfK8YOjb63pAbhnLiW0AHazKaceq25j
sUifuXXBJIhVzscDfW6lvOw0/A/7XghluUtEhc2GOthRrWRQ0sduSWGMZP/5ph/8
OIn8Bb0/EBeBx1GKWVnl1wDs3FZ7a4a4q+XVGqzQAJhZiGVm5Mrbe86B19D6lzSX
L0ZwtaS0nt+9XZ5a79qQVR9mpd64T1uuzsdpwsHEIrUjGbNzRZOIiTSOwCKYbYHL
svTcuF3b8Nqr4Jt9y9AjcHM8kiegtt8dCK6Z6x9Ha/JjRgbeoDwR8F5+vtFMXmJS
U7ep4jD4eK5/D2oPZpXWMVhlfohITvh9LI6aE2E/hUhgQ3hj95gKirS3bS9CIZRl
a0mCgbNcARPklX4SI0KS5h2q4gd34yWy0Kp8iINKqopvGuuivMpFe/oNaN41TGp5
nbcLsokPEI352wQQMvqhE5nuShlPqdAFx89UMsTDn/mZI1fq2LDIHsaUqcy1JATv
1WcgYKTiojW3luDUahJrM03kX2Lao/EKmEPck+y8bfK8vD9lRfXA+xYNlxSdPa9l
wyXvW11wQ/eX/G4bxq/9ct9TitwZh99v8aZBLWOmb6ImQ3tuIxSj/+H++wAKTt5+
YEDHCglp21VePkfFGRftvnABHx17j0GxBeBiu/PNmRSt7lNkTVtU06UHT7ka1nue
AEDNdbVGn9DWg5QzxZ0q+e61qv0xaSvde7li9zqAPFdKZaCxpotfyMLlpBZ/kP+S
LF2tKqawRxG4iVGlk+F17ip1vmxZLXuDc6A/tnklg94OKfB4khXSq6YdpqoPUn5Q
eHM2rty8OTgPKd3+cNKgCjVFRQiOaeS6EU2cdjo1r/Le5D9yW+Zjvgk/joTl9pwI
t3HZUQIYFoh7YjZRLeiJsJ6i0IjQ/2hjRO2s+hBar89BdeDd/Wg1ouhF5sKwt0Mh
jA1tEduBAzH+OhTAXBVsl+/9QveuvPErMlZE/8M8Wiyydtj8TCtmge/NhHm3D+81
5y4qiQo+54BiXyE8mk9xth2ynwKGXLw66FgYbPOY39oPfeHlUfNsSflwzyS4MXir
U6Cfrq4ShGtBKcK52ldS2a/O7UQMLwJxi2dHGowLh4aHG4VcAvi3u5PrauK44TJA
DjKss6UEyk/gnyytLvUNHcdYwg1e349KS6orvsNtW/sjG8DGhXwDkZiLMgd+/hLw
t9uWCZGcAdevslbIt2Evk7EUzNEHReJQ7cdrdjJrxhHDJkHFLkOp9HlndB4W1A3j
NdS26+WcDScqXOVCHMZHIq02yIU0Pz0LRnSD7qCXNLEqvdEyMGewTl72r/pOFcdq
8u4pvDZt4y+5+h17Sz0fMdEW6LeIANOaJw/1na2cNVvPtRIBzvCUFgV6AeODICSV
fbBCfF5qArhwcO2zWYgZet3qBL2MxpjzKEU1+Ym/8Z8grjdwZsN81edECU204Zbr
ji3R0A3toKqZBcczzBe/zBDVAvR25ngZwR9yl2V79jrb6Q/9DtmOs3XsoMLDBfYR
/87q1QIj/UhdDNk9lRzv21U/hLLjjLxrmsrrasEhmLP1uQDh++8xJvE3oPBrkFXL
EtbUVDedKopUNyYIRMnL80uPCPX0EUWojUmf4tlDtvtf+QB/+OJAS6YSC3pR2WQd
Hj1gZjCH0M6U616vRj9Vhfgvs+xgy/pFl3mgm7DcvsTOdHszt8Civz5a7EOkhJIR
gxxNSPPrVl9qpq4lFlPpiD1Bsc5YNTC9kNWyofj9Kb9ZCHh8dY4SXncIo8p61E7F
xs1cosd8iJcvsgKoFOmWi/z4NeIO8E7LkUnwhQtZ6YxWmjFG/vkwHILmv0YPWF1Q
mnrl/yFRHLgw3lQbKZylO7R9CeK+6EXPxnxq/AeNXtm35rXJV4iAVw3KuIOWfOkE
QoRQMtAUrPIoc4NWrM5uidzj4v/qj/x/ZuuCwQxXsO3xAs/kQvIqm74xyYp8/HUQ
JIZWs0bAkAkf2TDmxyLBYvxLoCquEXOunS4yGUfEnjj6kHuss1WDidPrKoywS+GP
9wVnmai6Y1GOTF6V4qjrYiHI87MIOnXnCdiqoWMNGtlzfOlChyoKk09c1TCFqPIE
gWh6J7DDYJa1/mycBNLJgrFYF1zuC6n+7Vq7nXGoYokh6IPzBJv3jAaSjoDAbrD2
GcAxch8K4p1AC6nGMyTEOSpGwxPQeQFKluWhurPajAz15apQG2Yw5yZNAUR8EfDD
Qgccvu1FgDOncAlS6/+wT6Qbt4cvLwakQ1A1edKTv+A1WQsmFfd8fzwr/3XUut6l
vACfVB5h8ebPFFySOmDenAGqelaz1gic5Vv35xAAM9hyTvPVPrw/lw8ysmixH3n+
b/eiNOXj1vcGkY8FLT17KchrE4DpSJnmUetnNndOsqDYtZQPJzzTFZ2A6UBsou5S
u+r2NDqFF3Ar/Z3Usas/8B3c0XochnFQI0i8Q7+1f6VGWWabu9692uWw4eEv8jc7
ii9T1+06As0snynCzBqUi+K1zh1IM1DX1ZmKWrysYu5pdDj3oe5u7wXtM2wD0e5I
4g6rLy8Cq9F1VhFvK0BEm0bezMl2c+CZNUq24FL9EFq8jvgGtbiZm4XpR2avDaOG
vUSHHRHCTWyB3s7smPyR82tYd6myY++VwW7SllOMsxQ6L7r/LD+OweVmeIs9vLrr
w5rdRWtNCR00y3vw+97qorRgbJ4kJAt88YPxhmk7wJspiZ6TNrqmT32ckJBDMQl9
3eEhp933Ee/Xf2NR5LhjyFGhK95Le977pndzpmm0UMG8tKkQzq6qHOTDOukMUL0u
SGUiqSMKvXZIvuBwZlk3xmDecSr+qr7e5T72/iI8HUb4qv++0DHiDEnmjGH0n/4G
gAtw4dIj6zlORkDmpl9DMwIAYItbhyowGhclfwoyGuGmPOtmbu/bzHT2ffU2ACYu
RNPHXnT24rrij2t5EbVpwG2zgvnVTxCUXiBOQt5F/RqCLJ9HI2PnCL8P+UVyQvCu
R4Lsgf2TfzN6RSf/bPwzF3tGPpSFM8Y0iCTWLKVKdV2n/jzAVSZ0DqzHYKfdWS7w
G5S4HNrlStgu2yzvLzTxatq/RYA5CNbDGXrMhzpYhRAletGUEX6yNvTqoMPd7sXC
RkHlTGY+0NUAKEis6wh6Y8iITkUznPeHvgyS0KbX5da0+AnXzKeBC8KesRKKbD5T
xXFvjldSP+68Xt6id0tvHWnxdINAjlg9nv8dGfy+sCcfbyFaJRmLBcvTy3mN2iK8
xN4s+6wNxYEn3YYP00u4w16qtxgB2RvWJzwJXhE57iFSGNY4038zy2mwTexcQDC5
nY32zYsyQyR9wG5glw7gfeY03skFAM1V9av60SPZW091It+ayFp39lVo0NMTtHQE
UFE8xirSGmterxJPmnylTwIEramTHdIQgrfalczeyFmhBIvQXawy7C9tscQa+ml0
2n1UVZGyXs8aMdKS/GCbUUkndMPcSUwreBUQN5cY9i4138CC6aFPAsCGU4CrvKfb
9lNNLy5iPVBug4CQvlWGmzArqLsiacn1KcbCkpWIF2vzd0+Zk9xkLdg10sI7yrxM
TANNV8ZjIOOAHCLN3G4JMJPuulbsxslKeEkwQSDp1VSGaVffwKYmdPL+BIFvyfHr
Ijq8dm4FnC97G8nEhy/zTPa3a1rG9f+GnBsz9FHLsxPldm0X5V45bqvxv8hVbhS5
SoaHWnexIoN81ySslfDY5lV5tQbRYIgrZo5KZDg6SRbXo+7jiPK0/rPOtSt/2QEQ
XXrck2vgo/eg3/U2CJhWSKvpIAN1dV5hQRYRSV1AmIFiihPTq8tclo2HkOuGol5k
60VjDT12UoWS4Co/FCGKNmZGBH4Xnx1swGhdIWy5YzHNs2e9a/4odk02V0KsGvq9
6+FC2ZUGBR1dNYz1338JOk1dHWufkeqMdX445tTvt1mTFstzF+LreZo5Brz6ndy4
9cwHtIthYiQcFr0pkyuiS9QcKRB9O12s/i+jWEBGoKBTZAdEzw8bx4ooz0NjSJDb
NPwENP5hSeQgdyBHAQtP5dQTzmSSVYB8l42ek7dvLtazTJJKX3rbtds6Yp5rUbnB
anMORHVTG34jOjd9cmJeCGZV11ZE4z6xi+nsUDrZfF0BODWxhT9n+cb3FVsx5OT4
iTTWef8GpVjj6oZjoQrjL5mmUY0dCQ88k2V379btx+ZitFvbYF5+UT29M1//iVvI
L89X1BH7UOz4FekSBxWRxqZE7aABni1z3T2TxjWJ4FgvmgsqL+KB9r00d7HhOxlz
BU6NkOrfu+ncUGKM/9uznM/Fa/8GMYDlkMNvsvV+fk85uX9iV9/azH51UtTEHhQs
LNyw5Npp2gKXOp4cWK9nQNNjPYjVV5y2R3nASdCIob7Kk3rFKXMyp29Sz0zXil3j
t/oHzXqgskiDef/zfUvVc54IWukZCqfS+Ilum/ZhpqH2UA7pIE2eGT5hg1BkXb6w
fZJglPTsvGKU/Vn+x7ifN78C27uzrCdYl5Cu6p9vPn6OmBSruQFoFFw2wc4SQa9D
RbV9UafOuffpsY1T4jH8rbEHpGWe6Sy7/QjYTSem7HLGtj/d2rCoWurraYRSCPd5
FzXp00Abf76hTDaBztairYGVsTZOhtcmHAq1fnYJeBmo8AMrgWtOsdUaOYc+z6Oc
3sSCWY3qz7A/AdnM3byCxDYa1OKtiESM9kn/dTYVvyNq9MzDb+ygY6Qqgr2Fe2sE
JAiaa5N9Z/j9hnnbXjDZUILq0665IuO7rARvb3oxEklhv3MetL+phX2BLexKORPA
oe5Ai1NsPTuHOLvgnt8vY5FdYyjrPLu/i4/XiSSQiBMyVkmy1IFx0ob8ncxvpKzg
h1a5tkXxVdu6Wgtj0z+b2udLm1JAYb0NgWUtleLrWzZkJzDDPyINwZGdZ0ADi/zP
rgkCRyEF+bR4kWng8YwDPPTuFtkehPkXxPjtymH8Fu/9SHFe4yI7W8ahdLrvtNhu
mnlyiaQB1pwYauxlxo+1b5vJDwWF3FzBFWWETNyETy80PPTs7MGojqtZZvJju432
DCKBkWl90YzlEs/1ZQsXBQ3Um6DiHZW2FWY6nMkFdQZrXcek39+xUwr+iuVKCDys
Pq1sqMQFs2ye0Bt5NNgKJqwhr948D+MBzua91lVt6/ugNTaBfe6/R98IS2KPzofj
9bTowahaFIKZi8BhmkgMrtG0OVveAMz1vwdrmRcq4R/x0ZB9IHu4Q3AFug/N7rb+
/vxnKXOTSB5Uhd1mNEt8gs9H+YUZiuaGXCfNFzbW4h49qSAx9AUTSUJobJsbk8n0
58ZG+9uxz/IU+6Vxi74shW8d/4diMAr7EfRVmhf3Qu29MZHHEDWualyJTXu9tCkg
YqbyJNcGXeAnVrqyEsySNgUjdpn7x/wM6bdEs4olEEhgHUrCY+trxJAYUt7ZsQZZ
3L6uPWTnla9Q7r3ooDlGph5iEkkT0sZb0NLYyhDTSuwc6CaGUSQLeS79SmsdI75u
q/r4iKjPjRe7/eaCN7yIPrPSv8tndxh1RqU8oATX1NCO3RPINcf09A29xy7jTyXi
fc/UNHtEXcF/Lpz7kkRjbLgnT1hrjMKO7awuDuWRVH0byssjz/zRUpwCVRsjw8sv
iJDplpkyqUaxlJo9pSSPqdluw+QmehX0S1qL4TUe3u71zupQCBXeVE2HYaiK2Bza
/UbywTDzGGS3ikyQ542TaTggCsXobCBbFrBPPmOktEAuN6Dzi9u+5/w1ZYms5arh
hSktt3T3iVnll3v+vCLeETQGBGGjno1/Mptss3PKSj4FaZs/b7i43/N5LTLmZZSz
bnaRF6fAo+8jyz9Tr/Tzm/mrDCTFx1W1YjybVgPaHs9PXNjDusMRJDaSorc6TKNB
AIuBm8HjrEYWA5vqvqiAwecF12kp1Gas4PMjjI2Ut4r7WJX/yovOwRoNJOCA3COI
RSjoTBwSOoHM2f12rZJ4aF0G/j4zu6G18/JueTfCeEXcmqAE9SFM2id11p5Fcrlu
YGNWi3mAv3df+TR95g91II94ssfV91CIwyNdftaQnvKWdI2GoGQTGZDKvt7+KAiV
XlNM9N7E04EtxDyaXiGkvngxEg3y0a7+6ce3Vit4WaF0x7aYYZMalITaeFLjFzHz
xV+9IDx/dS4IhcSrFoB2mrRJCz9SoHnWcq6FDz3E0rTIrjp6UeVbN7+EPHoqZ+rb
6gBOtIQM9r/D4yBKAJsNQKrfb7RaxxwNuoRPJJ9lDH+KWS2Idck005jgtppsLlTf
iW4Ap+iyNJjYH8rEZLLu1mslcehNbrKUua07VzZJ5MZ1cZg/wTuqiBzA6hyZM0s6
HnLF6l+/T9/6CyQDBUy/lL7GxGSm79nK1JHVWGrk8t9FVUYaF/t3wJ4I6JrjzqwF
deJx7if3sm+cD2ajJOm5kFhdHGLkJQUYIMJuSO4jBkQFS+ykylY4TFfoNqHL01MU
huHL3O059T0gsQjEfPK4MPTmzqHePuI9n/hiyIzI598F4NKKUAbyCxNzx9UZ4jGs
H0e2trh3K6AscO9AJ4XOEr4vCdSapwqRplRsh0wj8myg7PMud/G6M7UKhJKk8p/a
+03j5qmVzmnRMaNQcPxRLxjcb4Ibhi3vAji965D6/pTBS1ES2pAR+HqcuERTyb8S
kZwZiFMM15FzNwNLhLq6glQ4+YcB7fM0frKcCpFgHmKyXTXdDbbk5FPQgMIxj4Bv
8+QmoVfsBXhkODqcb33hL0Xg+zY71BsoPYCjCeZKtJuR2A+CuF5OMhNZcBIEAvC9
1ksnHvENQvEsR42pCRAghmcEoZcbxZFWxrs+LNkUkAdxI22Qb0htKGByqiJb8BQj
VESwjTqw/XXxv8z8BuUHrULJwquubSOjv1qls1qt9K06CfBHDKebC1HLxNB+NlPg
+nSa4ZTuf/WRhEj2kNR8pu7SDBTcSMJqLS9DkoDTaOBslykRYnmdfwscuLFSFNtA
GVxFL+H/YHreYVotfvj3g246OtbK7JXLtNsFr8Q9kyemXcdhYlBR4C6vAXdypVuI
4M0aj5iflRNhoI4ennMjDgDHPs0AVSWdgGMtNufovOmOm2LAtnplp8mIct5Lkg2g
F4Ol1VbjZbi5/dF4eU3rslcvhBWeYOcO6sLtSv4ls1DNT2ZC5XT+05dP0IZtZ8KK
fSRLH6iAwHxivOCXprTvbQ52OAPg8oHES1v5QVf0ZXEv9DzPs6UARVDi/+gPBLEO
xNFtfes0ao795K06CEIxW0fMGbCA9ckx0NPthfvMQZWIu9Qu80p0UxxCv847WIc2
aTh8IMm391A0OoNEolj6opS69nK9ZNJWLGpQfOlZ333/l6AblzsSXs0g8JVMXJDt
pxHNJlOrrdEkCYHA3sjCe56Jnj3D96WY1GsuO/T2Cpjc+vldQytEMNh774QoTLjJ
H4St/0UphkgtvdCnE3kC7X5O7xSAnImpBg3ngOwJBvl5Ce1kp7e/mJH5yWHIOttB
n4X7u+bm+A1GUIO8lpuvAO2t1gxS+XK8+UOiZUJK2UzUIa9l5IvHq6qyfu95SMj0
A+HoSBbOt2eMaiBsiaVCKXfWRS0eYPpomWYHkolAO0DqTnuRANsIqGD9VbLYbE/S
eWz0jSwdN+3KfLgnKT+SCh/vneQET78+yR+ZddbEbf+EqGks3FXjJGc+kYzF1dnY
lG7DJNfJQ+weGgBR4XT5ZF/6EAzVy+fANWUGoc6U5mvFbqfZI0gsOnAN0y+SWgCL
gVCxPH08H2FAGJnVU5aqRg22M8wjMdEaNTGx0ONJTETjJMgdY47Mvn6/sQyjlT10
qdVHn0MeWBsaN+g3TKhqYsVHtedHCkgQR1OJ2nFsDFG3m/kHjTK6vrpvN+uy7oCN
0yrFXa3Hs21E+xVd/Sm+zVDW/HY3IMADVIr3TlGqSm/q6/MNKE6plmONTJ0jqkoM
QDHvqLCmF0q+AQTCUcX9utTUGNua8hCGVHgg6xeCYfDyge2OEp7iUUw35WuCZCMO
/LWM2HVsTQi5JjOT5A458MjX+Gwk7J9hpOt9rkmIHBj1mQe1BY3GHwBXRCEcV7LI
qiNi9vnpQSkoS3K7fODyOOyEC7G/+66vGNJSkvQHMCK2lahYZdqB2Z3x2TUbzEIi
8dHvSu776raCN+wn174f4NACL1uofQjWSOVgeQ4dNKGjBD49sAkPiN5gBr/XVpDh
kMO9gg7dT6r4tmXB0yzP/cac5667NY6tNYS4F0vJzHbTezP6v6eH+f2jk07BYT1V
t2OVZKh+1AygGaoHLF7sO2zqQ2wcF3Y/OBbJczJojc6qNNYDdaiHCXkm50rETDWA
LaBz4eynlP5ju4/Lm/JKpW9+FIDVTnz2mHZx2RqwmiMJ8kc+bdBOp3DSBS7Tzv0g
e4JQKuvoBZIzlLWIbli0GJhzMS+RNydmRw5DMMCI5mcsJ4SWHKXAy63vqIkxvE7n
ccAlqLT2NJK/tW1inrvtOhaqp6DkufVyhGnT2lAl300FTA3WoKAxzN9mpDgE/BRb
hUHbykfIE8jv4CLGYOa0jazYpppslxi90XjDr5KRo9M3biWWNzr/dU6CgWGUbYtt
7Y9IE6bCxBK5RhxljiBhoAwxCQiFvZhl/SWXCQCFJg14JPY+T6ePAZbQinUcLuOn
4mnPV0def13+0E/iNiwLO9KeTkYSRL1pfN+WtIPJ+7oS7SUEC7beitSlulsee7ln
24coERGDezcsyBcGR8Cq4Y8QrhIBHgGo8vYYHClc57QFql5QjMLgOZcDCw9ZKl/5
tO30Av3SrJuvIbCU3UWM/GMMJ0jjQqbRNn/X/I8/F2jQQvWSOLlRMYjlr+PpTPvt
w2NI81CPcd4qdJ4F5p1JSyAzJSP8pLz4DiVB+WQIudy1W8NYYGvdpIDJnDPnLGH0
VlptQimyA+fRUOmKa2asqwJ5SD0exK07vEM54+Jf5yYixoEyHQzzO45jY5Xfn7RZ
oj4Bpkrp4Agb81NrEk54iA4b1UaZNYHCoZS9QdoZaqaiQo0jy6pE84rEqYGeKI2p
o8J95xpDCmOXYACvgZgs23ZFJ7hda+yY++U7MlfVHrLYSkD7x0gL2Gk8FoY1qkY7
05b+1ADp33so2HM2qpVVDJ/OWAT93OKUPcXnjj8sXrJVsPNX/Ll5VNe9UEmWKA4i
NZxAlxiHHxdN7cBbe0uoV09BYlYpZyuqN4LoxUaRX/RZdgwBt3cjVZn3E/h1REV+
F31iDI2nccQZ5La5rPp/j7eJAh6EquwPfeKh60Hp7vbiP+xV1Nl7QG1BezzJSDqv
8Nzf/gOF1tmGE9aDGLgkh7qZPIHM4jPeo+1K5IjFdc04UJsqcIIKauKxPovW6f8/
lOMBNJw4BQz2zkdbQ1zO/NQQ9oMSbw50KUfRwQ81g9dKK1ytmb9GtPCfEnzGCV+m
G5VqE1/q1LXytEGQtQqo4uFtW363XJrZv3C+ZdUPyuSCtiOPz8ApnT48EfJHUPcp
/O5wrOIeUN+J1Kex5EKJE5h791zwfojohXdz/Y46w3N2SHsmFNW1wJkwwlxW4pwW
PD+M0wdZsubL7CYkr6yN+21P5GekP7oTy+ZTiG5UN6NTYXKBTUMNXQilJjZ8G2xP
WEwDGgD3iQUTiEAyJDmGDrug5Hvk80nAXQSJraaT/8JTe1kBiOrzttYZ3d/saaLM
v+bBpNWtdtDpKY0TYQ6AdQ2c87vYVvvan1Lfr6wa4jVG/r4HcJzF+EgjlsQXUi8X
1YwxOnDqpFppxMDEAPXwgYSaeFlV0hZ41GjNpP/7iWBLzR5PFsseXTQn36htJ1Z9
xvaTc+3IGjSh5cA9bygmKyi/Zmdy57f2/2HkomI48HkGUEBfUNuGv9J+zgKHzZW9
B1UDs0kCA50BQOxewPOHa3e4zZku35Ca0tBxbCwzs4hNquB6E9ZkkD1pacgPKJWn
CokjHjW8o4K1cJCpunjdato2VEjGL7rMOIqpZfK+2cy6JhnO0jWnjlbmkbC8ibwj
pnyMPSOtuu5+f02r65aJNniN/MMjeMj7wpxyRypEQojh7nRn2KXSoahAFMkJvK1g
BMoSq8YCaKog8rjSDQJMbyEZhudogAKkkICwI+mZMBHdTMSbk5cNwU26x7It/PZf
Ai2w2XBL720yOz0Aw71B6Vvt1R2ZxzOKniIk/P8et2+XmAVhBOOsiTUln08khPUj
h/YzCDaQljhzE9Y8wy5ymqVmnMHIlSAa9H84A+ix5TPqogONOTDF/d2W8xCwXcs5
BUirsT9XPTb7iwjU6uIKrBZVWsie/ImDahpBzsz8LtJ/FZ+T4Z5g+eMf59ejlqXd
BGfhco+C3Yl8FigOYCb0yzJrtIqsJuOADfQZQJiHfAeKlOy7dLwJs53utIkScqAA
+/at+H8gbWg2YxQso9jGnaUlGCnGf5ZrCl9cn7FN9/DefMILs0N3R4kFBSfVgE+/
rMmJdoeb4B0SZRIwRMBLDHPPIR5uu0IY5f94AzcHYTEGoGZVV/3zB2gkQrStegWb
OTt85JR2t3BvT1aaO0MJzFrtV18JxoasxrH7nD9KDHJjrmnvW2Ev/QQ4nN8fKre/
qABr74He0+kX5/ZIjJ3kK6qp1xfDc8k4gwRHANJfsmGpcjrmL3gp+GFnW5lh3OFr
nrZYFi+Oe6ypFTM5ePocPJu+7asugNatKCcfQpGIq39IuKgTHQJFZS7Z00BvK7P6
TJI8QOHrCMN71/9GL0w8Uj7NqVgXu6BB+4ztgBtxntw3LCjkfYYo3fWOFkjWvkeb
/Hpx1mXoeYnTG3/lD2qLrUoYbrRgBW0lHh2EO7VGGq/8+keMVy0Q8+ssq/Z46e3F
7yFcamSsQ/TMD2abPpHpTdyZM6gAln8b+b/dSwh12l56rIyrD0uUrW2AT79GFz46
B5zNF9l0K/zy52x1UKnk1V8obFfDRj1ug8I+BMrFv4uEVAbT5DuAlfObMzTioZ7N
f5DJYYh6ID2PSjSlIhoafNaJnp4dHJjuj4w/upZ5CPMbffOmXKyUNcNoISBd1xsS
x7M/7CYGjd4GnebNTXMpCzulHKKMo7iJ47daXt0VVOABFz7xSOpmT530PKZiMx9v
uaPb6BW4pRJ0xVnWOFdhYeuXnOV1Erc4t7HP+T88rAJptfQQkiNjFMcLtC/Z1Bmb
i6L0r5mTUJqAzikMKYcofenoS40N1v09KfGGr9C6ljNCQw/8Ip+xKKT+a6OcIZsf
GJ+uLaVVGhORl+VPlQ+rWMw0by/f+rvoAsHzbP5F4q4P/0cvGLspkni3RiyOkebE
980Nd8cSMVGxd8aZDR6P7WE2ovxm+3MDM8+or6MhFEladCTQMt6A1JOUP+7eug2O
pmXKDUBxjA+y2c8uue8R+ZP6SXy7j9YEMKPvl/iR/xMCTkcJOJ6sQ9OlWJRJNdDr
o1Rr6+FHCuKdtWfe5jUwGt2jBDBK41mh1fHLhT7voyoVRgo2cUxocXIB7YwLdYK3
t8ZIiHHSci+MkTWLInveJe3z/RtQf8SnYVcHPIg2b5z8NquxMtvyu68zdDfEQWD+
NmxohoPvXvW/6uDMjWo33k7+6luQ4yoE6mP0i1dR+0CMzZwfwX2hIG32kTCsFNPN
SSwKV8dvBwYtsi14vFdO/j+O3tp7lCZyLjK1ulJXTULRE6KvBaIiEX+zTBzXmrnL
m5Yg5IvF9FLo6FMfe70aI1Cp2kIdWpup2pYvgTV8x++6de54R5mPr7FfvCSJqV3p
YHCdlrv6SsnST6Eko44wUKbUj2kDtgC/Up7SAxxSK+CHemaqOkDtJGBCfYwWQ3Uw
F+qZie2BsSfxZ941CgxfxzWAQhRyLGXKvtCtVUVdfajAONFv+0WR6Rrq2+6B/mZw
CZ3sfCJsveWz4ubU2PNUn/DG64ehS2TA1p9QR9GPYcaC91ggPTRclgnRD+Aw+uPA
tTFHZRZe1D0zt4s/wp1/vHxsOp40sNKwKPg//LBeINyGjkP2okPQWLKLTCytas72
3e1cDoz/n5WI1L3p4PNP1QNT2zrCIKlUTHDpvJnOkKZ5BSASLHAXOmP9PlCt2fSZ
QShC74StraMOzPEkFMkLjQ9Q9upOS+nfqGjO0LMce2HpxmSla+4p/XfwOX8L1iea
1/gZK98zFrtLp/bYonlsRAYWCY3oFRsU0tFdesWm45Yv+e8uTlmCLfdusV1Oe7uc
Yej7e+dMB2ZHiDGw6ek2sWVcLfCAe6YMl4PZYIuINIc=
`pragma protect end_protected
