// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LVLCN0yZEJNpbsKQ0Q1fyniWWtntvcLAVYClVwhMijvXcUdMFLCnU6Bjbi71+Pzn
AM1+AwdY1vTmY9G8z5WlnZMOjHBa9o9dilsNH4ij92jYjSDYFnTbddYeS/vsPyIw
diefFIfuGS9kiCOeiGF0Id757/UkTyAPwoTC4cDSiU8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3856)
RB+oagqbUB717lFofRhc0qSBKuD1RwmK4JsqYlbUFF9c+4/v22BCoXwS0FMzZzej
5TXcaamVdRmolSfBfk4qYP434e2QluopBbQU7PgLXNjSbNjzCpZw9TpTE9Z11wJ/
KOoNQXspWTuxBxE0qZQKQgA1cFfzZICOBvMbMYMwaU2cyHZYSn675BeDiLp0F9XA
nuR9zGqoZOzqpRv0xtvcgBd6F5T36jrbeWZNV8lG24gCImOdIYWaKXDQvgCLBIHA
0BfHDrA02LWsZ+wE3t3N3z0dHVHfeLti6zpGfP07FFCVk+GJhzCaTJ4JitPyadBV
NvDhPkFVCLcpj1Sgeqhhu15Tc3T8d4kK8+Vzx48ZauAvjvSueT0HWmHgO02mjTPx
9QhpndGcNc0igFw3UZyN9N1TpYBonmvjwdm7OaynZ2wHga7mOONVP8cxWKK+JEPl
y+DVQPEUa4+htd1ylRecuocRARJAwd17vfZnQqytiChGwemMM+uUYofZ2HxK+iPQ
wU7RuyqCDFWwK3p8swJjS2k063wKoJKSbuIHGNa+wlImiJ3OZfGcmrUXo+FftbP0
LZ7tYCIezHUcyskR8dbiaocQ3GmtGjzgM4wgjNIfLIcKsbM8XEshZARq9VTHWrle
yWgG0tFSKz7DySswFaQyYxERmdds5Ssid7RXaulrTTo8NMkigeklcoAC+fgPF8j7
1mWwQUXuleLzJd9L6Ir/HJGtpXvKo5/8tLhqq0QkFlf6Lg8ukSS/Txtbk/mPB8I0
ADD9My2QOzHV8Az8tscH1yVc9LvTkgmzW/b2hFGeAitaM9ndwf8kkemBDM+RyXhd
h8lb2MWjImhx6ktWlIWXalBeFucxylbrVC0Tjg0Dzlnu/oxaMbPez3TuKNi7qm9E
sQ0B09631yf65CU/NguXR+pP/o7hwWcWnrVj/itaXYcvAgjfbz6b7CTnGhcKuHQi
6yIimFzeotqzdnSYL1TRsY29hA7wc56zwgh1oX3tAvCUEosM/u1JZ3+PMZVhxvHF
gzMsCkFrEM52QoH5jHoGMrjScgqkkeEaZYGhIX7H8Zaq9mwMISQ6+IHq26YfdNs7
BJ1kzE8OmsjAV1L4jI+z5zSc669CpNwd0OwLYe9fEENE+FoSCK255b/bzixJWn10
7plxekQHgcYChswmksquQfJ20Ncw9R2w6Pxt5CtkU4J3EKn5XtJP4hI6+wTl4Hmn
U3Pyr6MsHB0+bcEkN7OliT2a3BWbFNmP6Zz65UnwZmhZ6JEOnxjVor0tZF3lkUfb
VJjdl8+oOaMjKE1WQP82eIbGxQwPzExzYTjSOv2Jmnfr0VQ8E13gtTgX5SIlRu2u
XWFKO0qAI9StaYMf7D5YVrnue0dIjjVhvDZW25grffrSPzglrGmFNjO61aue4ilO
enWdVNmJdYHUopyMn9qJX5avalw+TWNv4G4Xnny7OZJD/7qNzROGkRNrWFmeTYTi
Pzjm9rvlWK24DwcGS6vgMK2VGMzQnOCrY3J5KohnqsUS6+TwYnI07+xDew2nTwhq
xM4LRiiw/n6zAri5TZBkmOVTrDOZLF5Ybb/FTuWd1r9kIypw5hBjR7YGPyfWupuw
GjVGVEeWSM7MeFTnMgQk1TpFmwiOr13vGAbBEo4SQzhRtJfuPEM2TmTnwC1uQbhR
tw9FowChIYck8HugXiNdtKKgBL57UWNc18okLBmDK965Kxv6n2VRhJvC20dD0Ej8
x/WLn89UwK47KCy7hGBWcFSvF4U/Zf6TZaPMBPqrMlUkJtcLb6vMPdV99I7gsA7b
I9G4PJoKwGU3ygfYQyNFIEwGqke53xa/oSzXlY887dtGYVh0V2ROOBpTEjRPb6Mw
Qjt01xDPxSiBoJOH8ppuYhPDn5HiVN7/MERQTZ9HTpqv8tUor4WND5hUn+WZE/2T
Vgy2iIDsrGwpty5tUwL3+wdM3wY6perBkt3787oxPNGzVX0ogasdvvrn4lo5LybM
NatU4hbsfvZl955MwwyoxrunGfbw7OD8MQo0pXRtV5XefU99lXgiTzSPZLc7dZoR
2JMYlbz+sdOyrN0qxDjQal6Qeafjt8zBGJzYXDQ6RfskezJRUH8XlTrzeTjhdgfK
Wonj9hhtavPymVdEONAdaE8r52cpq3X2Ck/T+Lw/g631mtB5gaxonrecvBaBapG7
2eAJZIkZ7hRUqFMX+VDxv7dkAgJz2DaWVR5MmqIp1O0pnCepvQcwDiVENr79zHKo
HlTqjgM8bC9zLtpPAqSOOWvhbOiDWgiTpPt4QehJAf/i2dklzoVmE+6BXzTOR3q6
z4OcJsZpZZGb42iREsiaWUGrRkqlZFv55kliunXF8b5DkowNPW5QbCFMU8XyEM99
L/jyVp1hVfrFlPO8KlP1dS71hS+pU3xTs7ozYlZqEYdk2g8GwhzIq3BDhboVesyo
jOw3ZHdKXJav3uR9jdpL4N2hEyhmKElTwA2ZjHfZVHBx35qAV1+IEVpYHeILFFQw
kloGBmtG4nQOsDxxOZBGlkzwYEnMTSJZaiEdyj3gfOK7HsmOFB5CvyhAOk/KW0Lz
BM1PlCthG4rjW+rkcLPVsz6nqQpCuDEm7inF1QsYVz8/8KofBAuhO46YMdZhkZkn
1qfyk5eH0/n5PaOuE3Z/Tu7Zuq5o7SJ3mWYyNIYvgW18Y+ln3wVrKCqRMZeGa8Pa
T199kebusd4aoajVKJEFIchCdssHjGnLudsIDeVTkurCHgt9+e2EGhZKFOS2Sg/1
/i5an2jZ6G8nrgxdb8koBnxkkLfTa24aa5zgYinz2AfXRSRv4PVZFtIGCGC+2149
yXNnrA9GVe8IaTL03RPj72Xh07Z7JX4615fes2WxqkTU8FDQho6af7F8p5OWHds5
yHhJsB+ec6xvFZHMi1vIwTjWdohYGQYhBOG6qXRjEW0GiFzGUD+rD9KNaf+Kw4cQ
GlEOS8PVAQu2Qr0X9dN2cu03FhxXD7RwOM6Ay/Ey+4YmmUHHW3f0b0s7e3c3onjV
eLjovtk4Vt3MjtcwICyv5pyAgJDXVPLEeI0Ca2nrqyDvnwMjzKi0znKNqXrRyFOI
5lSASspMZjdO6+57rTpk9ScTLSpYbMiRBozhbonjdkJvCnK3IXqcQ3T/U2SVl8gR
e8mFcRraDnuKgy84Ld9sDF4KE9pdt2nEW/Gk/HzZMm/JDR16Um1lu+V5fGp/ouRx
BjP0ebWZg7xLaSxdITkYsFehGfmvnyRECo09+bXAA2Sfd8Tx6vdGsM6e/bic0wHK
/DEiQ29a4rC4SexNjpUQOL+z9N1EH0iGSVnoGa/rz/dfWvwPFgaQEtaO+UD/TVn/
FhCoM25y/hw8ty3lbiEn+Yqi+rQ35RtmVD8foBQUaxMfXAejV3JWrNoeHv+X2XlF
k9fLOcOS/u3kJAKsurSzMksga8XsXqScVqQumxNNP9cAiHXKu3t9Oxw6wQ0BLVyJ
nMw6rSU8o8b51YdIPG+2/C491iQjKUHwy+TCAhPc9wBhQy9eWKgi7aJo/UrwE9Fg
zq5OvsEIvKFJlfoDnrXrA2z8vkoS3Hkdq0sRXu+8MW9pAOHSDIGyymf+PUrIAgDF
upHiMJb+7rrqIQY2nxugZjFlBMva6XJHcFJefXxh+tTR6O6YKYMYkcXAaeBQMTVh
Z8zRg0H38mCvBZfpyLlsLhpXY0f95zL5jbviAxbSTOJJInQUPuJb0eCWJ1yvL9nz
89aH98EZsUcp2TJ36AF8JyHa6Yeutpw2xXJyA380dXKON3UN1VnnvRVKbsr0UfRI
AVMuTt1R3TPTBi6vpkvlRbHxDYZ7FjmBQHenWJoFv0FZhY/SPpM4/2TNEdSPnDAE
CvXgJiuNG17X20USqpz/rBF3BP/kHX2wtomRw0ZJT1dsVZ2YGOZ81Er/2gxJRXma
tmIC58o2qSW2KCY5Fe3t/76r8fOi6SDr1hl9dQD/93zmGCkMb4BxXPKHAHS94Tz/
rL8oykp2EwtHKxp/5u0427HX0r16Qe8rz/88S/JsLwyvPfIXvCGp2ZU5fbqw5/PO
AEL4rrXkizfJKtyA943dqI5A96lCRCV4n4GVsljqqradhPSiCodJbpaHEW27gD5m
xu0XC0gNhm8LW2w2ovNcSsHBWQ4h1tym8M8OhzRyoVWCINLd2NpvNkQ7EmVrqr8s
iLEop3UX+hSpv48yFc4mesqw/2BKFHoVGlBX8mw9Vus9oVrpdkVO5ZLwElNGtcGi
8d3YJQNZ5+liikQtgymUfYL/po+hMe3TGUwvmbKXSfNuQJ/n4z2JKE9jw5haOjeN
8NXvglKTBUvBAnr3dh6rXLVsdTbJG3gJEzHM62XD9jQKduwW1MdxjvSZfTXlHxpG
mq3SuYpjhCW0dQ7xiPc3GJ3dpHbC8L43E3F1twJBXqrgixJ/Lblmxhm2sm9UK7yN
EMw0JzhydjKJidNbRt3rw50u1SsFiig9YB305FBzEMAHlWsKsXiprD0e3ZDR2wFV
WAMt+X5NShpVlXrGNrbFr2LnpslkNhUgsGzWxZ2dWH6DgrkI/dR+aLyx0jW3KWfR
41vq21Lnd7sPsAFmKokHpGBrhtJA2lBSVaLziif9myDpU6tJ4HtKNByVxDXCbFR8
H9manBzykzHdSxRaHNrnc68Jj+3PxxNIU8J7+gYTqAxe4EW3a0ReC/1wnUD0vL+L
F7x9yn5nD+X0MssaNT5zsR6aLnoI1HZHDvRxjqwS3+kO3AH8EcinBp+9UD3gAsU2
APQ+OIgy/pyUvEpsDJLxFMPGvFYwjWbf0Rzme8CiG8Ov2m77x2XSxVFkLAmB2HjA
Hwx/WCFBik+lGWxcJ1/ysi71livgoQSfcRjsQJeyRbun7gaThZgtjsJjpMSc7aa6
zPupjRjRLkqff58cGmOKqdU7QJeBl+4T2v9qcXUrtFXuFhd04nKyNahJGeZIkE78
Cz7ggmPtpajofrPXyS6sEf7G1MDPZDhBAyqOrplRU/frNEES2VisMJ0j+MkFPHUh
uKClN6nlCTGFv5ObfJmBl3VGvtw0HMxt6+ZW1wL584U/0EikNPPg5WICaiH1KBkZ
siU7SSpt+mJBX6O/qUwb3X1f+4Z7wYTsiWwd6oBnNZ4tfog+WFUYZ0YKGWXLvRz4
HNBxnjDLDQBhnPnl/HVrSQ==
`pragma protect end_protected
