// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
efmqA326Z38Ztd7casIN2DkLu3sl2edgGyAraTAvgTxMtssd4jF/nIt30knQ8lMs
fIMpFqZzkUsjs12BnC3DhMgKOd5UFyQ4l4bIIKWGVteWgZD840d402pUXniB9eGn
FpLLDpl8ACqzgy25yam3C9LDNNujx0nqqNRSq5m2PUU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29232)
WDmdU3ZAUhg3Xef0vbJl3L9Sg026usfqHzIeNzkQkhZTDgA0e/tL4QftNdc8GCS2
56SbkkI2lH36vYiLesCD2UjflQnbE4qmCLW9+JXyNmz5oSHBG6qFMCOZdrf6NuLa
4N8d/R0rHBeDU30KrFt4yQ6r+jJaF1w4PGKJ5DcW7rqAjHTI7TAscGSCGBMKXJDs
sO7J0MZCtK483Nh12sk1MQ+aO2wkxoyRA+1mm+GUiu1PiwiMrQoz+VqUSVtNFT7k
v6UypugXJqMH7ntydhFteXYp8MMz1Hk8+lLe4mHwXDkcW6YO2US0CzZDSzQCjht8
2HfWx+Iqov/rdHHOJtfwj8iWdbbpuQEM7gAEKudhUwkYYIVGEsK4An4ZjrAN/W/s
8+YKu7X5jilXBTz3M3QLSd56eSy4oBzpxKom4OD8JpoJ9DpuSfMqijguqdAVSR91
+9mkgDFDp0QhN3hRg03R9Rmy0jehhni4mcMLf6FVRDDXPQNaee9fBG50lSdb/Sir
fC74ph//vh9HJRIzKn8VgDzaXGEj9nVwc9eh3nVGXZ0VeR7+rQ8r0m3B+Y/BQQep
OJefhDq7Z4toF3hmGJKyd8F8PifK8MA1uvvO36gyCTBpUG5OwZ+1ZZo5asDvNH69
HUM5ujblbpntat4220qhr/cAZnjzzy5GNHyzEFcZSUFx4vJXWD2F3dNuNVDDyR8Y
mvwe7T2YIDVdzindStc5GeWRQv0qFGAcv94vFkRIomVV1vk0RHUrXnHZmJnP1K6H
VxQjV3UJyROF/qMBYTGnOPNMNdZbTMWH57wI82YAO5beedVfQmAs6Y74iZsUor8m
JmDLmbS1soVxqC+Lr44DdF2Sdj3D8WNDlzUdBgxWxkvcqNrgf44MHtGRFQ9mABa0
FjRYhvD5DD9BGOBEfoH5T2OkjmpNAox2dPqsQM/u2E06oeTFnzO03bUB3HhRKAIc
a8WGAA962QldC4sfqKDEujTW8ebYWPrqiWSLL5uNoPEVakZdPrKttOTMTg81uk+C
JUT1F0TrCNEKPE/cH9hSETnXYfVkiiQl8YHL6w5IQ5sGWo/eH2j/GoNwzi1j5Au/
y4gLTKxTfpIbYz8xaOWpc4yiDj0Ia+78moGmuDtvJV1Fc7TPPL0FqKGbeJt/abcE
aYI0rBYQnqOh8oKHL1Jm47CQsS+0MX3bvjKrFAWApOPTRBLV3wbRHRtDC9C5vR43
d3g7doOv2IdXWXRGwt59l3Gc4H7Lf1Pl9AaiYgWPZpBA79S1+8VNj/ErmBC5BS40
jWn3K3ksc8ewNj2fX+iekncnLfvARmOww1Fs/0SO/bz6La1HXEYvCpgOPB8Y4XX2
htMeT/95tAstIHNS9xjrWHOeRKCBYEc1Zt486JhiWnLZ3noGkgesIPAO4YFczgHX
kwanKHXEynTIqnCnb6MBPP4V4lL2Jn/PhzPvSq/9C9/ok6JfthVpIWuABi1iNQ3b
aZuhMXwGypGob4Ht1Q/8Q0HyX3UwwFCDuHuCvWD/JNGzEUG/fYUXP6I+RI8z6R3j
OWvec/JOC1lErU0hdm72iBKxMNIG9uBmJuiAdMOkeEkiRMs/mnsIHDdaVdk5GEXw
F21nKyfY775Z02eA+PI2EIKLcEaXHLpPtMdb4xFqFUOBgivIr6CN4sG2CktXEAmj
7kQDfDw65raDrZtUCTQREaSYNPS4gsM/6Z9zs4kOBIusVJCwFBJRSRot9uMqODGa
2e9QLQG7UJjrDtZ69bygbQcO3Y5/APw2Lvgd7LfVGqZ1psHhp3YAVcSGPnhp0n19
R38ZyyJOKnHHHAUkqJQ4rL1im5hQzyndrAot75BkxrN7F6vSE5FycffipMMPEFuG
p4aWzZnDcVCarwlvSS5EbdqmWt+CBPUYL+k5EThr2L0aBauLMXnj6oUl98f/DVrZ
MB8Fb7D7Hx+3M0cPchhagY6w6pPdp+Ac8dk3oWW7rkrq1mr/CK+NCt4sKDVZRV76
rHi3Iq4faZrQqyqzG5dLsDdV54N6hHfui+P6bdeCf8F5bO73w/doCEmfS4DOu3jd
VTxsrOpOgfJ9jMmkHmVL1C+pQeMF2zLLamGnTQC79BMRlSZi1M/OcZOdf+nSDbty
XfUbtPrlEFs4YbnPDeWkS5/k2LvCYJk8MM4Uo43oC3eDZmPkjSSB6prb8GXIYAJ8
+kiXjcYu/Faoa/3uw/iO4FRL8DaLkQ0aRYI4aSN1R7T9pLocLFNIbJvWzRWaUtEH
gj7s23qVP2S2SC4EoIh9Idp3FPAySfjt6NYwxXm6JKr+Dx/YIdJNtc+ti+iQ0alt
F4+MvXMMX9n1BFuu0di6XBVQz5FBwEOCZtgQydf35vzfz/gLUBsSqYrhVZ8f2sBL
uHm31OqTnckEFydQhF2/MBQPmGtPDnemnome5NCE1aeNrjnetacSAbhOXQT5GvLr
Q4mxrCLRalFXRpZPBPoRRQJAPJY7oO1HbwIpiguGAW4z3PNzMCdCxt5uXKXezOlO
bf0hlbqyGSCWIu7mbHztKhZ8j1Ur71fot9XzzzLvD5IkDSjBiT3W72EBGwik70zQ
doiUw1oFE0Warxbn2CKtlB7wzzDVFyrW/nlMChdorBf7QzvUf9PxlXPeHBtut3gt
sfbTXgvhpB4oSknE3o/C9FcQM275xdH80PxqvKyD92iFnAvf6j5a9JGxA20IjB7A
xdx5XCV8DsPoJUjizD++5w01sgDCs7HqZaBLId8PcdkHD8ShLD46ZrmMQosvV0nl
eRNhUBbhWpyvMr8vCbVscmhkz7no489coLpmyt+YCAOC7ZfNCT4uW/B8GatpZ9Tc
vne32Uk7a2FbGL1Wo3gL0m+cVbdYSmlMxoMPP1dYXMo/aoehA4EZ7vVUxEDLfiNm
t+7YuP+f9vaQyLpPQX9NbS44ZUjC+08jwH9Q97qBnUmdgG0viBnnQUZ+oKcWsvgp
fshY5gs+lSy8waGU37btwPUHvyizuTZ/QeKo7vtXxev+HkEZ7QsqceS/4dgfd4Fb
ScC2y9LCbey8VVEA7Gm85KWXqh8s9i3djJizfJD+PHj9XRj1Wa2nKXKmZkQtpO/T
2JstiLsPz3hF+xmQLDgwL5VNANLLUgo1WEEgjxIYQoyPFg3353ZXtkVi6gvuk1hM
uPBfx5cGpr7CCXb7tP9BZBID7CcmdPsxrv9xvs+V8RkWqSBjzwyHAzriLFXMLNQO
TBWgwNDbdgXcoa0j9D8BSbdoYkC2keYlrjsZqDB0Libd6hVSgmqvKl0dNc3eqh+G
IZtbARfGf/d0qWiDRQHSgwbJwpuTbf4TUOuqD/6u8M1/UUovbH3/fM50Y4WxBUYj
XBCYVYsoDvGewvwA8AjFudi2BXrTi1wM7Bc29hUKPGKQUzNSXTZ5QbpPqzN7gmvI
KRlRoS/1j69dQWJm7ciYaW0RsKsgGa02i6HyjVyckaOUvLuNh4R8LFAks4iLV6XA
3tVZDtagUmiMEBj3D4pLz+V1vQIbKEhetKJs+CMOrsrMpWn/Kz0438NHHRfwZ5fh
S56m0iOtKSutYvg2YoDfRzXPZ3VQ3lFe1HpYBY6TySgNaKWPLx/aTvcmpWDswSUF
D8E/vT0+ptJZbrZGENu6x0KAToY1js2pKb99duGwF0my8yY6Fz7/0vxU8Tz2KFoA
ZQxuQXQb8vsa+2yNTunBIl3F+5wl4fecPp/BcwgKe+LimSJEd0udZSjWad7rG15X
5pEIhG2oRAaH/GJ9q/mX/0fZV5umrjtjdicEnVLQqukVyVjOz1O8cS2ivIW2ccMr
meBi6wzRR5RnZ42ZVrccAYX3Hf+mOCR8NHUgYjR1mZZjlEPIfFDX9fvyOmCAdeXy
ZopLhod6+Cm73bFxmHCt+6EXwuBnvYIlF78dF1kw5FAxXkvRgmPIEAj/oPcPxRIt
/VLrF/E4e0SKWhahZftAa2Iy6tVnp3+qt+VNxLq2sQbT6rKE5vMJhyvSnkZ8WH0h
L2IHpS68+sy8rv36feEQRo8i8S+7TbsOvkCY1qp62F5q1zNLflvSe1xikqNOu/OJ
WCvXC6E/3zON5wJvsl/DYXxCkkAiiJqR94PuySLGFSLe9HXh/0Kehb6vYghux3/w
EuaAtQ0viFWOnrryKVCxp2MrZD272v9GIo9IIqXfwZITXRgFiE7Hl6RJmwQapd2S
VLgslKPqvJkz4Rl3luSGXu/5YrHBJLAZ0aTZ1idrZgNnnYC56hC2jxuvbJ2HUoCU
P7Lv2qZx70wSEDkYjV4tfv1TxSU3D38kaYpmBl2STJwOHvZHjhuCm4XLE3Wu5txn
f2eyH+URYHsEYOQCj1Ns6rqmmLiH8u0a4xd2w1tIKrJ332NQabXkUnO3oXUj6+4g
A/eX75di16hDUkFO2q9P1V7pygIjrTxUaiWdvqVYqWZyxLjHhc55k7WLkkxYQZFw
Pa8Oh0xN7CyfqoQM5h6jeAZ2kSoim6+JVgW00qCuftlM6V6aj4GdlZZTy5ZvZOUr
vi7YOEvNC6rsqt3FeN7mbhKENtLKCDtCt+26Z2CyM7u/bvIK7AzhX59dxPOMsr4P
nnFHQ86rpRBJGqZq/eejDHaUIHis8TWi40l7uWMJfdAZWnW5xgOY08PJPhqMWxX5
wT4MpROZabLAFFd7Zdn3Xt4n3iDYpEjRA0hBO5FHhtBgpUs5rRcN0PIGWOU1d3rE
6cthTwTOhAX0DwOjMXtyHw5mdKV4GLrWYVlaGlBt7K2lSk7CbYZgzMDUR//mHmiI
+8ZcecQ6j+RY09lMs3f8AdfYJ8JTpBshGJhF/MniD5gizl1ezjgaxosu+exOQ/Xu
FlQBwc+sXQNe9RD3hQ2AilvOL3FvSbXBmef3V1P48Eib9Lx1wJDTM3IzEU/ItJZ+
NOq0esWJ0YH8JhQErXCXK3p5NDyHySQtUrl44vuqp8eSpic78ZimYpmCKr9JEYXm
IWJenJ3WftHswbstmglQQJjr0npvqLTyghc4VjkJUQNskyn8/tmj/AU+2uD9dDQ6
PSWF72Xtpg8YY5d/eSGg8onBA7c8ysOS6exkNEn9npS3+CQ9rA4jWiIlBs0u4rQn
GngWWHSnKskNeWJF7jhmG8PVLcSJgd1Ta4ihxzDOS6NIdTL9Y1dT8dUfUUts7tDn
3wTAVwYtfzAiKRAqs1YfZzf8EDDAAeFB8ymUwcSza3dK2RgwxdpL+JfrwpDVRIHm
q51auOdEds85Vwl9DqLkfyAwas1UEZMmTTuSSFMSXnClK3okpgl+0ZkAnvb5kir+
NAYyLfWAfPz9fp3OAglNoNlIR5vzbPSU5glA6iA+jrMjAUMwLzeHcEJe57mpEpzY
UM3mV4Xeh+DUnoLljuczTspA24LXJUwDfcGBAB+im3E+qzJGPud/VB/t74JScC5k
uMthLqGnk3FeJnaTCF4qkV1vwjJOMUQkwB3sBC1zgWIUP8670ZNSo9SyVFGnb8Bb
D75V7jlmIxwGLALf3arx7Il+/1WvI6+5u1HS0gl1Temsd1ykQS7XfrFWTXPWhYBa
FLjLTN1YYAfrsJf1C1ZBWjrASqVnuLLWtFyi29P76X53f+DjFUMg9h8heWSlw5Od
9IZmw8RDssqG4MiLwPbYYj18kNhRHQe0juSdT/omevzPgWvdDQSSQrXCexcuSFur
rhjlDscMHfGN4PjcjciHlvIr1vviHGrAVyTG96G79PA2NrZ/lCpVlVE0Ev9fFnZd
SvHayOkAV5ZA7vacuRag0d2KRWxg8Mbple3q1J/HxNCaULFYIUioaoDvIAw4DWyU
4BxV+RLdVuQMOJEh3OdB/L/9+RG3iMk4CHmreomcDL6p1te8OzdlHxmlLG2EmvIB
BWNkFy+xsNTfocjLlMJSPhoVop0KzfY8INMlArsWRaZU9qyDUcY+QNWS82TvZSgM
/fn8k98EyoZVFtoBLAj6586k7IuvR7veJVCJMC5P5HyCYnuePIne3X9Qeo+qLQ72
W4kgK1UnGOVpvD9WgwpHfPwXZAcOPzfvd4kmYuURFOifzffxQsvBFSmoK8loJ5w5
9Zop+9V9gtmjL7MUwOyeAhD12LHuQU7DD6MbNhQOPOVPeeWG+I0Md4m0a23Nr/EL
0T4svnMgN2N4y1u+GyVOYh+blO0xoADkuC3wDa8/zlU5uoMcqBJmVtcXzY5HDg4L
AT33N1imrKASxaVlYo/YHXR0m8Pga8t+4cfgK6BbTucuCDIhIbWrLJXxk9BdFn6X
Cdi42H9mDfqPK9eHGFE1o9urXvIAOcdiWiipwE6PlSuxIsQemzexPCqr9IPjo4z6
gXhXoAruiGCE+mSJ76nnmXe+e9biJllhKrRl4HcM52YT6K0NAOdRzEN8LlLHun/w
devae+ZXEPODBoE+/NUJ/YVwzWVHP4jHBm2bAdWCIgYHas21PfYukG0hv36sx2gJ
0T1unbamldMF67cGVsFIitxX4YCC4+J6/iC5djfZiR6MbfZuQECOwZ8ceBtgGzdd
NtoEVbsn7zcwhbKCKmpH2+SOMMznWEVoku3t7KOfBVkpEM2F5ubU3goJySytKSqi
UfYsSA7MqF8SOjr++Iefg0yLBRejqYFpIVOAsXp6OAfU59Kiz4tObppqI6Ol1SKr
5zZA0yF42cIn6nIM0BrVHA59dUFI5OPHUhCAie+13ieAtsGHuwxuIkumjUuILQgj
PbmIAEvI0qknhR/HP7GVS7v30dns4AJRXmyCVhpC/F2D7Rquu4b1t9A9oc5hh6Wu
qzEMEiop2KH18etzaNdwLLv5qijF125LTWqL3tB/8kwZYQ/7yHHiZ8U6pMpS8B/e
DmqQwQPXavmfOSPqMWRTmvZWCbJI7RznXV2Aiv2ZsjHYgBf3WV4aEHU0Shc80GN3
fgcn/kg8hGXWbpOeSfUrKTk79uDn8iVgkgYiIVRTxKDlEGasJq3mOYRQMDNGioa7
K5y/Erxr91Myxenp5Gb2L9VPuifH+AlvJXXC88HvdvWT/CWW5y1JBfNlrxlY4zLE
jM5TPkK8AXfAmhf2wznU2kLzMSz3ArINoYHyTntBVnWAevEySjSZPCieSyb5Z0L+
eSyGBdGOhc0ud0H1ivqZ4Gv8XTa9JKa7ofFDxz9tdTfA9O7zuIMqjYEyeQBvE6yF
NG3vUlS2QoofbEHkE/pw5LstpCXpPrG7CUmH1KO2ZbbVzK5dr/cnnfTbvNg4B0H3
o6B52HPhkshZtdtLCaga5zQd5VIkokbjFUzId4VfdRP6+Bxw8DILrvqXZeVukJ85
QXV99JWWhvTL+cADrXuUDU0G+W1HzWfUGamw/39MhpkhnFylMRcbvn177II4usWV
OJR4/avB6GhIuJIBLIIRojHEhJvcchgGfDhb5DkdQb0jUXqXXujO7zs7YF6SDBoU
gKcRqCsoduLYJot/nWXf4wje6qvWZxK3lyFKocZutiqxHca56HmQlm00rnxAtUzY
E2nR6fRAM/znCuodH8RcuZxhJy458t/r+QiLQ1OkB1CNOX/MgeW1WRl9Cb+zwOt9
a0VFBm7By1rhdQee+Y9ucZO15zIuHbKhxkomS2bz1MpYv7GTJQ7FjRUsN+FgL93f
l1/9Ek6U+Z3yp2CEVzMYEbuR7HP5ggiCi0yxldK+LEt8KzWJ2jpSs0KWMcd5gCxr
c9lF4AD3uCgluvotR6CMrby4ytwLe+s6xcb6AJfRoNCOEGfOmV+sa2u3QoC0WITs
x1UiaW+1As38yIMa/nu+gxSMB8Ctlm/hk1YjGkZzWovAKFCht4oQ5ChrlpOdRqW8
AzEVubOZ/e+31FXg+J8utnWoCXXqNYYJehbBA6eCeMdCQmDbNw+sqoZ0A6QGBYZ8
v+1fdb63fSfqL4MxjbTaJpGmZOIMGm6IjaF9K8nayI0B99GTlVIlXyhVoFWddX14
zas8o+Psg7BxM4vQT8f0fVD5JyxVVxm8SrhNDK6bzl7aC2FgrI8IDrsKd6GvEVS4
4NgY/LKIG68EXSb0UkL812N7K2bkVYRENrEZHX0P0kCBd5YrEjMVZRwNFi6KB8pg
HmpCkT34ZrxgQetfqdOEfIBBU8wXfysL5W/6sEX5DEXO+vhgYsfjvvQj3dQPKWI6
/LFhcmDLP2WtE1qTptYTccPsPM9h0e5N8sWYyTH2vUCJx2bKlxUzZJM7TIBWFEeZ
CKtc+LoGJzdRmYA3L1T+h8Hj/Qr2Bf41L4uOfOLd09pfEpDkJ3vDidqVCz/MiaP0
IEwvejVRa72gJ1S2fFy7cmle/Q5vn35eR2OK2AIgLLuZ+pKU2UelmgwIeEIa3UNf
ujM5Yi9g4dv+UKnP9TBQsquWs/c9gSZsz1JXGmoJ6qX4UeVyCctFyBfYJf+Dhp1A
1AQIwPCVE6WB4xzEncuo1apW0Rc4d9LmYJYRcTUVK7iUWssXCd/3I9828iX1tnb6
s/4afxKeCTYTQqB0AZ2OHMevXfYXHaIlaR0eoD/4C7a/vkuEe/fpmVqAL5f9xbei
Lq24H90T2nTUWgz0aAFEevCU/Wq6nSYNf5HcMO9rk3vrxhMsRvoghb7nCQDieC+b
32LhzJ2mDZW86UVKsZ3+/28rtnVQd6EiWPGKfzwkiX5UFWBG5WHnf6QMOLwiLNzy
I5jD8ezJTQBqaqRpVBZerzmob5ITG5/fKEEyIvk1XMzzn4MICd9Hw3k6pzFKNCpi
1lM4yd8Lw+mrFXpg6oYGMVIVlRh9irqS2mcuJhCxG/rQj2334x267gbXBr5U6Dln
0ZwvJNGEIb5gjuvZXtNdzGgtthoh6n2ExhkVf/36E8DKbS60oNq6zNCYJj4ioKSw
87+RU3sUu+ICHlqFSgYhbe0pbrL15YU3V4RLcq80inpkU5pOIGX5AO9043Fdigzo
2s4QWN4pie1uVFgcCtfs+9PGgWxFiuPLF3L1+mA3Xjfujij5t6tWM+Y8C6oN+qBh
MkQBx9+zzTaZke0ftox8BIay4ae6Rbh2oP1oydLjymjtVTx7nJTiAM9eS/QLFLxu
K9txBpIYBpge7Wgs7lWfozZXDf2X/MukLP76cwxKeOmSoR4wbipKgLUs4sfzlR7x
VXLeHy9jVAWRHPyUbh9uPb6RzAVlg/Hg+koWnSUv5SupgMlLZKcgNKyJWJStjNAq
IZtmAHNkr+omAIUontoCnkpOfSdumk5np2Je87arYPjFW/+w23kDclkdZZeytD5d
CS+IijRYv80ZEVz2sJIL4ISRA2kd3Sj0gRPs9WtbyRTVZA5pHNHPCGRUmaEFkfol
i7No5R803w2xZOOQX0jEW8HBtAAbVVX32+0RtmYoe2cKQ5U+mYV5sc1+t5VDsMrF
HjGS5FIDwiOVRF1LfvA8TBteUcZNuJH2cIEzCj4gprNUVKKHskQ5sXKicJuBYbQL
ytehhbF1PkM00yff33pRzIte059nP6Exxc3D86/OssN8D3cH9CNHcYyjc5m+q1Fg
v60jpUkkrv+FVTBfygBa2ujaeiQwNwsqcheIEoOhsBTTBYU6se5d6goGV+NM0ZKc
sagguYrhsRp2kU6+8wVprZzwDpKtM2MvRv3PqFjai2AN2dNatuk/peOwG+LSqw/y
Th/UkVIy5gbIOQw8ZncBu1VWy1Xck1mbXAS7vWCgniID8Iyewrm1iAxDaY3BpaEK
9f8KVB91vX6/96nOojwl4fmQk8ZVhtD4WFvTtSBg8fsZBXs/DNUOJ7zK3eEaqRIN
DvvL0w4e5HF+Ey511di7MRxTbyo4XIzSXLqzT7Ts36VGobxSA41R8QtUdHai9OLg
U1Uw0ShfcSUeiDq0bHrxirCCiULUX+ACKrnlTXBwdjoZDzKBdsgLXh73w8l9sNVQ
sBk7VyqkQLjfLsYGhnnaSDnmpnZ8h40T3ubW5fK2ukKqCKn5rSZCcyFbp8jSnoXd
UhUHpbzoqyk7VAVFQCdBuhlbvB8G8N33A0qkE9wEL6R6WKMtj5VG3DfsF3EWwvBV
f68SCuBA5M762SIa55b7E11oZF0bpw4J5VX+sCaA9FtY2NfV1aeZ87C8IkT9Y64o
EkWTZIucP4EyGb6pmvLdsWYV855uU5KNidKZ+JVXwHgRSm7K0saKTSL4iKqQpDen
v09ceozbjOxYloJ64dLjGivxXA6UGzB9oyWQJlCL8rGz76IcwT9FZKXJG2bnh/PM
7fsVeENtLkqx0R/DEYHyXknl6vV6BR5DBTeBFiJc1b9KbkgxPFcVwyj2Jfnf9LQE
GSMDTiMFzFideEjr7gTCGaQI0wBnZr5kbOxDaum1e6XC00ENe3P+QV+hOU3MDuft
faJrC+BvIRFWuzF0ttf+kRgw8+29YF4cxe9ouulC45ikXismS9vSPnj9LXWr8xHH
SeK6W873kpHrOxUvoXjDNuFDK1yl9yiRM086yBFR7443IH2/+boJ9rJYjaVTDo85
2h/V7pJi3Plv8I9Q9kTwXkSom5QToKIjx0l58gqBttRK32juT5B7ceNiZAu37U0h
8R+wM6tRK8ozaHmPKiUrwJ6GorNEdf+f4IbMmZKLLBsP6BJ9l1Ip4esQnp2r4AZ8
iK1Ao08QTztFQJLnXb5lQs41bw8QVaE9CdPubrwzjIZqdF4B1KSl6MENyc5ZSWPp
SzLisq1y08IbZU2LGsUjCCQBRjgu5Qrv1pdaBmQEz/T3DQY3gNBP2yi6Ysz+l+7N
FW15KdfMZfyM8IE4Ig1M3+OVE2FYNUCAnA4uJcgZPf69zvyaBx7/A5tSh4Q+ixTN
q+H2l7qygNpzYqdP0NNyS/amSF/JPnKXYqr5HA3kBFsWXl80bgZo3wiBWF5+DogF
EYHoyS4OIaKU7JcMJJvJHYfTCUjlNIH2dHhrRBqb3SPCAvBAgE+5GJJr0qgHUhoV
zXzVWmgrxErVcl4ADRGefSzjYkA/Z4T/7IvjoCb6FgWMUzfqAI2rxirSqiowosYV
f7N5rUMREgmnORtdwn5ywMfvN3A6FwGU4NInTDt3mTkuCNwITd6WjuLZMcyKlIss
Us384Si4OHpPOkrIJhKyQDqDvldXpYd9cMY343ZO9Ksn2zvVA6Bd2DY/8pC7d1uZ
IH1RE+B0xxUx2kJCeSiUbL0AeUevhoHV5Ic+XKn9jfThK5Kn19R4kWjvzAGpWud+
fz2x1gAfDUREagQt5lXpMMzM4bQ2kc/zbiuPFEcpnmlHWdCG0d0FNb3hvGasNLxa
e2r33s4oWPHvkG4AEtNNu9tuK1zWSrF5pvf5mZ0QD0J81S09OX17OTO2dk1iGoFh
U/hdcUgVPR55tp9t2drKbhHEocN+irF8IzVGz2oQbWlsqfi4+tdRvkFYBZcyWVtO
wJfK11DptP8fuIF6qVTulFJ8XEdKWAdjKCwOKXv8pAk6rXufaIzU9IozDD22qutO
t4sxyxGwvhkw97MCk3jjwqQCY/A0yl2JtJVhkhixg0XzejrMNJJCDCo2v8a1HazC
01Vpk7pOMSJ59PN/1KJWmEJ03YyeH/prYlgH8HTJ/RZDDImzIGJx8CU+yp9VzAHs
fcRcNIC4WDl7aOhI/8gYnhwo0dsmA6ynnW0pPnkIWHRUFi0UHO47rqUJ0/osQmTT
gk77pCD6l4NxEeBOCYbaNMKFwCETNlGUz+VGmWQyPVn3o0kcPtMIRL+YOx3jN6RV
4oOOTKCusuHP0MZECpzN8xW2B8svXB/vpOQeKZ7V7qnmycZ4qjRaFYtsxj4V8p/j
Y85usaibkSZYRtfxhxsuWjyCHvqxJv/RvPy04QkBNkf3JB5owFdIKErDuEX8jX3x
gnMMv9zLp5ELPIXKZ9fkKuZfKuqqTFS+DyfRFvpBHzsCRS2P19SHEFy0r2Nqf51P
XDRa2C8shRRxnUPmyOdTy1LyfToa13ihrPtY2a3ThG9db/219XKNLPk/J+te+1pZ
+oujV87O41Hy+TbZIM9ejPn4ZYHkkXeJi4VJmMgtqZgH7RM5PeF0bUQthRwy/jMI
b3uJrh+huYtQlOXwt3kWHNyUasq3K+88DaL5JZVu844Jf+M5sU1rH9IAtrp+W5g/
sOPHMoYY2Lnbztls4zLbalYhkQXMuQUHIbbG3iNgircwZc/gM6F08q+WQv7xhVp+
/v0lAXyM4qnnJCVZnD4+1X7YX1fmKAFcdGi/J6/Eu79KDFkurVzMWnHOwE3vN3mN
6u9cppUOQOcSjEtx2tgRSCJOD5q4VWlHULBiL70X2y/Jq0S8x9gg4p3auvi7jedL
/1MjcsFJytWPPl3L4or+R2rAV20qEIAlcvJmzH1qkpuzAlMB019q9iPSJNYOoHdw
N3ujbUf91Six3shvxKQJHKxTIXvM0ATgIMqv83d6OdlS57TN56bS+oJ4DItUX2ay
Icjq5UQKFtuBc277Xl4GbM3Lmhw+aCEIWcCTUunk+e6BiHKibkVqVzkU1WNd61rZ
r3c1Xe/G8IhSHtZiK+sYe+uK/ABGXny/CmtTioT8cy/8fA6+//U7/5R0D1/sDGOL
ce2sdq0J1XJnnFv2QQ1ePXUCoTYjyvATwuEHk5AlGKmqXLATO5fL1YjmT3BRVSSW
QvvnS951JNQMOzuPBvk+Mog4pKhyUP+5Qj4xE23XEhyVsJ5THRRmUKl5eBJSe6yz
+v4bZgMchZY4kkdP/teJr0R3YkdQJLYdOfsW5aXbReI2IzBJypKwdVzwKcjUPCdA
r49VhshlwBkye8oSknhaBXbLZXqcL6AXxyKuVyGZt1+xwG4pVX4JhKNtzArVZjAx
sZx1zsnNKbiWRopZPKJSwbRaiLhewxrVJ91BR8stSZYTFDYTpqC0lyrULp2wVXGY
n/dNnHnVV+JzoDckwSckmMgLqNwmjCbc55c+P2gvrBMkq+ikM22hFhNu0i1IOlY8
L67cTdlSo2VBx0k9WN8MOKpQAhq52BJ2PsrYFgmrZcQ/c3FWHUju8KfwOzEEdFUy
OWnkaH00qkxajCg0t0WMLK9RvEZj55oS5JDxOPQGQtQkhhS7sscNKlWQ6JnnrANt
O+3VNwsnEM+dYewVpPTRiVkYJ8WmJ7u9mlXisVA401jp5Ewt+WcCCGT6+BMQb1QX
2v/0bh4K9OGjJjUwPujS1GCNep7XyY8m1h/bq3c0ZOnkB0+BHjy3n/cwOEoeFHJM
EiEzU6W32JQT3wvJKjkKpS2VBau9Vq8OGtJOWrfAu3Ds48x5Q8FqN0qWJh0QeHHO
EQiVyAHxYDh/X7Opii7MdSJ6JF3qialovhW8Ax3YGd5PRmrKIRq0BYO9ozKG/SLl
gxtwYwQZ9IsoZZjjKuXZ9xqM+bRVqyWGpt8kulx3Jc1UPeR9VLIwJEj5CMv93Kmc
LXEab29OlrT0jrEg2l+H0hW4r8Q2mkaPbXBkip45KPINJXDQAZO2dao6aLCJz/3i
71HR1JBIOUcZwCDVVXDL7zj4gJ+SgCtef1R7XrVR2cx6Jt8bXUSPbH+zYB5eAnim
YIfdpxkTQHp53GmEfi3HRNrApBnk5Q1vZM6Q71FBdf+xBtXJ4YNkW6IRlZxRcD+1
hjivYQPm3MJGIUHhvr4CDzS4ku1FdzNc+4jV3Io/GA9Ua+T4ChxQTh/YB/CLPImW
aL56MQiH5eQGmQrjJ5kCeZRCZNDgIMajxqYyTyysc831S8qGZ+fiYSpPasOVh6SO
x19KNBA3C2ct2KkRgPhN+bIkIjh3KtoiPSTVsA4fRGzv/djF03y8Y7QQKgPWNjPO
q9DyRqe8X8Fb9tQG0ieFRn3AFGYAjXcRnj0h7FF+AcxkfoCOPlR6pwD3wfjpdQVt
wrLB/acEle/CfQA76hTzyNc/cnpKRios9ay3xaBX39i9hEzX0m1i2OWobEvP2gJl
FJjCQellEFa7t+NEnYBC9AYvSAhALLzuaAXnc9DjcIQ+8/Pkd3RsneXLKZrvypcL
nbR8wthNr7nXS1MDwap7rZ87HOexQ6UBwjmooDLlN8rx5o47rGepRdnxSmyL27B1
AE8TSOofrXYeWWAyKU7zBVcwngUVHsL+YXyfw2tVqK4pBXDTsmfye8z3JOxgHh6H
i4d8G7Sanxjptm7ZgYJhG6YoSaUI+0VHgNX9buHcTcb7Fl8fl3M6Lakf15YjxmS4
r7+BdppO6ZL+kQCAwNcE818xZlL3PD4uqcoADNFt5JYNqkKDLpCMBd1iHNO/HuBp
Rk2gTu7o8IJMcmfLt8zBf8xwKUidfLZU3ZNz9uWvz342vqna85aXCCK69n8UGQWF
cwd3sqfkGxdrFDC0KIJ4M/fiwANJI2QUXsRHLSZUl6jjUew+JIEhTmbMWYhpn57Z
k7hNQy+hhrKmIBX2WLKsKFefl6QTp59alWdgOR8AJbfjEe8fJXgNuRjrhvHW4wg0
vUddvwBlMU+QWJWYf6upB79svQCUWNUSAmewSsnRK19EDZIoNwW3lKfY2tLKlUBM
dJPB120OnuJJIJb5nUuZI4Z1vP7ok752OLrWqryQXgXNLY17Fq4Jk/5z3nSpbn75
E9xRWXu55QcrQE3/vAWK0vvBNBxvmrQrmB0xe9Eo05EhHwffrFocCgXDglQeL2wN
Diub2QNz1wwV8K/g3BbdiJdVhJDmRA7e29n6ZKzcrs1didiwoE4rhDjTb6RBtcSZ
t2jhZNBp2u8qhZhQaNePbtItwAB3KTef7NH5Xf/wXPtsn2XSvdHRxhqOQuw0dIFd
MHmY1LsncqKT3VQXY0+KMGq1XoNTQnPgGn+97NTclCrXQHBdkqurIHy/TrzBEM4l
x7nZGQraIcuegvEfwFHrk7MDYuG1H0T+2MriH47zrTh4eRfiQ9TJwlpCkomeKIz6
GJoFmmHuk5Nw0qqteV2qFQVbi2J01jziOI/ADd1KdjWXT93kQSNQHmoSM3FiwuQH
V+88dsZH1xGDl2Lr6CtPNzQ4V/AocStOIJwFV20UovtFJYFpTeDyMDCsB7dIZIUe
zFOIjJ8pMP61I+blQiPexjNhJ+4zNxNw+zGixLvO2p/o/P9YpMr1PcNmzIwxY6R7
r0BlHaGrcGDD6wgYLoazkx8sBk4zo97d9CMeGJx/R3Q3Z14ONy+b+HEhihBAoL9t
EwHtTyAstXcFwLmDbkFGsEBsAZp+x01PNwd+k6afAJfNzwbeqvyQtDn9MKiseqpI
ed2G4pCr+CS4OdVEqgxyUvHftZnBovNkXdBsmvKq/tcloanL8ampqmCizHZg/I+r
2gdwoEjEc3AMi3/sjY7gOD3qiKYeVEU2LjFXcTpHaufpXS9E/XJZa0rdttCDvkD6
pQvdqX04A/N+KlsL01V0Wtxwu73/GhzFWAGAO7AP9eSx7yg3MF6fQrai5pYngEgL
ZIGdRhR40XR8iVs6yL6yM9tKZvBmj3PM+/IxVXC0XPHcFSR44CoQERXPmSpAY615
922l8OcGjbXhCXIJ779qvjnI8+QGe9Tc4P46TIRGN5oPFwxmlBnLFPWp2RrsFD+9
EVBVIUl3JPUIF5J8SEO1tTCRacAh1QSH5sdla2TW8kqDUOsJOhwwHoQSp/7fBV5s
I35lWEquqmxySidVMaJmodFuAPJwnKiVPoak150ktmsXHkcyfrmW4cCNuHdQPN2K
VF6W7Sz7VgHaavNtjQO7VE25sBg0EZbO4CFfy6SmQ1sTEvLoBoXTxtqlePsZtP8x
gtcLD7F7BxoV74MYl6uxt65keIf6r6wDwTNPix1ZrwQTMUEoUHVKo8oDEBXO7U6R
728Rk+PPKYybmwXA80jyRqO4LiBKLdJbTK1hxbSQylGfHmqMQeVkEa3VGN8phD3x
2+cLVEr4xL9mjX19Ju4xAlJb2ej2DZL3mFXvNHaV2O2xfjwDGbE3nlJsKJWCNAnp
agBaEUSeCPGNvn2HJQ3KILYc7XBIoRM67SigNxN6c7oGhf1bzAq2XnsGw9/BaN5o
seAwVccndzbQPt2OdaDp5t6Dn492HMT2RpEHVB3sks/veaGVVTyvRxHJ8RobUVy6
hUk1PzhLDjZ4k0GEkLyNyAGkOBpFqWd+h4Qb7vqJVa1IMTynWP+X3gsdmoJpwcW6
YvpNls8zl/no78M11EOpk7Eg2YIE2HsymK5SCk3rWIMU3b6zYD8YpBGqh5/LTeSS
2Vy7IrCmtWVJajN1QQp+bzzd0HSmrLjWT73O1TYh9g2kp2pBFmBM3riP1DY1mDFB
2af19x3/3jlAAAwHztLXgAOhlp8uUSZ2is9phVC6O5DHm8C/xx/98vZFoYzKXbsc
5gdgsD1NAu/YTRZ9ZezdHgaCjBbT3oc8eG+6GzLmwbXGO5Ya6iFA3FrpJcjOz1xa
a+0dwEalwkYtw3+rbUBklnKiRYSg38cYHVKB6V0ZJpV7+F8VkQC1qtArtTEVUYWY
FoK/+UqVR6juwhb9B2NHUF038j0/dx1HU7XheZ1jtk0jG9VlljoFT9RO7DD3InlU
JAZsdcA8sgKNKxdlChuq6Lp7hC7UpybrjQLXgS/LbdNoET/klTtSGQEtznU4Gy4A
inKRGT1tEUK84OEsuU00IHbA1iWQFfuqU+3ScDxCl2YKucwrMqj9kf5KG4qMMrVH
W31jseozNFus9oihLmhuYGQHPxOFMGnNAuWbEd59smjjgMqM/2JgRWYVdyHsUrVt
fydsDIPZb74Jux8FQR/aJk2nj95sBb9Bo+6uDvjeGxzrNmuWVpJgYF4bExGrhNAX
DQ5TJbEZ3kLkIuD+tT+2YxzRh0g384gJQqlcRBHRr0Ed6SYvHmQHLu3xpx/h0KCv
Ha+FOW70KEbhFYZexjiBeT2bztqpOAcG+YAQ4fsaOEGM3wR17Idjtm/usB6yKxCq
4QQi11uKCRjdMaAeraIaa/aOrD+4XgbR42+6glZ4AssXl5qzjRnNYsRgkvhMDcuC
x9pIzngjwesv35IYqcSrxQs7ZfUJ5BHUFOS4r9aDzwmdVBhAnsUP9JBTjLqShcJV
YDv+OJEmGy+Rzath+1DxWFUIR/RHFgsJEywzRVYmbtUDn/2RQo4qJHnVgUeiu9nN
VwxL8K04YUOL+FLSny7ZirelMPxi/7BYc6mP6kgA0n1TmwBBV1UTT15PY7Y7YPTP
R993TKdJgmSL6EVH/Hk1QOUmDCrFKjBRCt0U/oJ9j4bCe/O7eFDlLaDDAbBiuq0W
KX0ITZsOhIqc5H3Lmchitp3xk9eNEtYl9pqbew7vv6hAGJOUyHJlpEHulgrShebU
cpn2Aywy5ptPchCWhAM20vq5G9r2d4mEFknjsqQAdwPjZAqOSrVWjgZDdscwq3tZ
2aHQiGoJ/LeMwzGMhqdls8wL9wm/2Ccbk2NX2RNA7ruNiYxV77O94hDQiptGEOdT
ex8WIe13q4yx5QFf56X0vt5fYjQQ3/lsEkKOKhyWoS0e7h/Vh8+fq8wu4p7+SCi6
LGqzWnvlKmnpWdXST7xHKF8QNbxdHsYCjrSXlo2zzRLrLwT6JfeGmt8xCwK+9IQF
a/efaWSDZbYKW8l6ldL20q6p4D7ceBjigCacyEgnNLC6PssXYwTeyyJyG9Y+nqHb
XYKOziiW49fxSkjn3GFNvZPNZLaKQRTH8iWHQOMkexOFpj0ImkvEjtRU8VcF1JEA
udELj4nCOz2KSwJygSbzZl2xj8szKaSll/rtWZR/m9e39Jtph0YyO3aROg/ZnUe5
mg6HwuyR+SBkI/+2BiNgPMey+Q2MthEUlA6/pSNNEjF9FOZNf19WwfQhkrcXEMGY
nXv+TGjPFyL5NjVwF7yJmzaMt6+LBD7QHvyyQHU+1QNCLxGJrTST9T7/EPHD/TEM
MPNiB9IzBTSW1j2GvysRlc2fwGZKsScDkPhzewarrhlaTbxN4fgIV1/Xo67dz/Ji
+WY/8ktnnVFpmO29OaWiPHckeuPdE+swhv4Utt7Qv3hEXL3nrwAeOy4gGYGr4qVq
iEDa2yNYDd+fG4SZAA7o/7eA+g7vE7Y1hISwyvGVzKy2ALJxHu96AJWIdhtoHHN5
7I1QgSgI2j3DbHwUmSpe+PuHgU0NtslrcmmNeUSKkLgjlh3ue8BsU5SdbAWM0ZWb
s5EbgEOwwL5yr6JJpw6aPECIkaE63LyQoP0qXUboChkASeOrS3nWiUx8Gm9bnFmf
q0WOYs2j/ECqNc1bQuCHDVjeAZqzcRL7uHui+Xw5LNMCWFfURs4C7saYdaDounKd
5jCq5bq2edMz0WsPxqJgBf/D7DohH5qLPFOthd9rIkqqI52PR6xZHEGS0yPAu0kQ
o0UlweuKvDn2emVbLwbFt3tB0c9BD8TWgY3ZqeWn1ndj1XJ0oyXaxR8HKGUWjRql
v9ORIjWhvCaClFSmG1PwfCrhFnbOcLSA2iCbd+56+UuKYkRd7n5A9rIMjiU4R0Sr
ADCXnzcDUa8weQfgfYFd6Eg4pFg1rwaRXJc1qIi9G4trduZDeXrpmFjCOdESRrEk
nn/RA82VLkbWqP2byi9vA3CuHJBiV8Yf55CoP19F/8Cwvuf2Ou3YG0wGW1DSjfdD
nWbpVzPel6NUbNu6mBfxMRV7GBP4zaXXcPq3m8LCQki9MRerdZwlT3EPDHjfA7OT
wqPZOOlTuAtheNmmZYYozWHsmsWk3mzeis7jtZqc2IAyE+E9oDSDomqQGGLmobvu
kksTjDCthQLi/UUEVLIafQoQ43DZ7iWQykRCZ4JUaEIEr+B3dJ9OwfERNeD57SGC
5wXuwIKvT1GVnC0ugiJikPS5oQdpmn5o5zGOx2iZKn6GuT32XXlSav6A4aF7vmLJ
5XzAcDFWuDB8XI0RrSZ9Xz90jxOyKiJLfvoPWMX/hOqT4nnjSHyG5VpqeqoED/hI
X9a8YF/Jw0parDC5gknyr6maLBtt2+CcMPv1ybpUOBMiTuGU0UC7UZCDdi68xUoi
N1jMGBM3GkQbwtU/pqazYs8iO/H7MSbIJiOZi+tSOdK2/706/yRPen1mz1gguE4n
L+qDDDYhq4YeIFSWjimC5Q+PFmrAz3MmrgUD2++lxo6v+YsdhsAlipINtAKNixJg
nOef4yGKnw5ZgK0E2gmODV5DGC6vY1hdR94iOUSzyxhpVaXhL+aZETutcqkaE8wp
0prxc/hIh3ZOgvIs7wRSdLqG0Ec2KjfCwt69IqRTIFSKOu++ox2vPGI7rqIN/M0T
r+6/CkSfnCWUEmofZftlIu/4SeVKU7BxqoDcLOR+CVqMu3dN9SdZKsRv5+fqlMMh
hVxeNdB6Y0B9Ms+Y6IJm1kF8iK63V4Fxiakj4t5QNw4yIBAVgbM14Q/iWLaOArAI
LDkQ1WPam3zszDHuP8t4rNITY+17DCs7JOdBuN6EtgDiDcy4wWu3bboSir7GJwtO
N07nX39D+r32fy5oINsU0LNueAXSiSFrdJ2JV/0PuJcqjVC1kDyd5g8VuFddCb27
w/SN9mbQfpaQDKfZIo2+5jll/7gvEhvxNCfMdbquV39VLkaWnT5A+iEpuiXlcelB
GTvJVwcgspwmJ2kEN/VFm8hcrUG+GdC78UGXP7Ypx04f8afgJRhMKklT2uODt+FI
+D8tp62AMO2Wy1htoF3FvUm/g9UnC4r2KIItrJWm8icCbEBUlIwIObSeSizo3O7l
Rz4x3nTAhFxhOaDmoU88Tfr75KUuVAaXDCeF7ZjkIOQh7rxEO4jCwctzt5happAL
mheSivZmPfxq0XIEpjv4mrECs2rb2uRy+fT+o9wOd7Z5By2qXmf3gxGRhLOcoja+
IdoRFfce2zPQzrAyzzMDZn2u1xVRHO9biYbhAsq0hZQlIXgpU2B1aLSm4XAOOcrd
4OqnpyNPvvN07z8r8IT7C7MkFAhY9WBaE8gbanGeopPv3+J4rHj52FAtaUD8we6/
t73fSIByHBr8pV45tgVzFcRt1y5X5bAn+RbmXo+GzcIXZkZalruE6Kf8aXI9FxSx
t5SzyQMBWSqpHCWb7QQSkx6xLD3Bwh3tToJgxCU9CX2bcODReA6k3e0d6n9TgNB8
/Fbt9MVDuqOIfJeLuQB3orVc6jHhX7lLbL16bH/LTtj1YixD+zuifMquw29vA2/+
M5lh4fl9GaYEqBh+XV1P1lAdkbGoYnSQtVUFMolDPeAf+jbKNt2QhpYDwTL0uGFb
AZxb5AJ8h6xoycQ1Ta83EyzRqGW9f3e4LxZPf2Z8lpUF9srOFFvGHiU8ZFf0/2jj
9chizc0CbbJNd7ii6Dj7PxDT001G6Y0wMApEIIVlrhhmDb8s2PvC5lAPLflah1aG
1ta0l9xrx8u1hVPuSZAfVZWGm/2Ot6o/2OmGZrWGQoppUCTS6SebKWzNYW/3T7Zs
aKdcHawCQ2ZyosuuZIpJLvB3i041pH8EOkLEi8g6XvrMmhgPNtSfaujHdbre+18h
WJy3gNV5xdWHqpIE0JkbwLtBbb9nxVNjm88orbf1IAQPOwYXtnUCrdRrK1WaVjeh
Rj43M2mXzFWr8AgpLZ/LAD8WmtDgLWC9n6KTMCcIXAfR+SlfvVo5VD/E5DQyjAQ4
SQ3h4A9wr9aeFMF2UTfZCdOu0Hejm9XvhKp+eJ5EH1V2tkU8JU9F5k581acK+rLR
8iQs41z+ueeQ7pCn6OD82ESZs+ZDatvyioh5ucjqqT7ilVVQXJmjoNz1XKHdxhKq
QoFXaVDPCH69bMgoQavxmZuQZ9BFJ35WazoESN3fxZ8GMz2f+idaQBc1NTTfiAx6
kQoYyC4QsqSuHtDcgMc/+11hHQaxYf2Yv4vSZso8NxIvKldfc1G5iJsoicxE9T1k
n/8qabPTfHP78C9Rd1l6PK/qGDrzS9D74mPJdrPwt84Y9cARBFw/1ILSkq94xFr3
zlEa6V/5g9C0Hbe1V9YMbsqSqCzysVt+2w9RdBp5xCVdjch6bxK0k43uiBh5iz54
kGzmSNprcfqTvUWvjLMe5OwwqQRKzdvD+6KhduCXSo+ywVdzbP357xNEm6AsDI7O
DMM+PTzSs0HdHmaNp2tlgdONJD0UWtL9T7DfRjGNAEzvB28070Dk0Ige2NYFbHxi
SPGx/HGWxHi+ukt2ZIKN9voJ61VWDjg5dLwFNSO2j/33o5byRFiGlmHmJfX2W9Uu
lnH3456S6+L2gWTZXnE4qriDLEmbNjiNipPsVAbHlcGRsIxGJa/RgmIw494np8vH
JIEuZuyyhZcASZz5cseWlfS+TArskix2Y09P3L/wcCPtQJThLUkPaGW0XPAEofRp
1QlaKMdOC0bEOgo88St+WMJxjcGtuHlYHCoSq55oreRKCqVxxWceNJjwsEeoU1zY
5JhkPZit6jQKQzEhcSVfIUUeAGZSHxAEbfhYfvLtEBiQg2sXV0G2FF/j7q4QBrvx
mXNVwhqo5IoKE6aYo2AL8vmHfBRb7K9LYyoO8xZR0VFtRqcnFnYN0qjJVpA9FBYI
I0FEn3KV8Ds9nBIPA0jqklmLcQmc0NlSgwmN1Ui/F6+CwmhLWD7OI3lh6Rhstz3D
/sLLIuh5qCuNDclI5u8Zx03DWdmkbmFSux6ffeev/o5la3QvMnCL8/NCy7IZ8fTm
og1+K0ANaMhGIdpOHrCGi8hGmUXZQ4U/5LGValpPzG8+YC1ETnkpeLhdMn2bByZc
lm3T3iIzYYlTOQPP7pWtqtAQTSnz13nPX+bHsq+OZN8naFsiUfzOrwCxLiA3tr53
IcGS3U5tZmcYFWPI/V5zwLR1PsH7wZbNEXtBB45QOjddqWIXBe02SzzkPYmqomCB
ggbVkN1yoVnv/Ojui7GtYVPVT2d/fgIi9j0gtjEv7Stw5sltvwcqwtVpiLkrc+Wk
O5fln/fjeKpiP/bwjfI9IY+9t6sQ2a4Yoqd1xRPJ4bbRLUfXtbPFjwnS40S7J7xX
cygDQkt5XZYG+sHNjBVCyHCU0G2KeRFPxvcMN4/g+KW6PbZo8dY9vuGao7ixlKIQ
piJXCpfNLUST91d3gDxvRFRLxpI4rRkuDt0nOu4Z2xcLjDfLwftZDvUxsmOobslM
v9AXvl384exgsoTD6ZsdFgjFJNeMEKfmSfuMdTFdlLSUPxGC+DS9lh6iHCknTja7
bu4suDvbovqLGqvm1aKXLm0m/H986lH8wHoLDoMJ/l3cYBCuDx9e05xVlidTeY7E
ULQ7cDVPiy9rp774vi0fbf9WxDv2QGjq1GRmBTa3sNuMA01kUTAo3lDZtl5MVyvD
q4X+vbbCpnwhZZeSDAqhl9wCLnGt6oBJDakswzuSGZKxwqoSs7cO4Q0xR2kG5x88
HqHwpImx7yfrmc+SUKR7OClD49Tv3yKgVCVmjfIKocPNkQqu42a7COqqH73+5Nyl
jRNRop7ja3jAzouWdf7L3Fs2QvX0px7Hf2X2s4ii7IKn1Yf6T1gfXTLaDtiy21SK
NrYl3nInp93Uy3hOWQd2Jj7AJy1HjeyhdEi5T37f0TQxsyWi3v2QGfasVXz3xDNo
p3A4rBGNzQrV72xwOOhunjFVlIZv8Fdb3RMbRBTfDnLoSWHAQg0MnzlP4tsS9vw3
dV7i+ZlNMBboebZIE4YzUt46ojeudqIGrIAptF6h+KauUVNAcFGsAARdl3fIJYPT
I8eZk3XctMwExqKRvfi50JQjRXmnCEQDsUKyBQ/YDRSDruScstVzQ0samoEz8yc+
PWnVJbJ59faeJjEHwJpqCW5dGrSNYiHL4+dag2skDFj2mVOgEWlyGKjzcZK7jpvN
/B8i35aw3//PsawlDFmu1h6S9g+I2T381QHNpwu2LzJ0yxUXFYXCfi3E3nQv4KXF
H2YSXG7QisJ1nDYcEdOCPL67+06tFX5X+6IQzxlK3PgyIsOoMmB/hOW8oBZXAWHa
7lNq5nRiqWHV3iyUOhTKP5krQifS3cyoMgEzKajClJ6BonHktj+Wg3C5KV8Vwq26
PbWz0BDm8Gx9xZwIY1WboAYOT1KIvpIrrvtbg3ICuxGp8Ako4C9aAKL7M7/7g+3Y
2ERJl+bc+cJET9z2R030jSkc/sfcxWZa/0Y4udtPH4QhtdXpSgkp6vqYrZ+jdaCm
bZ86ugKrAdo4p62/ZoUZcjx5MXhlcq7PkLw3xsOgq71Kkay+5S+b3Cb72Q7HveKh
BRW3GuHdboTAFzcGbMYxV1UHa1ozhQIli/975TiTvpge85sJ+AG8drC2euOkxvuP
Xa6905GfaaUsTDPVJQM8JG4+qJbyqRiCJqNBiIjZKuyhWezObKabK29zkwX/MC5x
kvyvhxH7KPxmVJI0E7eGvXOrWvDmDPqqR5n0/UCN+zZktckb4d0OAo89eJwc1mBK
EtPRa6DgUTbe/6TF9YWgOZyFjfK9nJnbofx9WUoS5qZsshpzwHcEl0tS87TRkKfE
F2dLBXUXeKoKwYoO4P8j0WxVJJZKSyIj8jFv64wuf2SRZz5HyZEpMmxjllOGKDt1
HJ9uY8hjXbOf7rhd4xcZAD3PXXj8Tgur0zbVrzPT5W5ZVX/lffX9w1dDui1F5ytW
rRjPN6je8puE8gXUkOwyci29YcuDmgSrJJ5+KZmkoFeoyGgoGae5no3u8MsSq8fn
rwvVrcdC9bvFmcrSy8NZ7r//fjQUG6pbGlmY4LGea+MFd+KPNaoIb3bFeGUdYW06
9LTwjfHxpU6hrgLBfPwM6WF6U3vQc9sHu2ta3DeU1mRvmh+hXD/x6pCmnP9vqHHp
V6JAP5mchedj2sBliNZhFl2MBo55EClh1l3niTWu2Ie8tI5YpAXgXbqhRRnz7J9/
0IJjl+Huo4uBFLCu168vTv0FhXs8630cC4soOWjFimu/MkDsTT9uS4+LbqogTUr7
wZTHHaPwCMeVnophd277I99B/70lalP2VpyU4ZXZlC6LYat95I3L4rDz+fxLD1HX
4j4QEt1/iwFsFbf9UhBTQ5DPIYfLMFkpVYes/AQBS1wCSQEZAzYg3cHfw2PuKE8S
f2febRYJpvjlLkkNSkRqa+3mV1UzSoFpoqkFJKCN2MOBpA6/VMF4DNDXocmkPsyf
f9ciuF7/uK6XE3ZTKFTrvBpO/IGk4QHQthltnVzA48mnh4UXC+U/M8BiqbC+derx
ChE6aSJ6pA30YGVhaV4CbIjsM8IP3JRNd+arW7HJIiyM755mRw87uFaY4JotumU+
hLW1GEItGkxx7YZs2MLFRDaoW8zM1yJaBEP9FIkRE6nWo2JVY3lh6yVIXpnPW/UP
3vLoZ/vUDtAwd/bHL7OOhI+zCjB/Y/mQmsdqWKbXyl1tVK9HRwCj8RaSQF1lc5be
Ef5kgRTRSsiUH/tWKdc80O8f3NbVOI1TUUx0f9flStTzQMvbHMsUAWHTCZjfvwIb
P1ilTzqSRP9+nUmBUcR66Fa4F6RtUAZPKeWnq8Dsnw9tK12z4MR1GR2vtYvdDByr
Uv02jXQx58pypDNWzAxWQrv0DibGsfX5vL4xqOE7dXbjCNxqqj5lM0Tu3SoTR4In
gG1Um8dbAS8SS+TEVapzxLz4iHy0rtzFziGC9KM3Irsbbjnu7tdCK2TJ9XLwbPxF
mz9T9R4+ucGI19Ll74cTeXLXjm5Zg7p4GxPLkLQi5XdhWJ9/EHYjJtkNOsENuMbk
MoeKHcTzGPSoGWKvqDaG1ORS4fIZmzDRXwb3OnrJs0pb9sHThiZ8UfYW3uyk7vZk
yFb2IxNNsmn6fEu192f33pLul9kuuv/qjsax10DJhkQ0QUz01EOtOY7EOR7rYhRH
qdU9G1et1UNAadByEGC92XLqzN9jsk8KJm6zgXPVQ/L2sdXd3GyyHjh0pIsR0LnB
n4KHRMI1SgbfHKpmY9ApHMw7dNWkCa8+s1SxA7oG00jcmGq8ZHz1lZNRDth1QA7D
7n+66D0JFeDbpxpMMNnEpikAwg7sEbfgHT0BNhh7w4MEbD25XVQ/JnpHuNNrmO3f
Rh+Dp2m1M3oqO62oXUzfzYSKI5X/jHl8jMZMJC8pGhgqWcVt+Xd+CC3DjpB9ZNut
nThMIIJDYC6ba5gi51aPUX3myjoEVZvOeML8hDzQf8NdhkSMSibCggOGgcUDo8dq
bclseDdDhoxaESWQRjavFny1nOCGWtd3iJebATvQSTl2TxpOxH9/BtjS/swUmPn0
LuYJpFkFndNA6LlKZBvtwZ/OGOC9Z7XYzFSl4CIsg9rzxNYcVizQW3+5kvB7dPnc
TYWYgQZLwWuWKV/tXjprZjKnZhHAz1dW+EjLDttq/gkh+F1q40uNSTuutKf6qK3j
rqeV0EwOxHfHYrEuwZDEtg61pZ64bVpjtCIci5JyiynVyiGnsojzP4PGWxTwVgjs
NBtEZHfPAUmFdEiaxYWwheJfH/DsdB9/61rFYFggclpV68AmDxXuyFFlqHeKyURe
ER29h4BycqENC/8KA1LCytfm0FpxcHrHOmroAT13gju1wFkaShHut2w1a0lrWEtN
irNRtlyGIlH9l8jFlRnsqvPWeYk/DNYKkt4Mu4NuteWOOvAaVV29+obxYth1CN0j
mMUnz/syA+tNJCWGNcksiWtvsqKozmPin/WBkIhKYq2UVvVgmsPppRJgYvZx1llG
5b07b3d9t+E9H3zvGeIXAlj+1wFLmVaw2MnROM/RWkJoYfXJoSpH0Ldfde66KHiY
hYLxEDMW4sOx5vEr0UWvIBtVfONXlVVLseNUJN9Q1H8DE1xHgqEQ4NqFeVU0azPO
tjyYkP4wMBumrp/9QW3MkeIziXArtVzwfLrx1hW2FOYGHbVXH8IL7+vjQD+eGW9J
xgqdjQsnD/AjjlNNr8SJG/fJtNaut96yVB5J+c7hm50Lai0A+/I5zkeFSsqxs8vc
dGDyvB5FyG1J0GKBOF7CfgDzJ2OFKGtK0WcUcI+Cb/H3svKvSProdyiEzJnRR9fx
L3yK6wyNjAkAiCRMv/8G5WKXP82FbtIZZNdgejtI2kRnRi6EOh2LzeiYw6hDoGTW
dUgK+lb1h4M5B9oEKBf0saDM0/nieOWJBaJIwUvBwVqJ1g13WwtrPlRYCRBDkSPq
cGu8d5gUdNk8CkrSrhS6duwtVUWKJaKwtEKernqnteR7dnfZDqxdcOhdzKv5egjy
KT6372Z/AscZFl/JTZJ/Qwtnwo9YqqSWq/a7YmzRVcvx9qp6iEC41N0G1X/SgpjD
GSxJxTJSiIbBmxEECdtcoablB7UAYUdVNMS+8wcXX1CbrwSaHiEl5bhzgDHRiIWf
Qle63W2cT992FUbt0OB8cstr5m4+Uoixb+vOphCdOi9N8kNI0HYpYoR55dkKmaSc
TLpL/gxSr42fCcKz7jhA2/1fcYwhCMTdFnO58wX0F9AMem5F+klRFvAGJxKRKTkJ
cqQlwKSIu+Ns79MTxuUa/Cp0iaGsPqKO0w3CYxSNWZUzDpEBCDydy6qDvfif+8+9
FsRGoI/nBnJEh8DjcM039ty8PEesoIMJ80DmjqCojlZ//bKPrap8R79QnrKoTPUX
meRS2ZP77lp5j1rfYeMkB27n3nDzJ6jwA105Xl+mHXYTKI8/vLVD8pdnKCVL8t5A
eVimoBM+PymE6GSi5mlHbhH8xfRpaE6v5oUz+L7nh1WA5eaWJ32iD3kzmXoYaxwJ
RPzgGIPnSK2P4vYnzC9IPtrmxuR3mNRt+OzTtrRxfbpM3ITErB9zD8fZoqs7IXxg
2uuKJsm9cdUZo5foVJchv6r/YRiqFROxCB59WsLTVa7rM8FJG2yjsQ1gpv1G+vLY
PrvPKHugQCemhuaTqFDcmRgo4JOcjHetwcsL7rSYrflNRqxk3WPWzpjvB707kSsf
mVnUe1hJBkTImhWf2qBer+8vmXYhXOTrIvYG9I+Dx8Zbwvr7n5tdEurHHivCkv0q
g6hlDQjURqtqAedHAnwLTOPO+HN0NuzxlhxiifOJKcYugdFpqYUPRZ1MBTFX9C+p
QSrmjz47CQ+AORuSwF4nXrMCfw0UZo35nPi6cArpz9UYTrdHN6qCuRsmZjgm2/VW
ImXpyGqG7Th36f1aLmDlhWundp35EAWzhRylnlopTFSJEqUaKuoUMGSu7SmOdkkz
Clk39vSiEgR5lWNpsOzRFD/0pnbmY13JHGat9ghiOani/Gy3t5ue5wj6Vo51NXDJ
3QmvfxXOqEy3KLySP177oL4ZXdya8taPAEeJeHQRatWMCX7BRvg0h5HfVUL3pLmH
b/Yeohkaw3aKVPk8RMA7fNKK3766sfCd2a8/xHrpSLIGFPEVq9K9+51A8xMFQWJj
jKWXNxagKL1RlTN86x8XVHLLjcCP7yL3V1FEsFb9ZZ8Lf3g8bGm3XAebrzsZr9Kr
HWauNzfKmE1Ya0G5UR9Ft/qPVtFjvKWNRjybqFwWNINvarugKZ7akszKTcdWSQqs
zMLDUCkY8c/bJXWEUIloqyrfaRwdMZ2aFLvxRMNTkdJSPhC/JG/3c5/Illj7LjrI
JZBxDgxp+J4gTwLSGVSCjuv0kJdHd+XncaCC7XHBe1NN7v98qiN3yALzWur9Z7cJ
pNB000kHqcAW4h/qV4SSM5n44XfMVxasrshUBFdoHIZaps8AQq6YIepO3Pu0eHno
boJi3DHFYGG/iBXkTtbHwSvDA+CFnZFD6jED9q0VaPLzeJbmHy2dFJ9CT5h0B5Id
8y1O22I+t/GB+fqezAQ5NTCINpzNEkA40UtJZcT7Mhml7RKgPX1MP6UoI2k1ju9S
DVlVlB7b0rspMwjYeGZLYNBA4ilJHJJ+lRmE1AQWz+1IBBNcM5jCh5SibmFBBFyN
Tv0AdRsmFC9txItWGOtv40j5IDt3fVKYT26v3pbi9oY8QTowCK4aLcUs64dX48Gs
ci1933IJX59M2pr7jxd3mN36mAUhHy5vIH2gRhw7Z70z0LHGI3BOLVE0iocjumgO
xiuPQMFZlGTy11BWn+4pfQ6ZlIr4DmopAL440BFl6F1kwfkKN8RNZFH/Fu0uOl9q
Jb6zP/0ZaXJnYd7Pq6Ad29dCPZ/KbtC5Zc8gW9GSEhRRhqZ/KAnlRybGQzBpSDqT
ZH2NiGwjk8G91UVPkhxLekO69AYmv4ocg48L4l3z419+uvopP0c4kUzthrwg+0Eq
D1SmrX5iyOIydQXNl1W+cDQD7PcgbLdhThIthzOSBYJZXZ2xfy7OKrAOIZSaD44D
fgmPDMz7l6B1STvX9fjaQnsPwQXTh5yA5G0vKm/n1aLChODXW3R5eltBb6/fEQDu
/IwBsTtgRF0IIfPptS9ZQzlbxIRDPRrITVtNCkG1alaRKf6+MBq0CyuwiEOQDVKb
BwN83PV24RdblRH+gqL7Eo/ozAggZ5JkOcSNaerztrLJDkk2cgjy7+FZIN+jeRWo
PlUASJznavqdxfUxFWkVW9THpt9YfpE5gB3J/O9OJI5SYJreKdgaX/1fE5qYo54s
Q7b6K1AaC8ewq428te22DPbxQf0KLQ8AVGrmdiGqLDWGHt2ZhVRIF3+cks46G/tC
0C4/6UFvyUactZVNAIGtEMFu1XDPZQoQ8dzVtZG4MU/t4BcIhpRuRoMGgNKoqxFP
1QOkYz1ix/FxgRKBpsVTI8sqqEYZn3q0P1quKMBeYtH7cfGY4xuxKFHsPEXLG5Ce
tolYXWLdYjju+EaYgBo1NruJBnIC6IOY+Bl2YRy7N1rV5Zq7JfI8sG/5gadZhytd
DThMA47DB/90o53dGapseumogAT7vbnqXDE8UQoLnmEGEq1ZR9HecK1mEGG9BZUF
nG2wl2+jzaCuVo3cRNCOPnUdLjLiyLNiTLKoRcw+LLUw52KpxCgnjOOc+V9ZempQ
lDoFEKn3cop2goFoOWpq1VYC8yo0CoWjdm6H44Fe9yb30drEemrp9Yh3hKxJd/JZ
0cuEBJPTYyuvWnh7lhJyOuQ7UslTK5JXOlAh7SgviiwW4vJ0Lr/VJE1KqgI3ydvO
pcE9tGSlCRdmFjpOYhGgCPKmbaB+Z9EXb6MdeK8DVegSA69HYxgubwl5eAzYX+bo
FK4x6e7PnA6mn++OhkI6C5bIJnj2L0ehPA4xJqk3Up2/YmNv4m78E3ygRUftV+AU
81xnlNaFUl+JvHMyPsLpQLq5hP1dEshoeboQWX8CqLHnBCr8G4rYnBJ7hDIEgZRJ
SoRR0k37UG2O2Edb7eUGxMu4l2HSgZ/fHehPfWOUO/FTSXpYcu9bKZfY/JVtBN+D
Txq3pdh9rzMXEqpFO3QfecUZPS00zGhi1on7dPbGA4r3WBJHvWxI8XcQq0eIygar
UpZgdevRYNdcHTNyfjh5VUZq45WGjW3CiueLusuoLVQGrGydO1EdM3nSsZrTAol2
hiRnWOyh4iVSXCg2VCorQpUv6tWDVYez3S9efzX/U+PrATjdu5fW8vnTbibFQoOV
3DEOy0xFKulbKLKC+H21exZcb0nkLMgFLxKvCN9QThw6Q1S7IxhGzs0Q+jwZ9tJ2
6wOwu/3cIT5iWPYizPRBZ5RwyeX2nCREFaQQayP9+YMINuRVR63ST0+fdcnFVkqH
0g0XUc8GmL5yk71ri6WoeMeY+qdyX4g8CKhtDl2SvfG272wq7X1nddUDl+TkWYuN
CdlUN8Uk2CqJtPwZIu96vLqW/iYF9qMbTMQybDy1JokrzREkCqHIqpk2YcMh9eed
Z282F2+Y+nRlPgPx/qYJRLJ4UZ4eNVQTS8Pr3Bk3JSlgKtPyuB7IKaLJiU6F0Sdm
0XXLMSD77crn6uoR+TT6o525vrdFEmlTwRJt+NEUDwnCn1MdfOpdBtoDg1Mklb3g
VUHyrdTnUoTtN2A76QQ/HvLGXzfj92tOc94ZDIwDOh75JdAgI5dCSXuLSTIR7PBh
WZJv5O7l3p7u+9yKWiVDrEw9rJ7Yf8nyfCTFoBpCj6gR/P3f4dgwrFRDO65Uhli+
R0yc1dHhQ6qGOOBoBWcNK2ZEUmotkkJ8AKAbtueqYtx55FQqZZ+74eIPdhGagWET
iH4PC2+dbgVFymcWiWqyLrVIYtG+wMUfMTVRWC32sqtFr673X17iJU36s1wntZXa
oG/aLZ/tXu7wJYWwXsLhlBk1RYaiQ8loQ3AeRaP+LVZk9ZXxgSgIuAYEf0I8EUKa
oschyE3+L43zqdcTuywGrpCs5G0T1M4ygO+GaDDutdPRSY8l64FcJh4/cPoF5Chg
Fuy/TRJpM8/b9nOYZPhqnmyw0ws0hu6bzgik1h65sEP7/WtlAnCTtEoBEK11+FPz
1GLGHbh7QXH+p9KLUW6sc4OCOdkQFnJ0TbA7M+YRT5LQvQ0DEs7FkZofYE/U7Pdc
9MxzWCklN+uZ6BwSroN10AsqlVKB8Quh63N+SmNxo31zdvAytPirFCcIyHUVZF4b
zzZdJOoGIwC/UVEoBT97VXQiDL81S7rYHZRQPkbwotyTUpyOH6vQRyIuxWeVoDvB
9603QGho8FTh2Ebcxw8oDJHCIyo8kpQ/CQvfBI57wsOTQ1ciZ+ygmQ0rKAEhYh/v
ijkRryMFt8dgdV6zJQcsb8DsP/rwwsp9ExuMbiEJtXeN+3Z0xMsYX+Q/GogkuwDO
99PJurTbAJbWw4M64pjCBWsn0G9vFkTtZguluh0w2G5/996aS3StlNp0ux70O41t
4A93lVkYZKEXLEqBdmGl15yttYqCmIiEwEUrXBh4mAKx1s7ZQ8vvp7Xd4eP8RkXc
uYpjQzhKPul34/Q2bJImrV+tMflflkmovJ7vj2vK3dr6unWyJcd6OTDefxlBhEXV
jI3ixiyPxiPxmRR6ZLHWSPcMLTu8RzlW9XYmQ5QX3VHNmkW9cC2Gs+K5ZGiTHg7K
vsIrjuqFt8pIBigsUVsyZacjVtI/dstz8R2HlmsdsZ1y7F+5y7EC4cJmtMiZsYO5
K2L9/YkNtUD8siP7d75JfLzEZ87T12Hmzfz8Uq5msRX+pHEXnhXEy25td2RZovI3
TXa0rhhrZMt1WSxMi0BqmiKQUdPk76elHzYTPIT2uqntVR078DO7tl6TlEos536R
WkqNN58AmYd2T+fgQbBy2LAyH2qXo10B6PNzDDVas3YntI7HyDQoANUI8dkwqZ85
aV8rzu6mR0thMRSFvCHpeyCmd+7vWt4bU9ypYVw09J9oLE0X2UR95HawRY4GEB8U
qz5DijihMF06g7CZ+RScvgZApjh7z9WiJGtzuodTQeK8N2cGag1QpKwc0N5hiAey
kPMgdro/61ZoizDdEceigncDkZXhDAa0vV5sj+zVQN+Tu01rbv/uN76i6w9tXRDF
8orbtpFTN0FiYHCPOHbgjJaJlfo33+1jCi3+kiKTf9K7ln5cbY8AVuITr26HdGjb
GYnAJ1q6dJ1aacd+VFckV+92fnd8THXE/4Kt/VdpUQ0KMH9YEq6mq4Sw2yD3UGPN
WO6+9ya26jUc31k97Dt2z/8GSvYh4/oxDP/UAHGt4CIIkkNgFG1GA5QYNOGSkgka
HdM7W6WCXjYmiJG2r2DXr7al8aZ+nrV3A0LDKZc1OU2fwDXfGAnuNc6Ti6l849j+
t8Gj/rnLnKEbdIyzwxaBezqZgDVxoozyT3xqjF9wvuo/5viKl+a1AobatxeYVSH6
igTp/YPeLWamXdbTD0yLoAV4w/jAUeQ5CAJeZ/ADwRnWeTBTMeA7x3dwQEBa1h+F
OhaFRlOZ5M1mBhAwc9Eu+54Fm9NAmtrAW5qvGI7ygN0pco3VdPHZJ+RVW0HKcxYL
jc5bh6im/n4Q6nP7SrmRtepC/KCjtQyTbRs3Ruq4xMBGW3UEVAUtVywbtUbHaE7Z
kOme+ClcnKOmkv2kBdo7Jtg216v+GKaQArUoKRJiK5DOIKo3mSMaEAumqSi8exWI
CqXMZrkTMDoIC4pWNJIPeLecFozBZB+RmFkE5rlE9vlDI8SbyQPtoy5dRMMSguFB
hraBA1W3Ryae7uS9LaKvBzPGB4sxHOrr2Q3EbTQJKa7RODGiYb2OZkg4Ov4xlT07
aujei8Ka1lHXBksryS4n9yX6XdIMWJR6P6OrN+CcsB4tVLEM9D9nuILKdOu8KeSK
WKkfff9WYBsSEt2PjwD1hRJ6PNknFTPwYM+DPylo2c33Og8ZbgUmo3kSEKznG3Vj
ih3JL8OqKgXX8JD/HpM+S3Zn9yS7u9eCQfNusUvwL91uFQ4Z/6/JS9KyfI1Jkged
gea4qJgcX79ZneMh1z81XrG6zmZqfwXmgKpvDoPVs5uLeedimexjEvYo8sXQP/Ad
+/fMD1yc5sz98DHZa0f1whDBrdS9QxB9Ja+yWdSpXARsV/Cxl1861XWfiyMawJ2w
W+NUuUOJFHJEMSiau9PAZvfo/hrF3h1H/Wbr+d+0U0/A5ZvVN+PpFxqaAfLL0zAn
0NTnz/Sw2VpcyUaLQZBz4pgdnr0Qdc3sk4KmUMe4HqVzGGbm8HyO7MLPwHqCMxpZ
+n0sOpA1q/yXmHj42TasVWX+a+3KNwyEMRWwb4Thjk/5n4+kueAv099d8Nh4dKyY
FNjj06TZuWp/oiqL9IQtSdcP4St8CeOWz2DR82WMYeO+Tk+0M7X1uYtiO3qdNKa4
FEBePa1yLCbbWbIM3ZCd3X+ZOSYIM3LvITysL5AEnJtGaz7preHQ5Ly9YriW8ItU
I/m7w0PecMP6So+LCJAm7dBTVoQXqzZLSnCnBl1NcG57gVg/Eicy24SVX36mPV1G
ynrsv4jtnuSBoJz3jqc4YXknejK6lGA2CGgPUVaT4HHItTA59a7FWt7e94dO1HeX
BP0H2nPgMLfosD5H/b8+t5qEtS6B/EcR9xaBsPHKSn6Mp/rJp1dpvH9WMo8QScZN
SfrNo/rPIscUPhkErCIH8U2+OLF3oDlaGukqMiGqIhwrhNuDF75NyXvIvjfviLId
3JSGvfAfbOn55AOqusi4dKw8h5LkXOxB824KrPwXxS7NwgqarSa4JJ7VWLiUbrfB
GerIOQ6XJ6bCacKV17JpJb4fo1QgfUfYZZW6RtpotMUeuS4pFHHlPDnqVx9F9SsQ
TV1rVpWFBOYk+AitTK58itfSSEeiVzTNXmC3iM3G8TK7bk6GaF54rtawQY7K1/rD
GDlC75YHjq0NGmQK4noxTTKnRy2PbVzL2Cacyo2d3NMnbrvjn2cPkl/WECl9Qvj8
8HDRtHxTgLuum56LIs9L+F8puSJGnVNRz95yjXeaRQjbnPvBaa+wOBVu57dDuVKx
cyIOeKsvaSs5/GilX0P3lMeNRJr1yM4FXYljNs4X+kMoIotQwtRN+pF6rHxoZnCK
y5rm6wuy/gI6UpOESxS7oSRxLlOk+uJQcDtAdqEDRTREv/9ruz4iZWvK1Q3Gs1SQ
NDTM/TR8+cdk/CHo563o6IwgEnow5FGMaLmFK7X7QAOxbz9JKsWC1SbcrXnEkhfi
I22st9NTdk2q05vxgBorV/vzsBABep4pDqCXI10HY/8EMqUdHgZz4Zu1Z+aNhPSG
Ivx/oyhEzdW1VQ9ob/wulnuYYTIIy5+d2ldMq06OFHs2ZGehiKBWZUhdLrQmO5po
MyW6zRPMXqTXu/6tsC5rINIQP+OQZc0vkIZIB/h3qT0zxSaVL/eXzEQtN5upmXx4
Ql1PK+EQHmqfWFwU7C25/cXx/xws6nJuUtO0xwJBm1JG9+arsjp2shJ71nontpIa
tJQcTVdI59hQEyd5b2rTQXKBIdVRc/a//o4NlwuCcWj4ldlgRPMfhtNS+hF+6BM2
UP4QTU6YV5Pu5l0GT0Ey1hT5EQLtpjn6aliPKrLkYYuYzl7S2S5x+fBy8V1uxUi0
NZ1+Bx2/RG9dc6g9h8fWrtoEqYhk5f+Rrr9i/lHny/GG9qfAGAF4JfUANxurienc
FAXJahFwCikr4RgFMfiRFZnF1Mn01m+TWsWre5ahu4nwbIqDQC9oOpi6aMO8Ri8i
WcTack6wAsDz2Uyc+sj7qUPq8EJA/DV8krWZbvA9pd6zgnxgcGUxBqnoZywTb12g
+XHcjlbQsIvvffVHfnSwjuvvUU86BdTf9gIgsmJ+fjDsZo5aTztdz1DRM2Q5UqVJ
Lx9WzIkKKGxhLP/99j2aVjewDdFwLz+L3EtBZKX9yVxxy2qRu9Zl91Ho59XO0xhV
zl8SKRi2xTIM1zocrOTU40z9dawPvAlDLXJMc0Npp5Qp1/hQnFjqa1DNx1EqLnfm
59GML2+YZBr5maj7pMb3JuXQSkLWn1QQ3aqQmsxTJVcowHG25cIJCXM2jmDsXp1K
+s7LplhJrmor52iV3377iGMYc8ixCTQT5oHzEM0OJLb06lB/Svw+0WDJnKZtBFOy
xgO6cc3MUKszZgoXmOVlW+zP26rvBwMhw/6JZ5+d1XWCKicOzVVqSeWhCc1mnb4E
w2ygl0DA/LIAO80UQMYD0D26Uha19TBpSBReLzLJfBXbYraZ2IJn+y+g8Q3AK3/c
VdALNH+hHuOMO2yh4e6ePgjaGxJhENsa416K8G0l724ks2ljkuBMxoNbaDDQ0nR9
9lcaCBvShV3COje9greVt6YVQTvMxUsN6IiYLSJwZn8KjUpVdmCkM5Rnb5I1u0E6
sJmkCvMuxJ6gHR5+YSBBmPD4FlD+dmradVblnwKug8vqcB1gR4vZ8or8UHe6cYUW
8ItYRuZk6vGCNxbaPoHNZR6+Aa421Mu28gPUn9t+WKTXGE/c1aNCoHTZ1aC1p3VA
o7+1YDrlxT5sGpNi6ZKYTUdM0eOHvdxD62IO7IVLiHpFAx9qkvfveBh8AafK0bj2
PLyCwGc4xkp7Xb2f4Oi3iaZpmsh60fD0Qk4OsyhexPGXmNySFt2TCI7Lso3euA4g
1B0ZcIsjYFBh6xy6xEGT6atYpfD6AIejDH4HRsSFCkGCwOPX8vWxJwnlFp9coMhR
bHr1GZpV3sPI4g4R56ETCgT5kj13iAihiqgkMs7KWaAcrx1uSZcrVbGoZBuMtk8r
mmAz1lW9t9ELdmaMDg+IzpPWEWPoegxByUYQNJuIifcLy4N5O6bB3XYcEnhqAUf1
1aJRCHddqvcd6+EL44Tbnaa0CqYWAFhZIwhBVgBea+Jv+LaBx1PpK6pX0JFsZbZj
ta7vGCva4U4bQ1tYLh51TjhRKtg1XV1vcSyGufTC+8oHlB+b4+S28rQGigH0PEdn
oHO/48FS8oHAX7LzS4W7EqP1sCXatAqa4MICsd+xio9w2jTFlXV+JzMV5D7L7K+a
AjxGdctUB7uzX0eb/AhJIWjDiNeZuMmfdl612lGJiA4QcDqPCjH0MONFhM9efJfu
ze+/awd5EBDg4mrSXJBw0/JdMWvd7OZUlkat6WwoEsu7D2M1ivA5WTgGSxH30KnJ
+feE7R3h2UkSw+kUC2FGeIKdI+YAK9QwQUcJPY7Q0CwSfRJEAFwJ5icQVs14OEcK
pPASb+3Fu/Tqwy9Q7Jm2E7TFd1JPOcqvBVbP89WJs/uD4o157J4k3YzTpgP2vNyM
D+w4paO9UMuyCloLYfkB7Un6lN8fiNqVxA3d+eafrkV3U5KR7gORuBR9s7LN1bhU
kynFxGRis2Wu7pICvN52aX7QL/TkaXmHXW+ryoWlhEKbQySgvoaHo5fzfHJtOu3D
HuOf2ZJMBySKAjWREMhZ1c8zUcMbE8YqM63gp6FiPhcg1j+B3/Ge/wHI/qsJ6sgr
az0LiTL0QMjvv5ORmAPeqw0yGw8xnmxxncRh8k8JX5PYXV5EFGm/lAktxyudNkge
0U5ndmO5LYigoEHulXcdQFF0HuMnEK8abgzwmq5++nPB6KRFT7XqSFN1fcagxHMD
KylfBIbcS6eOhTmKQvdAVNPTpHoX4u6CJonYIk6rXomBR9l114uNT5yiccQbjOS6
kFE2uwXKwset1AjpdoHMm1JbX5cU5FeYH/UJgOrMyErip8EJqg0QtlkRUYUk6r+W
z5JFmgm92xZ8lJkXJR/MpIQd+WBNUASPS5FSfhQWDzI7e08nCmjinasZ9uvntwFH
94lqEUE1TamiP/IV6X5c5/9uhw2tPmx61j8qdFWWOIwJCKH5aDMvn7DD1QNeDVe2
a4OcLxDEatH/MsSOv/C3dCady9sEJISCUwwGl60vHwUn796/OlnW1yyNfmUmG9jo
JCu3C+Ez63gA36/Q+2l4NdkRrqD3wL+bxaKZmqWRjfWXEnMF/PqaQ9oQwbjYE5ju
KUptnUEPZ9oDGtqO8XaznX3Ucdqm1sIPuGtjLG0SWYdhSIXSCcFcLx5DIA0RNTPe
qpX88QT9dubhYd6LGTSemGkENIYtaJlIaTQ0siUgzOsOIMxrigIi5A6l8k1AW4Qh
FaEW5ajeSLwSVqa7LcUC+I1VfAJhMpeHc68coz4m/IlDubruVtgek/6dxR7J96NL
eJtaj75U+MVBPlSUMMyFaGDjD0ri9wPFluBqOYLrV5mqHHk96bzHOI8VBwoMGzTs
Bcq4UwqDWDipF0ugqryxrPT80ZOQfvz1omzz1+ZB4jaazB6s5FNlD6EdMkig8RA7
C7Cpqw8antI5BpY00h0jLYB0flN9S6MgtEBXz9TaL2Y0U6MigLUsEFxc1ffmopsK
yE/KvSH34nZIq1p//qskILXonOh3xpzky5h1m9CUUUs65+BGVIDlALo+lKRLPx8C
d8/7x+noMIMTNxNnaP7OUMa++a0sbfy+y4xTEJ2gSJgdRAgpT9QdT9h/6VTvLtSn
nfh/C0qh0Axh/Acz2+7G6NWU5aY2vRqFM0jKqRMZ79dZRMnflbj+PKiqGbOVVSg5
mLaUl9YadInjBTf13mZ8ZoDwFq7g3WbgbAXEjMsUd6eBdLCpeRcbCVH0hJvTq5y6
4oD+NsUqWQfTj+X9YL3T9OMtPv8i/kSkt1MrvgZXHiWumRF02zQurfVCJMd5mh8y
1gu6IysqQC8MaX7efHnPVIM/6dX4Qvi+oOKVDin4BtHz4/SHnpFALDxGe/Le2F+R
g6L9h0vo2umDOHgYpK0a2D1tohCI2S9Vmnv9ubbQlwpWBfrP/ySJ/zS0waws/hOH
ZVAxaqnMW4Wb8N62lzuOEXGjlflm/amzvKDRCDhL3tuu5ckuF0Kc44MxMeMrFJay
dEgRCrwuXwPnvjh607/7Ys6wkV06dZ1RdkHja3ebI3NaYmC+JJl48BqXbTc6wCIW
aq8MJXihNF/F3sqXPFcogXklWR25pOjPQS3UvuF176aJ3VjhxMtK9eXoby4+CDbq
d2BR5DZAXp6bYa7ErzalorAT8gLcvn7WGxTVmK5WToTmQTO8kvPo+X5BY9VTxejp
3iQapa2pAuet9Ylthg2nuOXk62lKwWsQnjDn4MDkFh1MhwlWmouZyC9Nh0gg8CKt
1mKqPW7HZR8G4LwnBlhmhCpVsSuc2z33YlCA+q3ZFOE/qxZdjIDk5ioOsz4bXSyS
CYtC8zco/sFIN5knBeuYbUMk90UWCusMo79lscPpOUNPs44PaoZf/yot98tU7w5P
FTTFW8IVkpU3W8ybf04yZQ7ojEsxEPrH7OkO3knctTbfwCHKihmTl+oJJDETCSiQ
18VHmLCn5yUeTqWrZe0nlv1DJHDyxwTQU3zpvTrWEw+mFfp6PolyWKNgEBUUD2c/
Bri/GmkoooWgyz9PQSVRTLfexLoJ186ZFcMrUCVSuhKisV2te+E+4vIoI+cTTdUx
7BGUNNRkBwA0yAwd8eXJptdxpaDO0kKtZSWsxBr6u6WlBaeqoNxIbHYuf1qX7kJB
EV4R+wui+uy76lKpZr9uUFOim7A+ZxOsnLJbnDGEFZZZYylDLUSW/d36WdumhW4g
uIu3IdkfL1yqhj7QxzX7C/LVhjllTHEquQW3e0GpH/A057IsDQQ+cNyHTncmh7lw
55V9BwfACHzu9KOXz4T+/hqdtLN44DAcFqpmVn47oPdlnSBVtcI901dLF7c3cIFD
Fkb8eKxDnR5NYOLhFH36WL/sNJ6wXcl3zZko+vzebRWrwwezWTHlEJycD446OO6M
vFILtA8S9PT8qobbGEVKzeFw0GWThZ8NBC+JvMqcc30guIlYwOAMPSS/SRYsO+5p
yjFpCzB8iXCeQh6SyzJ+vgb75BVcg5OA1+mqWjVYMJ/NRorR8rewDQrRHo+jHGcS
1F+RJ55iK4x95aw81c1gd9uPgiaxfCV/niRG1zwUlVL2T/id118Xu13unyOcPjnU
QAUPcqF0OixMX8z3+s/n7JF7DIdLNybo/f17BeKUME6knUcLHb51PwlzhNK9LTYD
u7Dgy62AMqzC7E4TvvkQZaIVZ833FIw2A22PXeCJieOWAJhVFqw5LvRmHfgpkMb8
VwOwTnIBEbjlMaXX7yEBIBp+bEpUt4b0/lnYqxISXe8cxYcDrTkiyR2CSlKzDqN+
rOiOcMN42IXumQywZo9J8/deOTWigBj1DMxei31j0SqwfQMkCdrNLiC4eT9210ZK
641Q97eHsRc5q1vR86xURySNqqC4LHuNcAQreo+xW3B3iD0eI2AcNdb0c3AqSf/b
bk+pxoRQAAh3Wn9QQabsl/uuTSayMdIr9e2+kOwEmiIU8ekmGaK7UqiFpGJ0AI0J
sdQXB334GbeuST+60xYsqUZwgnMjXT2hQDfMOM1txglqikO1SuQOTbMQntosRKTz
Lq6hmtnyWJrUN3GbweJwSJvPQZjeFQm/Gv+iKVMUSW7kPB2sz5vwlwhaxum87rcL
JX6SSlQ9x4wrOzflP5pSgy45MBfdy+dYcTAWAhXfxOcfIbqy3RRpDEBFEVBFdKWl
7Uq38Rc/0ktN3t0FvHBTvyVPfEuQxVXQxZvwO7k/LpXmQD2v2Gfk5Adj+M8V3ohN
asxcSpuPA8lDjRWCLoXZB8R2WzMfRg1T9Q6a22M7ArXBP+GJXWV9OuSyPh2QvJHz
w4LGxOQgIQBx+MZ57pr/BL9rGwkWrAOpUaNNmb+gw0dgp1xql3SpFyy2PR022nU7
xRfQon9M4K4J5WbqApY26R90z1CB75Vu4/VKiuhWggpgNL9ndLivgd65csgVlFVA
lVt2sJaXlCU5T6E6tjyBcIlAWsggzuaUBypEdQXc4wOZpB+qRd+NB4GlkO82r9Ru
hBtA6Fv89suPIIv3BC2HTaE5uI698QdGDdh3f/h2/C/i9VA9hgIuXqrXP2lcu+Uc
lEAh3LGO0vj7dCCOaXqOMS7DGy5ogLdczB2xnHOVD2vvBcw4i/qIto6Br4N+vz/W
QgxrhbYqMQIAM8TzKTFK/xH/fO+kcaMbOvTJHd9Onqi11GtR8Pi+hzx2hwwUHLNg
WDZFR/dqyQJh9OUH4x0D1T64/pzCpeOypyHMlmxZUs6awdzF1d3KETb6qsCtL89p
`pragma protect end_protected
