// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T2isrnEReb0hc46mImTxNsa21UwUB0+eLGG7FPMZV5fnC3jFR8YMuqc5KSnlv7WK
Xt7DxKC0HuapbwQZTDXNz5YN3QZASY3h0myfwKx4WTtDp6eVN/FwScRXcod0WIbQ
C+aUCxmVsbihIAgUKhs1R863UozGncCi7DSgdeoRixg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6160)
pWVDdE9csLwt7XrAzGDhyv1bgUU9YpweAXINPeqMd+mwGPD8Q+jU7/A+MftOAr5K
h0UQY9zoZF13Xg6sC0NZDExgFzHg8dMG4B5s6x7VVcaPElMZkdpl0VsXxxCHqHP1
JJ1B099fL2liTGu95jGHVF+t91WuWK2S9T6MY8RjUHn3bDuOGrqIDCG0tNoEcpP/
lBQ1T7ho8XAgE0SS01To0DcaStqoAWvXTwbKhPDaZ+0Cng4eIupIwcLHkT2oHaJr
gXiwm1YyKQ82JEO3vl6iVho4gWtJmU03+jEa3jmLXWJJGlJBJAmyr92a3jSbSigP
qe0Y5hEfLx+mc6lkvH3UjGuYXUanFb6aF1hiAWfe/pwMK2AOoYkDeF8cxkPpY53j
bRYQpBZ7aopwnmNvctqMv+c3ppjtEwr4Vfpp/tRPqhwbPKMwLqnUD/o0m1e0bXlZ
0px1W+Qakbv4WoQtnwEfjTNLhXuy7d2zntb/QFmdrQ15VASnM98j/VsTpE116Ruq
rQEwIX/Veoz2uG7RQnMKt0Ea4TBBitaLLbnfBcU72FnPG4iBhjVPojKa0aoQh5Zt
tap8vyhz6A2GneJFsJJ8mmHyJ0JYkLRmSfDJGrHphdQ23C+yFPM1md9Wf+62oYTT
Mk25Mnvq65hRv4ccsTd0fpDZgfbxTiwPsgwqVSBN9GRiYWjzPQQZjpkrx4sGAsRF
elc1MAa89V/cvmBkN1q3S5iEGeypFvWDIk4PqBt+BcV/05zjiMLkvKrt4YNAGWjd
sNDr4HsWDdeRr0+n/Zf0hcgGrALresQNFX+v0WcoFptYe79rySB3vSVcp94fGNW2
HyRZIH4eKAfM992NncOhP8GVoE2AhIjxvVreytW3cq7ovVXFEmfEzIpg5pifLis+
tml2ERKldo+A7xdt0DzhjgWcmwwS2HXY09IfwmMtozuRS8VCnJ79fz3ENPX3sv2u
15ofTh4xfoXb83BBIYwb+c4DDIThjVE+elY+Z+8t1snsTHLTYGa1Ld/AgpF7FauT
p7ufNDn4yh/+TgvvbVlkH66mwZgLkGxZBym3cOgopv2Aq24vgatMLdls9gz1S+Dm
+vzSzWMSTdZy5/W5tyOURZ0vjZldAswL65MsXhX1m4jxZKs8h5kG+vUQcIolaTGr
2xpBFAgCW9kuhdS4qyg3nobxqniGys179rCoSfaUFad76458sGK4bMatjzRs1+Dy
q3ZnGHgmcqxNeynugM+z4QJurNQIbHtqYSyS/uYu14Pc5XXOcbIyNAsvp3VumQVx
3oluVNFxT8l03QV7+jvzPolLLixYzQL/8Lgtl2QK0Y0y6slvVFdG68EsDk/griey
1Fzt7jllXdZo/LodN/rrwgrPcRmn7rgbvl7YOMDUWBne8Y9EPW1dlsHF9KJBkfR+
MroELF0jkOTbPSO2qIRtZDsJEZO7v3kfmkqIvsiXrd477QF08fi7Lg9fiPPVFV0p
bT8ZFQUQ7onwtbKmK/0ZffNQ38K58dMfhIGMiewKDxGYEfRQYhHv/6qp2PpWrjup
Oh/OPemxydL2Uv17Gj7k5FtoBR6U+AhdlDt5SmB4Rr8v9CskU69AiybuYxy+XV+t
o2ZtxJkGFwQmo/V0C502rnqhjzET0Eh3CLf0EtCMelM90X3zwF81YGkGAHwDqHpx
+qsgwAzhljxaiu8pkYVPsLqNYw3T+CKt3QqOjIupUDCVxE9RmmvfPRTq5OSiUdzk
jmp1iXg2TBf2hQYmSjOzwEOnqdj9X95BK5tO+T0JQTAyOyWOvSdS5i/DbCdOobJC
08QduqVKdefpzEfNA7soUZxMFd0Vuzfqr7JYNaw3uxNbdobqChh7giKmqnB+2t8+
6iwTSoJqxlBMrMmQzC3VarP7XOERBkCT7pGTzYGqMOsYnReRR89hsAQ9UJjC7dh0
qfuqrCmVTrdLC+iqWpU5vGRa784L7wg4LPzzMHGrmYF0zb+Zk7JVX4HoCH1U1sHk
2ppCCH03jkW6uLeCVW4rxPfoxDMtql6sZPktHm6aqZZQcwaVrhYya9OKSnHzVsln
HuATOzbfQlFssEr3ZCnDre5vQq19HBtgjieTZ3LZ/J33gMaAUjjkMEYy3H5jyKF1
PIR2cDeqWZBOZ7GeSSp/TJgrggToEkQbICyuu5lstm4MtkrkdYqtPeXeqiK3ZRPY
nHdWWOB9DG4/Obne1J2xmPFeFR8OAvvQ6FyScIDbbSkfs4C1iNli0aXXOxlAZGNX
c0w/wnvp1sDZ4uAdYZTyiVNPtRgiv/EV9leqiODCdDJrLwZN7FtGqzZ4fWO88ENO
BVVKtjLHGw0Po5BgypDMNx9M92kIJPJZCabw1kto7UFGxeDj0yBiX5cs8xVxN9xY
FpGhsXrqZZcW2ElcT9cWsSPNAQ3RlHoYKOStRChWXiY5lNDTGuJ8ENSQ7KWurXQW
qJNz/ZIxp/7izCMSq8PgSdyu0TEX+z9JttwB1+X415qlUviKydavzqy6XkD2N4/f
tM3tB9YHSC+G+irz4zfBVO01UQ02ubzirkqz2jQVSGBSCDnUjgPyT3x++LRyoQJT
i3ysuEVPgxtEddAHDJF8UbpP0Jie3pZvgJDmvkrlppwtPWjuzcKqNZolGTUk95P7
XTKE+PRoy/SkiMotcR11tGG7XQnMHO3vBorFmZdcYcyoRyzBjwwpEwOc2Sj4XCFx
CsA01X6cjLxFsdu/6t/C6MxA7X+Ye1cEcfBLq/9WIA3voTmMQQsTLaamguBFwKeb
gJamC+asIwYWDoS15KaXF0uIMeIagEc/Exzk7PBYYsRYhVA8Jvq9cY78TxbwTUQ6
iULdNu5Zk3vzjyuwIetwSSmnPUNN8rqKDeVEJsgf54ccMsSDscdy+Ndozne3NW5K
H5f9lX7E41cuNA3J6nRi2Vy29LeW2kJJDHZ5KCOv+EoSwzZ+ELtGaFcSwufdOXjX
hqOE3RTuT8PalC9IdxdFP2Q30ptb6AMurPus2Xg8K/pP15TmU/7yB7gqGGz1EShw
5tmh01PyH0558mSc3HE0taQNmPqAWUhcBD1DhBAyAZvQRvjRcuZIqS2AmqUMoURu
vvMRzLsVzz2kLw95uT+Y3lyIYRqHQ1Rh1cw+ghF046dFCfXvFPYSIDAzSM1p+d2c
i+56HknXXuCSJzuVklYjy9i+JFt4os+rkBgjV5iUSlhEy/XTUwY/WSFVTAroprC6
O1Y51APP4Y21+zJ59fANs/W/einWOxH8Fm6iX7ClSKYDUvmPM7aNSeo+6pMu8nDA
nq8sNZggx5mHwGSNYbN1c8FjQOpQuD1mmnaovjpFyD/YtuQIYeVP4mAdgQR6Taiz
JZxPq9iFjkeLfUtNhwleftn7+tKy0APAV/44lqvluJHM1iQQLc1R170LhSGzXrl4
jgseldC/j4T54uoJnBtN3iCpV5HVqJQUyeGyDoZEMhkmSOSO46c/Djmg1WCLOK4Q
pdutWGD99FLdv5C8P2577A7kylmTqcU10bqW7rrZDUvNE+k46rL47Zmjuh40qRmS
uC5h/QE3dS1QR7ifVg9E+UcJJIuIODurAZ2V+XFVKtTjCPGK/AsL/xUnPlrmFw6W
MTofsUSrdtADOtnIOjijjmd7XCe6peQreTF0EHrDps7BS50Lef3k792qDwlWoiST
YY8/S67w3WTAIpqr+MD3mGqBesNECPi9fpUN43xgHQQyE+RN6KlAxnCAGI7qnF08
3i6ZFp8s566dMB0ra+x37g7h9mCt3gPib4bRYr48VvcEhKTTu4+q5Fo6Xx8kOVfy
5fD/5hwG7IzCgCbpPHn+XnjodqGXlc8RtxDGzZwH3PoLBhgA+KsCjS8UYjEtOJD0
IJTCytM/o2+GHlX1US7YkdMPBoJUfDaIlTd4ipmdNaaIB3So8Zg/uLKtpIf3utT/
YhqhJOajhbNgQgyPwYd30EHZMjdUVTIXMHavKXj9acFEiP7m4kImOd2xUHtyZbFD
usBeQ14dj6kmR9oOSy0qlGVVwt+3QvAWdp6vBzL95DmTl/3FH3BU5UsH+HayOSHQ
B2BrWQY7Y+u7JhGMbHVUawxVDDGZv5XfZwExyT/E1cI1XHnYkA4YfUHxBoTpZoRW
iAdp6NqtSKSQKxnQYZZnYe0MGQBuUWG1q8oTGHAC97XtltAusyP208+5gpCekGUz
r98VoXV3bws7YunMrsDZx4j//9I9eO53rZf/PgnXk+gQECoGBPFjq8DW/vFsw3cj
FVYBZY0O2QP23Sp6seDSQ/i0faO8tP7hTmahiPkKK2G4lB+1Gict2wQD0i8RTuAP
GYuS390QY0NFUYmDW/GTH6uXMZGqr/SkP2FqeS1LsJL4M5+xpYRsJjcCWrywwa+G
iQf/o4k1MSCmsNZRTsrzkQDCTeSZefYuOlvsTii1uE7ckdmwLRL2ylUWmWGnpT+p
pFB/rTgZmFqTlip1B5ZOJWG3Ku1icmN+6oc6b2DuY/sxcsYjjvQubxo931mQMLta
88YqIYMHkUX9fnuWGN54ENZ5YTEOylks2KDy8vwbNou7OTGOibLr6wDf+VQsIuvK
3AyAQSsb6GlnlTRBQ86iE85TYKLlV6FHISP+RF1X1R0eKriAVAmXkBqABb/FqHPn
laRw8DuNZFJ/ZXhql6bO4edvuw015i9g7uZ5XOi6IUQFtKdSIzkpgff4R5eUdXus
dZGB3TH75R0BsHn15Xm/aM6fYfCOvYaje+Ve7QESj48Ja91L+IJ3X5zmEPPp54Dv
fIvBJ1np/XpGL7iFivQ0QLDcejDdkmWyjdUnJNuPSLmR74urjpiDPqkEMj0bmJrV
Wi4dsD9giucCt8glSa+t3yT+dKzC+BOIyp01v43rIBmwzBsbu+F661sKDfqEqPZj
7XwPUFWLWJ6ZOOkJsgKGg4O/txF4OW5Nk2aoJfC9uqGuwtTGH39Bm28z3RU2gGw8
FnGwCTjaP51jHAGp49zMzi5gJS/m+KW69+oKHlDdAhT3swXTnRqFeGqXizu98P/v
sgdrcv2akU7iK6eTSAAa9QhpAnv/RktyTlruUADi65H7pdtbGGTLc/XBLOkgdm9I
0BvScJlA0A1m0bRst9AFbFyeERXi6YPnG87GRpPwpbTRfUp2RyN+mxxZe6N/YJPJ
SKo32GnYSOmEcurtU06cqfyw/SjoTsplCfBG9f7qc2pOW6dMteexseecTQOkEmVr
vITXs2kkxqoobl5kQ96DYwXVficsGwJZt2J8maLbMPIEMhnFo4vjult6/puYXCGZ
fXlQLIYx/gTUsJcv1+PvDcTdbz3CC58FMwgtr3oMAEQPIRvoT8ErtdOup3PcQ0KP
kTPvTruU0nS7FR1E6aB6mVSOJEPHniDDDePVDu5Xt2Qhcr5xudPwZcrJlFAyCQXx
yXMn1DRHf44TLopT0vwHUZ2JNV5Mx74VR/0o3xriCoDEG9md+a6rA1uU+MBxgDxz
nex7+m9hdBibzbr0k4oVErvMOocVr94p5wQa1uQAq/jqR819Ogp5bZmJeyqRwMAv
PfbJ2MemQ7ff81LwGnMXzQR4sus1mHIOqeZCK4VCV9r6XrqOI4m60QpXcXxrbeqe
NwvCu/vZA6CmJRcm0IWxuZXyBP6dF4RO3kCrdo+Ws/dQZgj1matVbWJaLHvFGvRA
1clY/mjuROeCZL6tfTh+ak2XyVs0J8SR7skSCJz23t3P28wdFzOLu5mNX08kAR5R
E7Q2YHkPb65qyhn6YrSsrjacCuji6xVeOtTb3A53g+JC5rimtenNH7Cbgt7GFWEF
9hPmVFpxY/jjwPAGpyC9NjmPBZyGGgqiZKwosISgp0EWVXtoiV04Uaja9uSsGHut
7xhmfdYBmNyOx6dBfDfK5KXd/gy0ly9YtNFUaa0kXXl1cCrmjrMxo/f0dFmMdQxa
BKl09H3iQuuvAcQOWYpscuLX/GSlpuDIpVKQPN3Et/HRVEiY9X6WO9+RB6UsrQyt
FVEfKZpNRwgaZX6JHjQEosLruzICEbowLszuPYsj053bTKmcqquw9PiudLCIIRVg
vLPV6lcx2EwmdByReGsYMXtVU95JVDD91dMu7f3rTzDS31F3diDSxrncRiUjxHcY
TdBJcG2XxG0b3HtZEyZuTn6ampualdmqTAfI0RNJ/h0FcrYmVuq/KuvOai/CcVif
x+A6I5ahdjHh+wsXh1SFxmuhVX0XAkfRPmsTAfgqEvnBCHJbgQygcZF0Rq/812JJ
zTf9ccTVfsBM5jvERwi99I0aaeeBkuU+0y6pqb9QXiuCISdBc9k33S+AKmTsh/Ai
Nx9+6jfIAH/yMa5nCB3LkQ2wpZehWtvPG11f78ncE9wATLyX/n3uu/OilVGdcmoN
CbOyuWcoWhzwERdpl5G8UGjdXgIX7rBzqjZa4R1UNThITB1Xis4U5uIiVQ0swQTd
pOKdH74TLnxE2ijiAmSiqoK8XOllYjzqsAZjJpi7NhGviLTcsOwjJKt13Yq0I6HK
H4LxIiqTPf4hQE2Tty6UXTVAlQR/jo1YWukPAL9TR7NmC7PYlmy3miI8nlXYB/v6
6GWT9zu07Q3QvNZLCIJ7sec35xh7E/mcUOmQtd15Thh1yvfqEL+ehh+apaQbSpK1
Me6YCkVGEV2jOsRZgAEDK8tWIShrMyC+80CVC1wKzyG4xYcIUymq2fRcK/A94Sgt
8zbBgp7tLcWp5wpVDJK2znrnzrgeCzTZLKUYwyIhghF391U+D11SBBLF5k9bnjXF
bxfgBEy/VHuC2cHWJ9cdZ89BRRebAkrFUWzu+7SKkqvbnMGBCzBBFP0+p1JNGXgF
xZnKUff2BzfjMbM4SYhJgpoYctM2dzkSVYTgZbADV9w2zt/lexNRj1Qa0J5fHku4
FePE6Qm5la12S0K/9UxQCnsRnbmR99tY89uhFpy1FHW7+LKSgr4N6AroDdb0bNV5
UUEA7TFh1CYoMAre8bkqmfzqnDXhyOlOMkwtLRC+MZNeb4LfxD40FsJQo+OEv8VE
1KtUjZj72mkDr27p2E/lX5x+3M/1ZONofCUAbz85o3DFAXM5qo0XSeM33tw5Oi7A
G17n5GpM5FAyh4uFzDzmgl/DF5ogm8yAAHjuPnwuwnmj0J6Wbek3w1W3FcAJDVGW
9PdJvLGAJX88HQb64y7LIDhPpMaEvM9E3pTeYyucQ5htCDMKQMo5lJIhn98Kwsx1
hkrSZ84rv0Mu6Vj0fr7MN0uyhCFuLG+koPp23FHrHp8w9zpiBUzs9KMlQKU66YUE
0+HWCYsSV6Y0Dk/EqQHrrS9qf8X0zT0SFxCwqfjmbpO4le86nrykeumZYSckyyNG
wnMN8iYkBrWmxymreTBJq84WUWtVqQNm5ibI/R7c1jspbAWFvXt7CMLggB6VuiZl
ruP2UNv/K9VnDo8164Od69dNEzKBWp9oHxc7X7dVZlG9wD9bcceVgzKgtZO+H9Qw
Tj4qjp3NDA8Yxt+U2xQx0RIHu7sMwFTM+LsyRPb5jyy9ChF8pnVg37BgjhwsBl8n
6ExyGQtk5agSZFOifQ3gIj1KwoiyY4M1wvWzTxIUVh89afkX2ASQ2b/+0SD6JSgX
PkAI8fbhrHG9VyUXRHG/9nLpAEbFMDQaROJbxzOTb0zuX2Br8aEBXV6G956zuMZe
Phi3J+Q8OOEsWy/OZLDDluLsC9rN8V8KsKWGNBMSDnwSC2gxyg7prhv1lr5Uipni
wQsHcopAnePAGE6dnhtl5llT9HDITaC8tjE8qThq9K7ypcOLAB6yr63cm5J6MP+L
o+A/F8HesSm4T1mQid6GXwcaue8nu8q0icTE3Hor03ybxrMfsOlMXlGg/xkk8wxZ
p1MPcOm5fpYQTdbocMDundOvV/Be6n8Bqk/h4cgnHBQqSr1GjKpDevkWgKzh7rma
TDg6jX77eH98ihj7bioDn0bA4SmwHesSgjaq+AhplYduwUUSQjDk5r4/8dcIx8rs
OXi3DBBcB1J205Ia7p37rxPScMXqkvOo8xcmWtniMbPOfLgh9hGQTV4sxuZdQDNC
8f0v2pXHks3ET+EORzQAy1w+eUYNSY05VcnRc98DLMoruIvHyKN769tBcWXGYL4S
xTSx28w6PreWQRhevK5uMu6Y1siF5ipLuIvqWEzB2NcXsVdm7/PswY7GBigGWmOY
w6PSGfwu9T1RwyG0TF328SAqwpfLOtv8DaXip3akKCH+mBQx9Zbux1fNx00Jr3l6
Xe/HZQfnzi846lhlwdIP/w==
`pragma protect end_protected
