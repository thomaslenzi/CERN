// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:09 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cUqlUBk22n8EiRi+wDvO0RDs1lJtHP++eeqbtO8xvpMZmUuRHQdrvV7GrV9IEPqn
un54suwB0+u4a+vg994vSHuayKh2H608n/anmF/0vfJiwu/o3vYfqv9DowmMFQjR
hDHlnvYd/CVF4SmeRblp28lPmXdLwV23Nwzbk8txBSk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12784)
546J0BWebOovuPuYfshy2FgZ2DuAg2iO9PMeINwam0+u8MIEZqzWHQRxliTmJgKk
mPH2n4ETtvM7oJ7CFAxOxcKciDSzVrnE1g6fbyjDKIVgK7/EGJo4BWs1cMMEIrBm
AaDoZYm4HGSlxqz2TET+EdmpBQ13pgD5BQE7PTlHXOXkBAV8ktmmf3E2Hw2BIuwd
Xr9HCVhG/z3b1G8A6j/4JMF+SivQxL01U7/NiPXRkftdQ9PDlEsPVKqolLkFYAIe
qHn7v/6aXIsFA2dC7deDHB34IrOTTblzpECvyUOXicI4pzeVKaFTkwLPW2ulKZzx
JmHWbZVblp19fb211+FTLsBq4m4StUyNQW+/bL7UzaK1bgfd5Lzf5tgJcai7psiG
OPzajTAR9D0t39GJOFYrN+J/XYtmtLhbriV3W02faD+buTNUTNgNbrWiURnRVNRB
vwGoWJMhXfnGUige1Rq/MLsMadAKz+8lEkCEkqAaukZai6rrnqVI/ovESB7LyQuN
3XN9qL5LnJkVH58McalpnJil8jz7J+jlvLjn/FBcxbHD6gm33Dsi7HV7Ers3T9QO
d9UT/9s/lAMtBbOcrtiIB9D2ttccrnutFI436F9B+2QkTmvN8ga5YHhryaUfuzjB
GQj3frhgmMzFhX+NTsBYR1my1Y+WUJXVibVzOiYolhJoBV/+Ei/Ph8VRtl82KTo2
AJA7Gvyw+/eNDprZJieFPDcIsxg6eYChIKjr8AHoTbSvRzrKR+ROQUN3a+5GlijC
O6wfP7vbRgxC/xDHbGX1bdEbpkTWafjyw56S+OcjpEStP0Yo5RNJyAtO1sxXxt95
DbbgSvooNk7vhQhcIofXC7Tv/LzfCPW+9bB5veeVAcpPVqkBXFjJNTFm71a5uzvv
eqb9MwXoy2VN4nLiQrwmM90TYS6y7vIJFWGJjHNG8f1dEzUi5WutG8hifRMEMTWt
hWFgxLNUGQdflOhp62iU1Xa3VOUu5h+3IPq83tTNz152BlWBrzHLhq9vkTWy5I9p
B7wwQCESD2BWS1DZAlcyWJck1YucYbqQJzLZDBeHV2Dn31Lb5RgxHuitpatx9CNB
F8+YW6jdKtJfCNxGTJyw1XauQ3pJdYyRPXFSU4P0CVGK92ElJQb1v+N/V2D0P9DX
lBaJL8byTwf74enhlAZDkD1d1kTLT04W6n7uD2b+FUgmiUUMf49sPdmLDXtvncj+
pHYclv0391CtdU+npuuOxbJnpAO0YjIhNaE/MFWrCo+A3NiHrQS9v2riQ8mwYfdR
OPrV4lN0Li1Tgtm27ypmhCi1VnN6xD74bMqJozCHkoDONek3kxQl5BUjWm86wzbo
6p+MUaYCaE1Bd12A8I0uujxQ2ZXNvq+Ggvp5558CaohWGoZnMDddHDa7Hqy2ke4q
ZgpjKQ/e/WSIgYN31kc2JcRZMlDYHg/LFh86n4yX6dqHyxyJt53YRZGsXAVvKoRD
iarV/l179/UZYfWY4yjNdmw/DQvBnAsV4k9I++mpMzQapU7VdFQjSscVpMZ1qQSZ
msH0ZzTr6def5BvFoC8M5FumFK42DyUIe+6FdWJP2a1xgrcCy6Y8f64lAhcIsB9e
V0OKmvEptBglm85FkfhEUjDtt/Qsu4FM7/0NFQ4KX3IcDHpCw0f/lM+FGKwCmkuI
el9C/QPUEVs/VJ8U6VgHzgpa+4Wvwisy3i9z7cen0IhpVRtoFw9YDHarTfCG3J9M
Hib9P/dq8BV6QRN8Iefo7dUdXKIvi053lG1QbV9KaSBShuRqaK0VdQ/vWjCa5k4h
H5O1gR0lMjMGTIvxji4YE7Fife730NzcAmzQCD9eGIdfI7bindnGPdGCyvv7RchC
TSmIRMpfWAB53Yr39TxwWrFIfkwoVeq6kvuAFP5jKL7ZhMS4chp6sP5PhXJU6u4U
tLQs1SU4uOPY8W+iq1bzi7V44kyBCCHQYjdUy2DS317CP85NgclHTywo65iTSGS8
XQ/zMtHLk6rqj9Qr0xGCByRC9+num2KbRFtfZvSI32cnVt1PpRR9Msr7UOYaXZtR
RBuceW9OtMYzKALlBbzjz3+q/RvKZp6rL8x29TKgsXCOTPGl7Z2PTHvbOACqSGO0
qjZI0Vjbseu1JkfHz7DwHjHwT+XZI6WF9UTtTWTnxxcRKokSlE+eu2wEodbC9Q9f
S6e3IxD3N+VitURtO68fi0yp9WesIwcaHcv0otsjwJD51tFBgnAVTT0KhHCfJufA
Z0v3GageKBnOBBqL1iBUYiFTR90UfL2ZPX5sSnxTZFeqV4XSmcM9A89Zv6RgVKIc
v6KnGHIlN39AQf+xW3fNklIYUi3GaVcIss/QA1oVWmtZUYQ7pDXsgwmWC1XYbUbe
h8OUHZw0bHxdwsZfLT5sMP8V1t2ebtD8JZTOn+abEWBfYg1aK1m5T+t9yU2Zmh/2
FFWc/5FR2qcTokUcsgSpWSUkBczuAIZtByhWP/9JlUlKT8mBQdRZwvzbZQBYbAUQ
PcfD87WMhLbxoa7hpOZFXg4L0CJQLaixmVQCVNyRcIhofMiIt7OM5i5epj34DJoF
kU5mGw9pLCO6Mrm0JlATLs//pWotnHvyZhvDkUGgR4745uX0zrYuPeRUSU3iruhZ
8VXEVUWr/QSacMiDrPx4aWn6SOh8s9lIn/YDyy52OibIkusY7+o58Qd96PBa7yb/
oq8CHahIjBD6ocDoVbjCBHhbx3DgBwtMidlMdMPrQ7n9bL4lZ1ufmDnACO8QluFc
O000A3KDXbp+NMvyMxHlp3lrtcSptdh2ui2F2JoFLKNwCsbtvRTx7GFJ3QNUO31X
EMKWSnocSXC7d0cLMTePBlSnISQus/nLrvSHSYFo4U42CZfs0eXmoL3XFqr+MTuH
xHWf9mQLpq+QeBxzgcTIKDTrpJaU1hK0OQ1U5gDB5GqOY80lcHWZynw745Zm02FM
zYHAYp1BW398Oj5AIdvb/Ew817QxEsdlWkxNMf0MRSflGjofTgCQyrU6ZHG9x8yL
EpbgnbXMd5miQyuM0qRfGOwnyXsp29YdPkTPKMI0lLu2o0kEwrQ77lPFRWcBpjXu
aiJpyn7TcZl552UlcPQdymckOy9QvyNjqnUaaYTe7vOrqf1D5tDjre1wP2Vdj9q9
LbAJWhSVGXNCVygLKsJ9TmwHbSznwnn7RA1sNLgVtlnuz+7oUBlA/Gx26nG/02ja
l4AW/C2vyPMjNdJpH00q3elfddqGj57NekU7J9+VUGWIaud+CwdFZtGsBeVkx0Pi
w1dovHzyfZgmAvtpz60sbISkpg3/XFyWxZeJlbui6xLadVA41Y3UL0R2O+DwYTbH
+mjcBzxeM1bgsLFTCMRQ/jzHVYxhGich2qqYPzGn/6EorczEREu3NyqSZCpDprkU
E7gPu3AqaejyRFjfoUY8JTFSJSizPn7UVAtQN+/LckqhyhrVC8z9F//9Q9Bz8EOX
rehKWt/4DHhwoKtMCMyCtSZgKjX4NcHO/hkdck3SAuJEDdgrxIHsTccvHSzfWcYK
QLns4JWEVV5XoYbCOzivnf5PPtM5qfuwzNE6QVmJmZWcW+Mvcqh0Sp6TMrv+hotV
jPmoJk/9nWGuwO0tz4pVRaHkRxsWiDk/pNNGhWSp1ekMnaBoTovS2abEvxshbKk/
1Ha2F6PvLfyUf9Xb9en6mo0wWHMUbu/gQAA+2x+pRlQkmCORgvNcu9dnupIJZIoP
6lK8qG/9ftdkm2Wxb2s6DQMMjdPqsT8WFdCmnMPj+XohfRvSB+gDlDuniGq9EJMZ
plDbRBRCTWkpsO3EsTpV4LnmqYtcLhl4HArsHm6112IoueZmYKx9KNB4+biXDf+1
zTcnkjw649G/KGCma9ZISSJE0M37Kw+jXotA7XPpC+h3cKyJe+PHbPfiHNmF8Zjw
DMmORic0WILsR5cgZo/5BogyQ/HMnpKF3ghR4ATQvuKRss4FO65hzPkVqiEntZwg
MWi4PUYi2K70RgS7nVAEJtwjjQS+JkCLlCJ1qv9c3KoZbuXdS4ZKjVBVm7sPko7U
6vLFlsI6L+suY8voNbmXua3gLhIalJt7FkTGn+s0RbBVbM6wbsEwkIEujmksJkir
qOwlkVEMkHjgt6YRvqbYyuliQ/EQroU7XWELOk75ToLOBNuLLyh02HOFGyoCZZSK
vrVmmpc2uu12h75MK0rO2NG1IQ17fK1IbT6qOaugAM5eS5CcmSxVb/zp7askxAyk
0ZvwM3f3sZxX+u7lV99haI4UITz45BoYLV7KAnK96GCmn84tWShngY171f7OHf4U
Eh8wsCCNtXh/Bc1SWW+UK8V8re+M+4M76OdpCN/W3RaCNdFkufi3sIzosTfsp3ep
2KHsALyRBVUH6WyGU32cjypHPp3szM8dklVp/MR7Qbf9A65aEvvb/526zFjw78sk
kGWIkbOWDgz+JKHngBZbXyIiQdU61M1vK9++KSZ99FJmDp8IOOxoYPIQ7WKCTF+B
6ytvLdrGPYAVFA///AfTJfdiNLR1df2YGxB/2u2RuKBkbjsyxPlCQHSh3FaHaPUc
1/RlOQoWv7II6zW+rbi1zRU+//iyeWBJ4hVaYLCmN8PdrQkcfUMOPoCsILeZ2H7x
rHXVTt1027fLsOiKVHRYr9Ar5ChG2V4FcJvVmOv0Xg23mumF2TvPdZFctHtSha+M
zGYcpgK0wi8OAMzmYsOlJKUZAR+pYzUhZetyC+17am+6HDcKun2MHCbkh4YMpR89
zgF841dv8AmVOb/+ucLEDyYFOV4NwI8HR+Kjaia8Mfwueuj7ZV69odTW00lNmzXI
YlVL2lTt7uXiObSzPgpHtEAyENqR5HYlhQAfrioAOUaipgnit+RQsXuWuoO1hwtw
g5I1pVZNJeNnfhFfs6CVA19lllxaIcsSm7jqYCVI/+A9RpdyoqFp/VUsFte4BDxC
7pitLV6upqROyF/NBsUxDS2JieBBhae/V15bax2ezYa0LA7gmnDfkxrp9JSVA16e
tEpn5qIQbT/yc4FV2DISU4ryZyKTRfpSWj4+6kPNvXOJbqcIlqnh4AXdQey0BwKt
ikQOv9qHziAFgEnVOoHb68f8dZc//nSYmspe5yOXpE/UlpFjZBfmC85WcATzlhYh
YB7mt5cU01e0BRdhHVRLw5QmTO/O4iU8EzRWMOCl0ZcDlmpshyaod0EmwslxEOqg
Xyj7u5EYUnEGmoqvi+JZBhro7hkM7DqhBzperRx3GVGICEzSgkWoLjqi5Xhvxzo6
vwg/EpFJgufOWZuNqHZQ8HpAstKeZb0cHV0C0d3CX6PSgPMBq3iGVi89ILtzTGKM
yqqBhNSk2/selK9zraHnv+69OFvlAiHET+APFGnbW2MftkoL7v98/L2WjF3g7/Nk
34pFkCLzGvQGpCzy0eonUzzSjOMvneB76vjlQoVfy36VQtJwU1VBRRmHvIXEERx7
7jz71WPdfHYMygppIe6J225kqXSKY8ju8XCNql7YE1ubQKlVhMyztoGRLPy2hCCS
cwvfFDm3Ax/58AExqfqq7J0Fr4JAT75Vy39ezR3z+LH45BIL/k0ds2kkWVMoitml
VWPTHdbfHonS/q8HfyqFkvaowa/rpHaKKp3cTdy7sQWckgcJ/M0o7+EjgkKWkfbB
pWtjPxJLLTwUUfViwNKwsLkdDSq19wj6M9nQlJoMp2LdgeiVFvCrOqCT+w8SbABp
3tTo0x/IQW15dOGJFW5ppKzpgzOU9X5Tfw2PiQsv93z8YmrO8TcwzOzgueKPQXfF
kdJerdExJMEhjrGuCFm2h3LBNKBWbENW7eK9zhgiXvK2DTkpJ4R0wnUds34tQum9
3vxZv/B5/vIofzZE6p9lPY1KTFwZNms6hkd0xAvGgoGh+L+FDUxa+O4ixi4mxt6M
VcmUBDCmO1iJI11VDZeCDoEeZtdj1scAq+fZRu/dQwbAhmispElyVZCaIzCU4LXl
UHas9Yo1kApoxuCuCo+H52OUkG0fEPnGBwAACUfW6483SJX1EC1ns3Otj9yOF3a1
xBTBhrvTBvhcXt7gv4hsXfXL0jb1BDfdYJRG5Y+tv+O/geKmdId9zDTwwLe68uQE
rq0cs5BXvbFXpE8Mem/vKY8fdYkgTB4ynr3tmzcg4lPUGbi43kTTjc8Y2nGxBFTK
+qwu0dsWENODHaRlyZ+m2RZu9s+rwOnBxYE0NnGvXVg8pyzIHAXL8uzm1I3ONsXt
zdh4+SadY+wERpmn3K0Tzx3vZAKv7A1CpEneBW1jQ1TG+wEGTj2d5M5v3MjbgQt0
to6DPlbqTrpGbXWdasQthWhT0JNdc7Kq/onBDkIgSEFWNxC1s7jE3DdyyOE1RYBc
wSkgkk0GFX+7YizjnfR7Mu7Km6gtQ7aDhIlKhtIRfqgqN//OZaLvymhw+siQWY5t
BfSMC5s9jde89LgChX9gS03cRlT5jidnRFdsfaDKAJR2wIshgFey/Q0uVPiKnJ9m
IH+bRIANs/AyF6pORktS/8ThFdk9LITnM3apJqwTd8Op5bA1zsQQdUr4VHmd43H9
OlNuYSMrKKpYQl6vIJ0qoNwTvpjf73EiE1kaF2l/D+fxdQlzWB8WgGgDcIqqqi+2
eCRwhpNZSUkE/UXQLE6L57f7rvg6BXbQfPfVQ4p2FC57FdaZYdXXkpblL0khqhfr
GGPSYPtpiLVgtHcvGsTiale5zRtle63Sd5z0p3Ao3fdeVe+nBerCb5J+aLdO71yK
pxKdXky0i9uXysxK09Mum4aGEm06Qt3n0BAivaMXCbCmKZwS4/Shk+JTLSSxUSJd
ZLYNQsvgydWSRdJj3vbNt0s2r8TIRoTN4n+AwdpmgT6gzRzX/DvpIIr900+ta78P
Ts/xCEKswGKVExZRXO3BjLHBH6dMrPgeIO3qknZ/OaZg+DQAyVHWfP96e/krVtyb
K/O3NOxULxLc7Yga4Djw0H5XoVXEi3xzYjrhqD7t3H4mKFyhS9nlzCtW72xYblho
pf4MxiJiQR+kdo3d+hTYO96u3jcHjrgsH9yaKRyveGfb4gGDQEa+qQK7XVdZzWun
f1MBXWLVJFScs1ClvUTSven2ij7bLXekZ/LpvTxt88+GVR2sSH3JD8fq7XM8kOjE
i6Ot2hmug8iNyhNc4ulSxo71rP54GS/WNf0DmmO1ksfLmBODCX+z9smtg88Dvjdq
i86O897AONuV09F9HZEU5zJ21cocn/VZtjuN4bMOliNMZTKlXJTnjJ3Mrqkmdpdj
xn/4dD5oLvMsETyJAAavi3WlvTpMv5ABTGlYMvwSoNlJLXVg95kFwHs5VDu8uh/S
/OOhiCY8oT8OBShB/IG39GYVzJG9GXzfLFRuWA8x544yy5jk94MoAtvNaKCf72T1
TtyhM9HYz/Q/4YnEPCTsXgWggR4TEaPZRyNovxzCenH/S4UJXvsVBVXOEsRcA5jD
VMDXimJNQlxrEWNXPW+0TQNAM/TjO+TkFVZih3Lqa6xOnvmbF3jLb0L7/KAjczcA
a3tpM1N5furyrMApOybbbCHAyQtUgKJXQQr3MZIeF2kl9jAmXb5MOtxDSNlSnZ1n
lJdgvd3C+fViJbBzuCc7LYVlW6I7BkPt4dZXU34rTrFOb9K3ZWtUwLvYNHuRwizj
D+rqh3IWqWVrCtasrRh3z/mwcXSN/0em6e0XFy81lL7zxILNhRlnayUe5rf7HCUd
lUn76WbhZn7GfoLhLQ7l2TIo3mVvegxb3YBkv5pkbSOxifpfHg08YmEuhBbBPCpP
mUGE+aZsznsk/i1WWkpMPjrulhkpFnwBT9qP4iMrjkwHqHFSOYkNlxL/GG3ffB28
oksxyFlfm3I/VPgcUWbRgzUqAYZhtzx2gHnFsPIoxuZtDM9NdyRABrKU7Zn4dsO2
AyeNaqW53MhASSrG0WYCOjqWxmJ0rjScU4WyFth95XbMNw1/zOsJFJq4Pd/z5f3b
2zw3OSjLh7Bz/8xcFGAf4EFp7LMU3MvjkCqGgwsLeQ17KhhFEVwcwERoaDy69OVz
F773UbctDIxp2kUqVF0XU3fY4UJSd/bwlHrfE8BijgZUoYJaNNc69t+WFqApxtVV
RaSxmJ5Jdp5LB2yUs/jOIP8ERKUdloLMiy+D4sqcl7IOWYfLSKim8ClTwHeZNk38
6OwZU5yesvgk7aBBzROaRKi9V2QxIXJcG6CxsTCCwe6F4zJyrBY4ErngO4YgjSb/
eZYcKR9+8gmm5oe8zUncbn8sChzhPtWdSc4rfDLT8UyuhoyEFYxFGGpFHtg771FM
I14NPQ7Mfvmt4Ynnc2hhBhBTiD8iFE5oXYyUf5Jwelp/bMIGofsaTPRGb7yUjNZN
Tx5hYwrBF+UWJ711zD+EtroKTDbY5b183lABSCG0X3k8XkeoeqN8h7L99/bPoq9V
icQBP8AHu0xEOmAw5zjUS2m5v96KTdIcjCzKM+4qNu7q8JK3fj0gaXOy+vKsgkOC
uyo0HNA6Rvz+I7E1cdRvCCg0YaXPaOj+2AWBePrPDcMQ1+pqXvNi4soe/DPvuSGK
guY2eXrzsE+cT5FDu2IsUWb3UqQdpxd5JnPOxYEmEmYhM5pgXtQZB9bX0s4aBqZG
LbzVXV0k7viZNMt1r0/RqNBdCWozM7eMt2hlAbHySD+E+JEXbEkmbT4Xd4Rg9xcT
qGa3dRwSEA5oYyDlzwLkMWgqTCkiNiLAWPoHbBdZ1FJBn36OVmd4EPB1B0hDNWY2
bB6KmFYMWhmSM+yegasE7qUcisJ9HkIpHGZBmE1T217IeY/fg5pN/XHAXJjfTWeq
vzsZW6jTKkxYaLAKhaBUX+TF19OEqozjPhs8Huv9irnLsEThmpRPkinJgQNKAFm3
zHETaYddZieMUk05J+I0+0CLW+iZHG1FzEnBFnnpse3wBlYWydtEswiI96EftUUq
5A5t1UcVz0fXzSAb6UJZFwBsMK5X2bn3A1iNjLpnkXSyveXs710aUkE2T/VZmLRF
DxPRv/Ce3vBkELxp7d+/zD6Qazpqgf+YyAPa1nU4Q7A44le279UKjqld+Vqb/1yJ
oCGiwoi9HfjE8NhYRJYafzPs6V84D7fA+06tKuagcULezDff3LmhWVjQ5nfnGmGX
ME6TfvMIPnHpTr9kjreaaIMQw0eKs0D79qmti3q1uP7gtTLiNjZXNxvTzlUhPIRJ
i8dPHFx0S0opDT3P8o6VxyCazdNWDFvKneKAonuKl8pFAl/bqq3/x5vfJ3xMUeAG
mJvaIsKOCR4ZBEtBBb8m+szlpKEcJ8FQf/7ivxvQPwn7xHmgxFGq/nG7sRA+t3sf
g59wyiIBcUPyDZtci3XJR9rgMHoSKp5IKGYytVLuKFQKg1ElIK5njVoA0EOHq81Z
OGY5DckjQA5YWOFoP8NBeKKOuw2IVwCS3toKH5F4Vk0bqft5fhqM8jA/v6fTVHxG
Gtdde1W0Y5RX3BqXApDfRIDi4lslqRGDNsVD+Rv5wrnn5bPjgxMZ1wLBHYL1LkTv
k+ct9adZUZL3LUSl06/GwKKK7bTPtzOKmkGtiyO+vBl1XImdCPLoRjJtIx6mG2CU
K2mbr61cDMYp/t6Vnlmuk87KjEhof/iuJceGo26eC3i7lh2QvaRb5tFy9Epuussk
UU0pZmxV+Al27KrQeEohbNkvm79x4jgKAUtk9nEDynh0ZlLcpz95Id5G33Pj7IR5
neankeuC7iIrEZvum7DD8cDftoif8US2GwRJQ57VxVvrh+ngt6h9EB7TOyG6ZPL3
FCGdmpE96go6mzmDN3kHiCTJCbPv4zIUm0qqF1kSW4NAv5G/+G3opEKSP/tksUu/
hZRIl0BbB/pvzS9NqFeqLqu2jKt9L3rE6IXnjZqfNdjx0fTNc614KALjzE9ESA3Y
1QJIWmdU/SSueNN/xEak5eNBqtZBzQXwF/E/U8BvjhUaJcPvxUL0huOdBe/w5nmc
xvFBnmoaOlrGekDO11Gw9tuLxQCvyUWs4b6Ad/AMrx6UnXT4qyflu6sjFdWRVIrP
m9u6L1nnt4AB3kEgRN8B2IcfmfQKazuMJV0Dk1P0MDPAN6vUkd7+Ckn9DtYsAzA7
R+7iFvX7DHtfs8seLfY993sX0YPuBVZdCEs07WXapkD8GbVlWLkJCW99LVyevUsh
5dHQQjF1rcGUNwelyn2i0hEP1zkP+s2TjGDW/ZwmC/uBFIKBOmPtn1I+/TRPlGh5
ESL0Xe4RFLhckmKkUX00fvisUdnz1vOUORT8P5ljFBe/Fo30+L6WkLYHO4X2nEEa
Gt4nTTkozoyjisK9sAZRFUSES0KHXo/JDlU/Qw39NhZy1h1DFTPbYSXWDeTxQSfy
DmMdBjGgJwvWR35fnRbFKuJnmT5XrPfkL+tAJlLRLbHPIb01rTDlJqQsicfHww5g
8tRKSU41OwVI/2t2YUKq2VVWzI+90hhzWZhk8CGxwhZo5jwhpXyVKbNEiRIzm0X0
vBU2ofj3tsQr6Ywxy8y+wF8WyQVtPhMiYC9KbXx+QCTWrtTU8xqtKqneqWfXodpI
j99kKuWOT8SfYV1XgI1k5Snbd7dSb5bTubgyA80L4CPbnRkEkrEKQcscTMyrVnkt
sqkz7PpmzWkXvSt2sTtQTs9SxL1ETZ0mFA2x8fhAufxEnW085O4nlRJBZAmL3nDX
xpxEkFTcWlEiuzltS+CewRBKcRC4hRBEoriCsnDF/a2V5v35ZWRiwWWJE/VxkpwF
p6DobbkGUL5Zv6VOZjJEDkgbdU3r8vwfYvMMJdrVF9dg0/ej0AzICz7ZhyikRJ4Q
xICQafM9A1HL++JSyAlWDegmHuvqf26C8aJfhis63Y0R6bV5QYZc7Vo81hEqErOV
m5jRJcHco3bMiLU7XZkZjfsWoNEyVYClTenLmP/Dftg/jfKqqlkLA3Zcn66fXZVJ
Xc8+S3BvLvl7SB4tIZtL4GdUlWth6YmZHvA3RRy6dZxd+rU1fHHrw9gsT0DbLys1
NUzjbUNVUe88QGvKTp+iBM87wQez93msgSfQUCPJ+XR4nmJhc1mfHchB0ARd9PZN
amOATJNdsLAg+XZ1Ue4RXRTQ6Yr6lQreaH2TJ7tGNccj+uKZcxun0iD9N+uGJ54q
kIfeROvMNj3Z82TAoX6q4yyGp2V58j5jwkSVbejU+qahWwdh1ZKFkbGoQlGJ7nI3
Arw8TQ0cSBc2XBBwENAEPqu94jXhFJMjWS6XDAHKkCWprrx+8L2FOGJZBM34+fxA
OlNBmUstusUtK53n4FKJr9xCZTxvUoDcV4IMI3pSNMWNNaoNFp+LuwjiLrP7EJb0
P2dbGY+riGfo15tUmJcntgvs8MYX4FjvJ4WKgn9rHEH20t/mqLsEexyDds5aoFPk
5WdYplW/9fF4cNVpcXVNgFStvsetyjXrQUhASc/j8PrGPcscOfzpP1MrPficZBbv
sYQdhUTbOBkW/VxaNMyYF1zCMX5zxhWDldli+N7mfoJMPSF50ve5UkYDPPKfkBla
5O8sAaArQsuLouI9Ir6DKCwLGtzJip2Jdk0tKW3HGZrZMk4sfRknaosJDt9h54dq
HZv4z5Zrj4fLkW0AmdYaxev8lZPA+7mM8ihiTmBgTSrxiTRuX2sq9UvyqHRUkwTW
a3Kc1gu6fXELJRvlMBAFEmt9PT+gWo3olB+zG0IgcMS4IAFakljcQkRV+MGyl2Bb
6t7L1RjyyMEnYjZqGQZDFdb75nGXg7YS2VjrrwF6vnqKqQBBTuUMy4DbuXvyre7P
XfXh12QevWfIQGaDOungUEFKFKokFBvVbPZ/XjkjEW/r7pTu5UI64wCeC8sLVrF5
EXuekQJQvK2G7Lx3vGQSxZMJXKalQ9HXcE2Px1UIKQ/ZNooHV0obg392N0qc3j8i
jXVvSArY/prhjaIpUuIi6stGlU3P0QkBrHbAN+qS/bDRxRphx8xoPqrUFykqT1s8
gR5nEBw0HaeUbiCXllOHv+dZNGbB8a4TTjAfsEcUJag/x+0tlJy59xArhme9pN8M
Upk2fFEaBiVoTlcK56i+QNMyxE2kEIoYKbW2usythPcwUfwYZmyytI8ImgNdDFbB
LP0a3YSloadLt9LHeSQleI+/xTB7hVW43y3O8qKp/cVilfeo2EnrRxxHXs6gozX8
UG9pUqycDBUcSaB8vVJW3KCh3jXEr7nx+eIqsZtchWsV2tXMfDx8BLecYEYKsnAT
gWhjXS7KYwGt2yPy8ZGxe6QgZ0uAjUO/UOLMhz1fI3nhjU2H2XXiFpD0Q6Yn+l38
hjDR1Cu4bJTUz9MnObnMKawPldwbPZ/j1ETUXxyqfcL2YG5Kp0xvRGJ3xF1CxP52
Y88Et3fdtQzqdyHDMxudGtGpMW3L9564gEKVPN2AtQ9dvx68+m+C5zi10j/ggLlN
awCRrg+FHNwLC1C2lMQeyvri0zC8F5t5lGlqEvL0cIIJ0YJ/HHI/LWhYl2broKTu
duUwLi+3BVv0rdPoHiOzrvMPXvtq92D7titc9RNHJ/8RwMveGcYoIL4ihlzW+f0T
iGZz/X6QDMtWA1B6xcFg5jY+djD5acVz4UT0FaTHnMXffGVZyeoZ3fPl5lNhCU7U
CMyVSUoFmYrC3x7YkfVEeB03+v0DK8f10WUhA7v9S78SD5jSa9SNif2Zak3suEBJ
ltU87PC2H2mfvaTulm2D9k+gxuIceG4QZ0Vd5qfaRJBm3ZKnWOszo3mk/FDObuPK
ha6vQV0T6LCj7Rr297mg90LfutzvLZPRpcYqTm8DZuiVHWIuCuy4MBPyvFXXHXrd
3BuibjO9GyE53oBB1JFRh6U1X6F4H1Wc3DmFHlVY1kF64qB6hT6i6DZknxj19Gm8
Y3XynjzdYRjLKY9j+B70ER+iDY2xNfOnwx7vyTEcchCOtB46XO7Vitfto2tcF/MQ
83ulvpyMYOvnUbNYEf78bNprIcSpbDIAzldJSIyUZfdN1ynwKcI6eNknI7PX/5cd
VvBkp9ksKLDFHxLWo/85AWlgBHiDupswno+nM/RAh6jzJnexEwnYVg82H3fnaiWv
y5Zac52cqC31IrsLn0RWoyJ3/5taefOOpB1qknmbslLlhK7NbpRnTcrNtcbvaI8o
U10hBwRA+J0abhW7A1goO6c9OqiVk2fLXjHXTodxT8zGkQZXnnB0L0P1uRrYAf8R
25ADs+1c4cqK10fktiHZquBHCOF+MUovbquW67LZMs9WQ23s/nYNA0hgJ9blZc9/
sECdYzXPM0ZkIN5wwzw47F09+T3kv3vGJ4yrDCEftqfwEnCaBt1SwUd/I2PKDzy4
FIWjUzhf3bFvxxd6cG3cFLnuJgGikmfDNFgFjTmDBm7HAfMlowCxWsmDXFS5J1fU
FQmtFe+2EpKzweet9Xv9UDD7cXmFu0ioWIPQH8oH2hGUG5cXUtJEwXJ/EKrxvd9b
TIdrNb4x+fOMb/B5+Z7o1d3hebzGSJVhAxNQyPp3x9Vb9Q1KgIXxUNzikyg+jbyF
UdcX+NgSfgMtGSCFBWywxyztnvlwcOm2h86iyn8S4Ss3s652OfuvcWn4HXAzbglx
/OA+E3LTb0G/aek/qrWH6GpHxksrFZtT/EvKwI10RHNjX6/lFSK9LgwrrcfdrW47
7mu4V/9Wm+r/UktCvVuUy9WhBDF9LVGI0vfJYvMKj7vJk/pQk9o2iEj+5IODdHXL
R9luwbk9V2OM0XmVaN5IpsauVgK7SeR4hdcxguLm0Hz7Bh9hzsyeTStSE0NH1hCe
Hd8ZyGx+0Gpqcq3+fxok+/Yra0oQchLJHDGHHpZ276W1eNtnlz/ynD8cTfC+lp2l
jUaNO9Nt85DMg/j1kdqWcGmAzTPU28t24PC0M3YUHgJjRpUhIrEdWwxSK1PlE563
dbWmajKUYWLMUFqwH9DRIg5RNYGIhw1FxUuYhCodAjin/OI246qwmrFtdvH+KBZE
cs04Gr9VBhYamhGYuZRolhL7NFY89Uxdmw+6O8qQ0DykwX08SnffkAQofGVtPnxG
h3MUzZJVUsdh5vVW6ZOFSY9sHK51k/S/9SSu6BhIWTuykFWBGwVRGpeLHZRXmgY8
CG7TltEaAdFK5aFSksVOppoHB/Cyhp7jVAtNVKeA7qLFc4nu0+2/Gk1tUL39bMuO
wfnEuHvuD+5FWeZcA4MDHzFDRtgAskV0uSgu38aRuxK3LlpjgyTB3cCYhcp1Hqh1
1+lsoLlP4SuWeEyxv9vWEQGmSasvCb+N2EeaL6coyqXhCpatxNiAgYF9Y9ja1fH5
EmYgBLrX61MGrLL3RPz4QBF9PKg8XLf/18NiXUQs9Y0Pzxrs13moHyvIGcztNIbj
KXOeVPRvdxbKFlxvJ+fiRHhwrxFm/zQbBhWbErwQYqKRRgN/jpuLRp4wLsXRfseY
XGR7iXDIt5LW7OJJ0LRbFMxNMacibGIWAicCo7tckRfFI92ob7dZH3e5wwDtNqrl
kMjhtEJSo6EhQHj3vospoQleXDsKtCAUZ8CH6gHgkYf+io15iHhaDI+KF/n9QgA1
dmgt9ypnyohAcm5g5CGgVsIyux6v0GLBtiT3OTwwZvBb6K1Dzt5V25lkzfOr4/mk
6M/BtXsxU2bsSbXFUtj3xYOpMVWjY2mTZtCjW+j/crWj0K8qGyb8I7l2yMbJIBxt
HZ5P24grMQoLBy/HnoWqhR55DRhwbVFX8dX+g3uBCAOL1djoLg4pphWbxxyUxRFj
X3r8mJB1oxidtaQ2U0FneOrJtVJQO6Y/vSO7tZcLHAD+9sR4DtqnX8N7meqA2p5s
DPH6v6OHKS3PRQLsTq1BwbnyHiNz3DFLNKGxqVTmDL++Yd70K8G+ltYb/N3rp5yB
OoBtXxzlE2MfvjPMfQpe1ydiRtI/hAzovpM0gepr1sm1q4XcWTv4KepUEbVzoGQ7
qMTNLwo7wEhqkhHWYTb3PaAmGqn6BkdfajjUO0LAwLwY/c1UierHGxmOSQGlkAxR
qyvuziR1GrvkyDF3AfO0wJ6qCftpm5y+HZD4qbM+YoWPrQ2O8V6Jv6WFfChwU7ul
m27gvpKx3DFy8GV/yiNlvX3BYPUPx79STYWnc1kulxet/4rJY3Nh2v0apPGJn3ti
EBjLEKNG+0M/jBZtfiGswuLf/FsnWQlLuJ2ssVIlFPqmbcyfsvQENEZzzpatNZhA
Mj31ydOX2H3IUsj77ri65jKiGWLjgV1Ps9TNmNbodkRBpM1bglL6IPh0VoeKrFBY
JS4Lq2gixqiJAORE9W/COl98wLGoiJLOwaF1eAZDhnaK/FYds4pFSuaAP8yYnOLD
33bbUdKWQSmW+EJ/A/FX7KN9K8cEErWbkeD9q8qAsQXuS2hhXOBC8W22zV/1fXvv
noMx4fjoGxUGREaM2JxXhtJASdc9sampKyc6cC+qi+CbsPkg4hjxg9bPaw79HBWR
POPkmKJfa8jg6zjY1xPpQje9owJ/tGjNDqUuyA6ZSrk87YdYY1dA1TR1JeHhvOhR
RlhJtU+5Adb3DTU22LXnkFngI7NUkOQ4KkiXmhEiXQHRTbY/++NrKlfEVhGD25W8
qMvHirzf7tiHDHuvguT8vwSt9PTiaTfr4txuqJ4ngFNCcpv9HivAwi0Ls8MHux1s
9jJ3YJ99zxKVEP34XL/DmlD+JX20U/SMDtvhrVOJMIJtTd8PLknmbbG4aMiAgE1L
7nH/1KdTfWikkY3bcjDVKvAETiUcIK1XyEM/TFipENRHjF+jVwoO/1vZUReGAmb5
PsLrmGJX00QeyouKoEOO727UTj75Sgryj8migavMjkbegmEqDWBsPKj/Hbk7QGN0
IEdKFer9Z7Pa/5A7Cb6kEf5rGlKZRUedrFVKkTgVLZ3i5ZBFcAuaBT3tx9tiSHYj
18T4oZdajbahXLXoZ1pgfCC1Lbo3aNJLyT93eUp5SvNm2nLA/Cl/H926ZXYt3mCa
V2xtFvVnye37sX+DhAjE2H3DNZmWHKSWEG5TnoNaYfyEFbaiGumLtBqfkDvqBn5b
HKgBVllgKIryQnBOW74knviNiVrKTWoyIPhEXqKakijash1TdXslNKqK2n1Bp43c
H1sLSewFFK2uKIJvG38QF86T3z+E2Ofgf3H1Fz/x5OcU6GiC2P9JW5mFXcBmMUs7
ftRwq9PXO2Zi2l/ejy3jyq8kbidYoRteOVIkjBEalYfKW4MW5dJyiGnPwfnAWtxE
qJ5hATaDy+b5np73G+CJM3IVPQRwJ+YT/S3HpwEHKVgV6HbHSLJoAJpddh1xHge5
8VFyQy0nYMg1C3M37Oo1FJeqFnSP0f6GjEdJ7q0RDZeuEu2XQeAqovWySPJRWzFM
3DvyL0BzO8PWltoiOj7FXF5ueckVsAiXSrLW8+jLtbYJ00NdQYghXzGR8tbWzBrO
PkVaaQgftPmzAjIgyBPYE9HKLaqcZu24rmPnp0VYLpD9bwwg379G/LExcnHpY14R
rBsNMf2qSUDfXIcscL3N+abaWF37Km0OXQ86siIyUR01X+G9BPGakEv0ahSLm9zZ
C6uun21rKdNTMKVWS5Z9UogCK5mqKJG/82qWb3GRb989JwV7XNfe6tZ0/6TwadCf
Mp9GQ/DgD4gEJ2nXFKpdDcO3rsLlC7ODOTjjAl9Grp5UJb1UcCYBBh4qkQ0Dl+d9
5OOuzhvQHvHxuHuWeVFQ12U2NVlqnw114QrJSbUdzqb8CMpZ+zCUw46YA5WW53zK
7Tcb2fdFrJElK9H57sOT0XEBT6BcuKO8sEpget4FWGbvvhTVTCNT6nycx4eUTJQg
ASV3u2WnQgptucCi3Al5SoKrtp276g1POi9lvzFLO9T6V2KODVaISKAJJ0S/uT6O
S99vbSGlvxnBSkUbe0E7qyrFw72GEl62/LSgUJugQpL544VX+3fVlIXp9SOJ8uuX
+LwjZrBX0c6uyE//sA0JH7t8ec15BJZAf7x+Wdd3LIHxE4J92h28jvX9yts0c5Zj
fHE+jseuEpISQEf0YAXA2dT77Ac4PX4dO4UjrCJ8Ea9B/tB01Codf0LxO8MU05TN
z83SnoDCRj+SYxjTnBZtb5/gl3cB3VLS8bufoZ6XaTZ8mXU7WLLqacE1koDQyfoB
/2nnsQu0fsje/+cnlNitpg==
`pragma protect end_protected
