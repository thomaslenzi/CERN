// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jw3SslIVTkUlRyHaaEMGk5Gmqc96fcR+8qYXafAHrcO6FhULtEZXZpPx50Rlc55O
6SjVEzBMIEEmyi8cnl1eWqSrl8Rs+UwC81efj7WAYyQ2X81fj7lg/3KX86g9VF4b
GcCmIQXUKoth4ITo0A51fYAZPOn09rPVPj1D5XvDv64=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16160)
6xSqZbYiX125mEW7i+LkUsUkyFUdNPiU8OWkqSP4o6OpnAA3zEBt+bKYYHS+Mfrd
OZSwqYUPti3zN/k4lG9IiqHuoFtL4oqyIeWVIEF7023VDKFDDrYfrxvMyL7bc6Hi
6/Df3j/1NSffsFtNM5byer++8ydw4mIwxA1kOo+kjJkpAgwQ12PDj4ziTimEWjV4
pScmZkMptEtE+76+jhSc6eqmlRO4qXOLR/ekswoawdM3TyKJabIv2bFmwKOnjRvZ
F2Vkz4W9RhPtNZqH5/A46zYgiKBHvSvMqcujltawiYPsHmRY3ioYYsxNwueSENty
at192PIj0I+TLwYFI0eO9Uv4Rc8PZnt1TlnfRYRdFf9FOj/VuqfzMlMdB2a56SCi
rGp99fAZ/2D/vTQdPlclCvczKbRE8IfZ7gCPt7g9NrN6LAegUSCA760JbyabzPr4
KYAdx2swHqo+hAq1QQzSo/TL6y++RoK5xRFYuRmAj647yBifsQ568FOxpPGg6o8p
oV45XCDN63mdiNTsSQu+IaEFfo+Os8dl96SaDr6b90dlwHF3MDOikW1GCSBxZf6u
SbLfQACBMZa1q8pdjcRQ+PJ1IO49yDHH2xI2ivNKhW/LVFBSqIRchYXd5uAw7DWK
fvcyFjpGZx0dTd+uTvSydmmNiOZswlw4FQt8IUnjv0EzWYXcybkhwR0AqrN3xKXd
fB4BcPAiAf2HgTElYVyd+sf7N8WuoL5grHPU7mqjKUX6auMV+BHXBx0cNRDFYdhL
1DtecjjXxnHJ8615aYsM5H4n1deeQC8A6v5Peb91eXqmw9/EALU8xm9bQVTEoSg+
+K8NuQfrA16JV2hQkuBtk9ZTySqcoYdCtpffeI388cEB0ytcHUNfiDBJ9hPlZ5YQ
G2rhB9yQgKiwu7PeaEDlOEVGPhZs7vKn1BsMdTs1UoDw24ea0CMzlBNmESwFeTld
8/O1bIDmnGWi9Obu7WhTzIaOxA8tXujed5ikxlw/NN/hNEXVZ2FzCKshQ2FCwu94
SQJwEQDp7kGldDMQwsh/aZxmZ3kGUytTJuca9Vd80EaUr+oQI09d1A3/zUezSEeX
WHbYsEuVttFen46LIGr/zaMwAG1avoHSQc8FfLBGxYXW2SxkO4wI2EHSD9nhhtP1
yBIFxoW+LlimoYwA8eUlk4FYQlBHwRdmMmY8ri5Cw1pXrOakjnSoCBL1tiLgDcRW
gAQ7GKSb6xB5JGifevUS90FIyOW3THalbIxrVJwJ/RlNRILqSVdfAQyURrhTrsqd
qR4YbquQoQf10QcIXi6iCeIckoEy920/yKh4En/KjlCA8r2gzr2U7CDdj4y7fos3
kja3IcKyHJqywwQhdXm2jDW28AEcBqb0XdZBBzkvcJ6tmzloLfFxL7YbVExmqDHe
7N/M6RJpygK+HWh0i+pZia6nkID89CmRR/fG6B6DzhD10pzFuSUOEs/RpNO2F/Mq
Znt4LRId/6xWzMzCvqZe2j+NfYRGtCy4TN+ueDASRM1kvVov3UgwUU5EQ+5nQ7zG
aZd9ERJh2ML+WnAiqI01UqEDUKb962ZGZdx0zwWhduEA084iUt/+tQaiYiLIdmrL
cq8q82vI2/0tU6O4KU0mkoJ5ppwZKgmRNw/JSxhjbAU+4D5QORKR8Ze/6eRDPUPL
02qPuYFPIL1k0dmXwof0CWnBRrMqiS0tlh0bIUPbGnpEg9SnBAtox36rkhIsLgjW
kz5t10Qk3eBQ86b2D6YMhWr1i8yRRiZZfbK5lrHkYK+UrbK9ybUPw6dTzpnaP87W
BGOiRnIzpdvibX//kHBmrJS6Og3tg+ozkbmCh7gJ0kVEBxXq9Tu1GGsU3iK+NDqx
pVjgKBm7mNfoXQPp/8UtSprZ7sAsJbWqfLjedDnui4AppY4vJSkyRfGqY1P9ZZ7n
ijVugjOVSeStapA8J1orjYvp6CtJbBleewfROxlV/VEAMsIE5FL8UAn08MZdQq6M
ZpJaIZgGSzv2bf8UzxF+CQd0C8WBjGjTCF3p16/5QHa3r6/I7N1mfRRAQ2EW6HGC
QDjky7vW6Z5ShgXMSpkRwT6xr6YCDgDGv8JZTCj1Ukxz2UktrBynUswsiGqAK8TN
5IgGvs7vL3MwKpTGnH7CURrlDKMvxFNpSA/zFE5zd9X+DviMArY8nzN1j0ak31hK
7kBV9hZEW5JNE9YSAcsM3KWuQqJmVdbMFwZha0w22REOICLusLf/dtd9CQn2tgXk
0GUSZw8ckgApEYfaQuo9BLE5JhgPOXINvn45sK6y/TrjbXzOlYp6qXW/xw31RhzD
iiOE0wqbUdnmBI3hLdTmcsR+Ff3tH8gzpEKk9u1paZoyr+Joc9fm7JM5WN/0R3XE
Gs1atkPTobRek+rFo028U65aLfbmWc9pQ0u22J73XWCoqh+ldynxQ0qGKEDtcmz1
4Ws/4cl5I2K5NSFciHchM4ArWeAJ6F1SdmDlXVPQwkVBfgSSAIYTSOMiZWZRMFoO
6QteKygOXl932bzndKCch9pYNLr+cfGUwefx2KpAW2N7HubEhuastn8cSAULJFpB
+Is/2YkRCPBa1NQxJaLJp9hGvMt2Axp+UJgC2BmqZOqaHDZ76iQYXZBFKtvFskE9
Ov5ikWTQnUqxaF2T3pNlvAYUI0QWg+ihhTZRaNAfub4P8VWGAacwtSDcqHzyNMQu
yoqdZHhpz9ygvdJlS/zNz5e8C8V5kB3uBpMczGCHl+4zg7GhNGymjm3Pd76YzlK1
sg6NzPBDw0dwWNb2GbgMV6XhThDP+79YCPP05sbNVRI0RZFiF2wGXF6jaFhE2EQK
KkwGoCyxkmCiRuJ+bNo91bqh8XonMqjxHs1comF8p6t9CCVVY8cbH6Y7zizMXZtM
Ki8hOsni1ltEN8OU6qSVED8hFPaXLaa2EeWxvzEWVqMkE5e6e6bhy1Xjh48u1ftD
WUWbo0KlAe/DWlafW0Iavy5thoopZTWp7YmEvJVJBLRUGxpRE06F3Dzlr5hZoVY9
8SpsnhueDtoftZX9U8foskLpol7ZYvzjdF8PxWf6JrCuQRreY0XYkqm39kMjLC1c
hCbvbBMGsIOrEV982KC1mbxNNKbL0MOj/NbUkHgI1nBD/o4onSUKCYaWyNbEgTLM
P0XhU2HWovtjXFNXNGzVDKpAlbe9+R9aJNW6tGmbwEnFtPvsbPxtRodlFoLfDzpy
zm66EW+K1eLxxHEL5T/OUKQuWHxa1sG41Tdvx5JHpPcSnwPNE/SiBDt2Xs6CVBmM
1OXjpmZEFZlrn8NJ7gzW0TC9FPUlxZFO5j+OW3BkEVrvWJ893E2voOiPFTfA02Jb
yW9uAFcTa4DsftSOdRGJS2Gj8DTaK/cI+FGAOonKBoosmCNneEZ6aoVyOFo22tLk
CaABhwuJ6ovP2Nl+zIWyUEmnTsjLEX2Qd6EXaMllDnUlLKPtHhoHbHEf/BzZK40y
+UABu0iZa/r/AGAJ2hfczyLGN4Z+Jt4En7YQmk1B+cXZkKiVAv7sJy44QQf+2t37
XplBKcMukrIaz1taJ5FB1dA8zPwb7IQ8mbOLIHDf1ggggiHzIi99/yJIUROFs7IB
ZgAGzP/rHMW8FyxGNlltUTndgub8ExYnQpSSjtU0IuPWdd9NHNy78Gm6o0Aov11M
M4WqIc0HaXFfN8d0xnZ1OIlwa1oLMPZRZTIRtDkMMIma7gEdVjw0OgcGNo4OFUjd
lzud+tyMyns4/DZyFpSQHcQUOOchIBmir6lWUiHuT3tG3AaHO+KjkjkCTjtr8vaQ
2caz1PYbLEBCvLlXfUeF5xxLGgRvCKs7xoA+LLCYGUm0l4x5hs/jHgakpbVlvjuy
4x107JyfKnYTBwzwihafywpM62rDClBArU3Jk8PjKxaYnLXTljP0KriXodr0DjUn
tJllB9kNITh8iKl5du1yVr0TDoOihAxzTIxLNEAA9JaEJmnqmOk6aUV+Lignu1O3
ea7SkxoVWCigmOQfePHNj484KzOOeHPmfWE6LFf/0x7JDItp35Q342AuuX4J0kRY
5giSHvLLTdgxzBaeqhHEY0+A/RlZrUhG6ambRRITNYcoSSYXa1w+Wf0iVFh3qhSL
qy0LTu35zB6lTSrO77WvVjlUXHasQudWuemf8mRY1tC/740imdDdpF1GCEH7OfRe
SUEyVUwlYXoAUwnzDIAy7tUigaqaG7CGGsjTMXMcxSIYM9h3AZHqZnBYpY/HoQFo
59n7K/VVEoyPos+iLC37qaFOiFwCLARI5o/lbrxNk+7ZZ/B25iE0uqsb7Y9XzU4G
L7XXCe5g3iFFDTplhR2iHDO0AdEFsAwkVWBcepX1y5PFU3ky/dYZStZq9Ions8fZ
jON9VlBFZC2YxoAc6BJYJ8zYEZH8nUeCY7qmn78uOvj4HdewTJVDn+E96PI6+8en
CbJl7dILuSShx/ieysq9JzJNcFrXwN0+zDgJ/g2RcB+0W1rBfS29gaBlU9litbll
yBxi2jyAJ3fjNkGfwN6oRYOPFlYQWlWDRPmaISzlttfpeUywlf2Qm3shSwxBN7Py
SYPb+lVE6x228biCetUnaRq9/yRkZPvx6PpxsU/b8LU/t/i8m7OQ3hPnWYZgSetZ
AJM9xs8/spgCNIK/8Cq9zDzE6uSQhrjmCm8PlVZX/FMyajBmNadK/l3dQvilmEDp
snO+O1OMI0DjvDNcNjZNrAS8pdx498KVr0pG4TnNxRvf/jIs241F4MmXHMU8gfDf
ODxi8ZCeDI1VQV+9/zC9XkcRrQSsTuxgfs0ECb4j9JQCPWVJ2VqBk7t14Qo4Qf96
erVRPlvcyr9YFb6d/qPDG91xHWNifUwZy0vUlhmJQTWOlQkwovxzauaR/dZduwUl
WDZ2C021BKuSajKkA4tZbBo+yurjClBnlJnTUzWtqPPtIjI/c3DDfkexThRzjArD
UFk8iRhG7Z5UklWGolT6h9WrQkVbJy6mm0eIZHesXce6zrglRvnzF8IxAr0AoZIL
/Ys5WGR+NBxOXeqHytWbHq7hkJBoJVsDI5eUis5VvN7yTNgv70qggceH7lbRY/k1
aFklgvR8gfTyVp+fK4nhw7VTVHH4nYuFySVnELyFmc7mzxXUn4pUOzBNaPUZVInb
M91SHbjausXIJi0snsDnExOshcH/fnjXZDJuHC16onAmZs9ZbbTs6yD7ETVdf2TC
7Elk12KFROVR9/Rq+jPGAqIhe7h/goa+l0TylJOzsUbmAAVuXzoiUvWgaBhE6jRe
42A+6zSmwUsNxiEREpDridbEJmVtibPxjM58CILuhKHf2fjyX+KTE1tBxCLuy+xo
n27o/fZT+oQAhKEjp+eIdMPKX4ryDXv7xVUyIrC8n0eLq/2LsYw/f3viIjE2ydKm
qBD+Og2tUwW9U+0FMstQDqWrEdeu05ECYBOygFJN/DeVnEVkDd68W14QjeGUCOkt
zivFueEeXXgRuknZXlRG/Nlos01acJylHDnqBSOYnke9QcT66MTVQKAVpZYHB0V3
tA6Dbegh/lRM8xPF04J/5rlj06emwh3f/r2sLXCv1Ls3o42mVun4S8TxfrL4D4Ej
/9ux2AYHXIw7aOz2QnTAfOjAaLluk+XFooyCArpzaLliGIqcymefCxdo83k1VQxe
tJNPSThNKga3rta4yHgPvALF2JwMiuEow/I0GJfo/c6bg5BeRMCNHvcPDH/gB8Sc
j5RPx41QX26Ldtqcnu0xqka/RbyDf/oPeFUc3orKsf03H7tJbcJa17n4Bc4mVgjH
irwcXyb2i8tu+iRGS0jW1fudM3PlPzM0AASZLQ/GojYncciFb9mMkj+pkEoEaTGu
eE6FVlLwXRIA+GPpzLSWfvUK8WiyqvTEb9bBDNaF1rvSlmeUHrAVnUaJ1R6HsFNl
4naBqPqPQh0slKHpYV/HTaOWQ2z5fUxb4LPY03O+nY7pWSSi6nXO/NcMPm74jzvN
fVVQnnEGPDdaA6xuH9kzjeIxgPXpBkf+zxUYeR/Eccabb03RhP0Rc7+//2Cd619M
YqEMCOplcDRk9O/Rq/K39fs9hR85e1Iu4QS24ukU+8wp6M/W+t8XnNtb6LXFpC6h
KkwWPQyPYnIYQ2JsFxKl0OrckKaUmW87la68ANWZcw1Wg8R5tGSMMvmmdBbcArr5
cuLkLyRofKdHmV9iJK8Jpa1zdyUXUlSDh3iihGkYUMw3sMo0abp4r08Ya+CxMYyB
YyPVxv7pGzJqi4e7SrtjgUbYyAJi8zUtmHQ9WWCP9aORaSLbBhDyVWtgAoysAfLD
7CY2yirB45ysaOSVmu/Ku5Dt9ur1NjHGhq+Gpm5jYI8e7jWq06fbOrgRT1jNhtIz
s9DnDKW1viAQEY5ZvPxTafphx/WM6yjl8D6/Bga+iwkkCm/iYYKSLA4wHPMqG0xA
G0KejSdK4r5/zPEjFHLie15FUE72lZTS7ysDcbHDLsdcqnOPKHDno1ERBi3zZ1j4
Im6XSiXVDViG2KEsdgKG2X586sBGd0MI0HA1U+vOReacRXM9g6kw3pmBgDpcOvTx
YiWABPPUF3ods+nMlLoTgJp9JBjqYK71cLP/8FMb6ck+BG2L6EsIXplyyILY5qP5
82AyaSUlLcuDXqCMmW7zKVaWYTYB4sy2wBYsT4t00fk5ErDQSp2nxlWrjVve2agi
KjzBkaQ9u3cZYC/Kzhdv+EU0mN8NzgRErDrmAGZ5TqmZh1hewTXN8CmcPyObt9y+
otctrk9Dqie3iRz0BcxLA8Y6gbZnELZW6KNFcj6zBDjZNuf0RO4hHe8z2S6cUP8B
+/C5U0Rc5bDkfAx7J/983P8NkqvlmK5N3l+WySgK2cJQ6Ox9seCFpes8ieb5Vd9n
N8UsTu4ZUMH9supTA+tKEJ7xLzEQNeeSHSy0jxSmTh9eBLxNWjwG8rmwrT2IoBY0
FAva4PK0duuqh8iyj8lb2Nh0I6kmURkYwFlQ7L1eDN8jNVHEnJUIdQKGE7q6sxwx
1CC0PFB9Q0sYPGJPFn9GbhuKaKhT3JrPeeAcI8FrC9Ym9pLVzDTe2OcLwfEazTtb
ZCByxaW6gbNOJSyTfCdLHLp6XrX18L1k77IOQjIaAGtDIq0Y+W65GMXocClq2XQr
fL0p+AyPEyPsXdLFRuN1XO4UD3RlrhZWBcymxH6Ug6ELPzwkJdvSUToDm+0LycXP
F/fWZedB81HTVi5+SkRIdsX9XxYxLsKw05fYu8ANhAPpKvC2XhxHyKy6Wbo8v4JP
ik71tfl1uIS9fYxJ5icrFmwo2PtHiNbqeppfw3yrxDOEyOpFBOqbcTkAlTmd3yfl
Y/N5p8fKAMGDNDsvpFdH4eDX5PIsyWOIgu75z8gqfrWKHV6YCgFeuDFT2OdTjae4
nI90m50B9H1V727UAfngkjPl39kr59M3h2fH6dHjV/tgPzwJuaVvklSEWfByeFLz
MwFJG3SbSJZY1lGctaSNcYo+TxcSJ2NIveMlO/lCEG826UU6S7CGx8aaIXa1TXhv
Ey0ZrEjRNbUoH0kVAPxqF8W0Ju+qmksLcGAEmZuKstDe6c9Aop0aoWK7mCkCvbFa
woqvIeUZin4BaUu4tAN6THRutHoBGwCV1KreT37DGzUZcbVsQ971N9zSgfAgxK6y
wXfSBRK4Bbu6kcSMuCGJVS07SgA8ZYEWbqqqBNr3MkvGEWURSPujJz+FIX/+Rthi
//GfCQAKkpLz8tGZTxkUebGs7WggsAm9KUq9+/rL1CkigXWIBCD7vNUDkL6LgZfh
eJeDXGBFVIjdnsYzI+hgt5eq1Tq+3Xv1igg8RZlTbFO8ebC8ZT47NYznYHUbWCru
XG5MRk7rSDB2uyHMpTov1DNunsfYmpyHfxn++M0I0pfMKjv9c6lYhv3bZugvrr19
BvG6CX7Eeot72kBnc92immUkmTPe6myzWBo2lHgbn1TS9mqv6JXkQ5YKfr37cAFu
OSOJM7lR8ZXK69tMIpQyiHdZOmdIQaZJqZH/scC2lGePG/kMWfCMGV/N+dp6bxAn
bKZoWyrU0Lcd9FCE/RqpmkvDJz3eKJCKYETmt8kMyX1b9F8QdSYkgXeEQ1W83opI
G68WC1deQAUArYmZorXy96hkbb3QoLwQ2UvoDBEQswtWhJd7HINUTdbYawlsmikE
QvTfmhiOB6NcjAnocnSAsjD/HHBnTiHX5uAoWQt3lJ4BM0nMSkCOV//+NnA+B0oJ
ARBeea45NCBqX/7I1hnqcEyRMVG+a5kdeACMn6o0qsF+cEHv+HEfd5443Gzlro7P
B1qyLt7SQxm8D7uSsB4ZKsC+QbkAOwFDBvI/7+iIe9m9ATust+KbI9fTdX6i2z5B
9BX8llymvWn+jJzMwcLtz1BgxyxTTTnWEv/Q0tNBUNxd+uBYgHOsX+n/Rt9eT1Tg
31if6W488Bs5i/H41xsVnJWbv1XL6Vmi+15UIcPulsoxZUK3e6JD3vK3G2gLVZqP
ySEW+qgxQjZ40r82f6rT8SMk0Z/Q43kIj5qFVJ02ssY+utH4cQHw+8Wz7HwRk5am
DSzbfDDpwDP1/ppmfV2Kx88uHpYDKjwe3P8e8eI8AdGeuUYmdmEFram2xlgR/gpN
gRIXLttao+xML24xaGkL2dUuC1lu9BuWG9QlrRIF/xtY89fPqLACepS2ak12prL+
9glBKZx9AqdkGtEzWcL2AfcLyLHAJrjTbHoEDvrrArUb0J5GBTxsUKyUUD0KxGaT
vmxvAaIomw6X0frSI+AWVPgjPD0c5XGAIl7u843lWVWRV44J/kzONZbIt2aEj3nV
f/eiX9ZSbEzxKbd3bR8F9GPDAiy19Q1A9Lv6knkTi1Nq2zNXsg3QpmVheLh3zKe0
53mu+QlxCz531fB0aqzJVRptMr7H30+r42Ga/yTNuI7X4JLCT7YJaSbZFT2Hl0VH
IoJ66vnRXEI915p2yIai70bxs8OqBoT+mKg0BgMbpjpIRoIdmzsiqpo3up54foAf
oystlgr2oLAArQD8i7K5onv8UYShh6qwbNjfwt7Hd7I1iRtEDNeFk321vr/lp+Uj
v82gUDnTmf2easv+DAWqW1obLtmXIdwE5tcYmEEpDFpvz3jo6NlDjtQxTEugXiL3
UmEwO7ZrX2kRxKMOFuAAayRMq5e5MP/Bw4Z1prOmXiQNMCykTLmN/vbvSqOM6qXA
HL59990HadvaC3pMuJmga72/QcO/omig+/79/9i6NXC0X71d1MlEJqXmitWTLR3G
Y0+n6vGHDKoTjkhKBCW0fdZcoSQA6eKScHcmpAHUKFtk+QMA/u0q8XZI1SgPLBC1
CinjGrgbYCBuy25OlsE3XrJhmO9kOMZ4zLvK9mNB9qmMAjRlj2rIdNAXxYpGIaIi
AK8ssAPDnmPR9MTL+NNds2OF+5By2Bgm8XyX+a3Ccef2E/+fHnN5RIwGe9DxvCJJ
MvHjxqZY2Gi4jcPfZkI9EidLlF3qiiCwU5qIw86vhFc+I5ZwhZA+UdCwzyHiAyes
QoS3OZU7N01BgQB6fJ9ND2DrOIP2uv5/ntxszFL0vIucph2u8xrT5DgN9+jWT0U0
Hk4y/JzBzolktBMC4aZ0yasQNCDqBoZ/BNwI+r1myCgSfbmMm8zfoF6gCUbRX5qJ
YqTPJ0CHDtvdb1F+nrqZLA55HuoSVmiEJmrs+I1mfaEPMfc5p3kEugFLZpbEngBc
GGpc6mNavAUmL630RP0MWtLWDnhZ+Up5zHyve5hzlqbIMVtkMmPDyag9LmPfvD7i
3kF4eRbR0zM3OblKdzn0QktbdUrWejPbVjJJL46aHPuy+twepIaHJ2j1CTY0Ye2i
H3IzCfq1HXYCOsPLpur7foisRu5A+Vu0TSNgFiaDKXxHslnBRTrvo1h8bj+n1vZf
RUAZ0jWmtHaGNdxr4se6eL6dtEGu2mULbfOQwcIuJ5+llwiijBFM+ABtk3AKg8Nh
GPwVVWkoTutHZyzUJ15+ehQLYY58y2RtPXhc5nSiwKUj/TsknWRWxTAXX/jpgPqr
PmiuY+3sjbiDFN7JusEd3nCqvscMWd+CsJofG8rWs5ElxblCxVmlA6Dzsbkg36ZH
WbgF8Dm4Vy9HMB+ATr75Ho6pX14mI7pq2HZ4BfrFbMzDK068LjtFn7lDMfj9ueHn
7VCVrHPLgxAiz2eHpIx7inVxi15xddTJLZoKvI7bLMMiAIiW7U2gBAWLOiVDEA8p
d9Yk6Po0NJPrvv0YVdHd4W9VDqpzIjGH932kWfefNr8K8Kx2qWFNDQREXBCpSpC9
bnOrml333tyqa9C+rtOJOu1OrSAT3MqIn/N0sEsunLEgdNXiuQodMkfmovw7FZ/G
jZTO9bHVmROVXYB12AwDStMyaUa8qWl0S6va98Bf/zBHzb/QQDzZun852U7reGkY
jhaM/H+1BUHPu8bJ8XAs0fUyJHfjr1Vq4Bg5AlHEEqlEBx3fBXjgWTMJ0U94KhYG
ybaOPHpm05zdCMzpBkebdit8tXvS7ggYuGBv4JPCaswPLzPZR/kyxLou4L4zRgDm
p9ijNa0u0HuOjyKkvx5lwoP2GWtqPZGwQ5uvZ7P1qV2VV3Av/yBAEw9iSiFr5NXp
T0ffvLNIRXpNnn8XLS6snz8MwDblRQLYEejBcHT6USzVEDwGIkLXyfef92DEj4lt
orAbFQnQPH+3+OJo+VPza71hIt4AJodKvyqKD1GaJ3DvKQ2Zda9gIWZCDAC6M2j8
pY4je4e2+bhLPMksg9uz+nmdTYWh2gxDaLr7+N2rcTUxsVGXDz78kbPJeFaDhQ4q
aPgCyNW340vsrq0bFS+N2oXbK+nEZfRqTQ51E4BSaumoh/KbZZXTXY216cXKgOqU
N2MDkpYTxCx/EpBM9yxfD70TteZiKj1rU2hdD8d44x/l35zsG4jUvwMjvrL8SiNI
ASWYJtHq/6UuOSSXZ92Qwx1deAM+w1QVmWD6Zvxm8vmkB3GUusFpl3O2gchgwf6K
CsV9n1m2zrwcmtQB8f4FymRcccq68MPcsQ2OIBsQ/5UWNGvvgymyluP2qmbog98M
TORo4KHIksB37OzOjokvcGxt6jRWK5C9LQqJAVOGUMa10J1SiHWrR1NGvCds7RCc
yfyAdOxgmHZYF6qER4+kOjG1CLrCdB+1rY88rUkFwOsmmoPgeEyx1OhjVkaqvwhX
hPMKTQhTI9MI6mNcyPjR25Y89SNVIXLKaHI7xHAQP3YJD7sQdNT5h70rkgWnkQNb
rLTxOMTVpiuOK1l+ckrpH5WMlSxanXRKSNPHDYA0hjilopKal98aXpCNnWpKusjP
QkYooFd84JhHApvxPl3tni4P/tiG5QayrM6omszUZjQjTM0RGwLrM75CjLFQK9qa
zAHd5ry+B6HCx92CiyZhgDGz/4Dn2Y3ZjPV0KjlegK1mUVKCGKRefNqC2b8pm1Lf
8OwJlF2LXDv8i4gB93lWwNzKTRUkFmdzkTD0UIgun97INO7RtpZaT9JV52jnDdqG
k33+o15TrHZpIMD/kIuMz9H7LUlBsYYvhRCi5kzhALkaqY/48lqUyoJD4pOsguHm
rL6UOCuiAPNdrfxRd3dfC+506hETbUmyrXmt33D2LfosQNtzJc2Oo8AR8CqYJFaK
rELPBIF9KWqaUFGnkA5Ut6VMEoHgNZXCXWQBcpUdhqJC71GDv6f9Tya5iisbtAAN
PrKYit+NCEPvu7ci4yEv6Ez3U7HkYvtm4KjzkaIvLhqs421T6EWfAauruW9WndL2
ImBScBA4cE9RWEHu+tqwSgtKc6JFhuKnav7mpT9BtZOzOSTYxIPqFsKdrA/ZiyzE
GNf/7ePNM8ZKXxLD490sQA5f+dobwd5o1NhCzkkuIAQ0J3YDtcMXrX2fNvxoE+Bz
DSoWC0/eaicCfAlousoZdQRFJm4K5W0yYkMZ1Zlm6RVhQ4luaJDN07KXbYsxBG70
etOW4e0nyat805fA7Oqr/4OfJBRJmpj9nvlFv4Vin74i4GB3DLHZ+wJ7G66o+krj
2GuPI+j0O9/L3oO/4q7c9L+EP3ZHqHOC7qXSIjFoLkWGn6Eb2Aj+bHYIENxP1h1L
Y5GiUEIAWg6jgmybIlOOKVVpeJIi/mJzC4Rfw/LQeQZznaVVaF7rXVVBNev2kYyK
vE33nu78U3G7KLEFMNuqGYHsPNp8a4bM1cG7R2JdjpeL4RQmS5L8YUK0ehErDg15
lL6Qcz4trcxIL5Fq8nYrFSAYVjybEZttTAReUV3UQruT6ws9CJNtBRH+4HSyvB7z
FB4odduPpLOwZOyj8DyaDDmZItXNVXg1FXGGuk44g3H6UP1gyKtNBpdkNYQiFxVf
/1wewRAcEGbYHXKXgu/n5ethoq+L2sBHQ5y2ofnXlfqQowX+fzRcPjgShTPTk3jU
VzNmmeT9V4O1V+lkXYNY/IiR5rfKRbVzX5LY9W6vGWV0Lc19MksbDjuRaNhD+jYD
kOrMRcrF/L7188MMxgLqFmZhQdvpq0rk6H76IZhNhr5ZM66LOXY7xWh+89sgDzhg
ikmR3gHt0bL5dmW3gdxC/hw4IQ/EUiR1daQ/cJeL9W5UqqP/cJfMk9A4NM4tlcx1
ow2bk5l8wIBc1mvmp8CatltJyHQbD8tiPcdf6b+lPUdYgcm4ZhF/PVxfq9+ijmcR
dc8TdezvH+EI+5C/aGKFfbBnx2Cj/DBlz4Od9prjNZanVa5Kd+oVEcedEkwq6BGA
jfWc8Xd8J6I2c43rXN9bGitzO52BrV+iTeKAhGMS9s7nFTXiZWH5mCAGCXR+MOGh
Qi2ntLKDe+pA9SCs9g8DVRlc2JOVbJpSTyu6ZHXFz3AkSbyJZnZe+GsFuTm4NiuQ
XXdOeSspV/baHFWYrDIJ5MuOYodxs2nc7uauKa9t3/bXxvuZPngAGh+GG+D+5AA+
+qOok8U1RTLok8ikGQ9La+Z/T8kAcYte3fFnP0WocMQDv7xjIDjJu43flGgbVz+7
/Wdf6/KRdYWexiX9YM1EfIL6NS4w9QSQhw48jvpKn5sbLfimtQOOC2EzX6ZWI23k
8MqlIZqwks8XB3MK3NkfVRSglnyc5nC64TvQcU7chTI/Q2tNamIWGsDTrX8PkwFx
b1fjhPetPx83ABNh0e1EMQg1Z6fl8/555CbHpwEaNhYdrofn3rp6Dhj4oO/gxwVF
Flj8VwN087rVYndWQ5mLivJt36fAa1gKjgyHu64Vl2p51oa1EkTmK/NbLxinFYVF
xxibUmDBMIXABatBv7BqhPlWUprmdgTBYSrkoRl/Dhn8ztKJ0DQVO94vKbq5UWwo
BgzEuBA0FIF+QRn4FE0MNyBw4vPK654IfvJCMEoDtNfNrXdsBoJGSJGOBvnHOxDz
LcABhAqZBKwmUExKRa45N6UH+2WPNR/3jfsaa0SAT48YeA5QgJ8/nJJ9dZTFmOv9
E1ezpnVXujzntxKkXUSXKSJj0CjStsXQFOoR9fvbVK7QK5iehtYuzo4JcFmMFX+9
SwHaNEY9HcB7XsKaIonZsh2oLWplpD4Pu2/VI9/KD8u1RnheIRWzst2W8dH3FRcS
XcVYpXrYdDGOeAR+eh8vwCKCiESkRUUmCd3hu7l7ByU8CqvqmmgNhYkgMowu1B4t
4zhe4nrge0mIgA/zEl43CyZ8UOlSeucOTwmeflFt/BhcMYQuvgZpB418DtSRXtVq
iTBIZPM5XRibGA27nmuZv2tYa28RgCSy1X222BgnI3MlI5r9fzzLHrP++yTaLHDW
RpiiDItAZwk45zBaPm4KJ1Mg0m/6jLo8WHDV0nIg3SxkGMSiOGyoZNdzFb6yxsS0
U/Ck0LUVVgUKQ2/l9xztJYiFZktLzvXfJA4H42Xrzl8OCRE4OyPR8rmLjULsfJ+M
V+t/YpwCn81YvS2h1HbMDv31USu7fNzipd0x0g//gWaW/pw41Ktn+YHaIFxfkbO9
/+MIJZ5ayDzTF4xH3uYYeVsDqvxnrI+gWf4Z5r4JXvF4Top1kg9bjonHFljEGLS7
9ljw/eHidA0oNisVgugZ6BH5ATiot/KhhV3Y/ntk3gkJdyiQgd7723+weyahj8pH
jJOU+qEXqsSkmtFYX13DEPE6VoARbMCPLlnOYZAH4HCDZzFb+hW8/MMrLCj2voZ5
A7rah/kPa8pVcKR+jZz7fYKnuY6ma23AtHoSXZW2rs+TZMjfL8fPLwLgd7PmQO56
KK0pybArFMlpQb9itnGzuiNL01ZHu+ZnIPokXOhAMvyKrsNfs6i7iNIi7lO9nEIu
kcyT7/bzuW2qC3sxBdnu8IOMR4h6p4PliLCQ4MgncJqBkCkkEV/41hT7rOsCdD4r
iH3swesar7qOhizKO+XBaMSbHNnLpqJctXBYI7ozmmCc0dTn0oluYBBWQH2Ajp7c
HO4aMevnoBXYl1lY+92GgLF6PIXoLtXmZtbjxqdUg1Dt1e5/TPj65z0kF39b/yp6
AIySKU0zm5KtrK7E3M0D2tWB+h7JZ8L4xbCh/eYMdEMk92puuzvkPcBDmw6daebc
DLLUz/F5tS8J22EL1l7qS1ZwTS4T/RoapoBNkTpWNIyo/+V7mFkVLV+2w8ilfzVc
UIXQK1E6ZtVD6AZkqgr64COBvh8vko7f/db4RCabfug8SS2PjcjN0CyeAuYHQsoB
ggdiiQB9Hxtp4hPFtNEmuZB0PlfhnDbDy53UKaGBr3nweo5jgQOQroNlRQFa1xTZ
12IDaa5ec3IfLFZoWoYENhtTTmaz9oco72IBldnN+WakijxoEObl2CX8MAvaih9M
TdjSHrRXF5w39za9k8OHfGlhyjVdTChQfKrML41WtLuMDWWbJ2l4YhSJyj6kuyMf
dE7yiFuAauQ6SFJrsC6w+0BrnP4IGmw+f2XGoWSwlV8eSdrPlpCEFKT269OniA80
6Yv2+TkuTHNeY5qDOffbN+Rh8GbIbw3Dw/LaMN3AVzn87BE22QGiJWW4+Jnazyuo
UvfISscD/lUdK/Uy6ODhZT2FBOnmMWTcdCKGgeIvgxM9W2p7qtZNp5V5a+QSf1Vk
Ickxg2RvJXad/37ApHaxEO33mAjmITRJK18UkfZUBPCdmD0+fzsoA3JwXM9eF+Pe
d95yBkN3oGYrmGlbgbpjez/4eHzdJwAWhIUY9emMEI+6FqAhAHQ/Fz7iWFulTnaw
hKSW9iXhSmv61upLbc2kqlFOuI5AReaW0Ooe+QzjF0hAm4xqfAIheJRHDakQbGPG
kTULl3s+QofppQlst4jg32ipO31XcukO9XpO35GsZCYcqZ0scAwNOxjUqPRFdqG8
bRdEP+iZjSfQ0K3ezj86rUJP5G5Zzg8hTkSSlBbK0YB67dEtyRwKmhQE1CUFEAqw
rS36O1XOAEoWuDUbTwGdcho80bvbWsyI1tFc2CIZeAna/xFF7PENNUL17eGlOkDN
0PVyIpvEnFooOE1bXuFL0AgN2Eaywo7ii4bY7sC1S6rPxHZm5Nx1nWicW+OxxvGU
HQFJSp4xG/YgEaRP60PJcaRcDoeGn7iQyfx2JXGoCitOy+GfN+C3CWiIDtRyC5Ku
rqstujkw4HtIf8DHrYDsmCMXfKGdsxQbjOBrJzJykS/KidEwHZh9keKcpbdHimMF
PzQJj/r3gyUC7ZHnaESr6JnCDdehIkbIXKDPUwr6t/Phres28DC25KMhVfUCL5Uu
Lqvq2g51X0TxI9peMRcYfVHKWNQVCIm88TK9kx7+omMJvccrE6cFQ3EiGUE0XLlv
xlRm1XMImU9uwO5R3jT0bxfkIiV4BABmYq3UXhXymqE8AHusBlYjq0kSvUAHruGW
t6OxUbq5aMAbUU3HVp4evssg6JoI4z0zX6WMx495RD7B9Gma3wE8ekwuX1L18gFG
Wor+SBoZGCw+KIBmE8pV07V4yHa+GFkJAXLmMj8kwIJ0sl8HLaBc6fj4e2R3lvcu
TbM9l/b5/OmPAJ2DoYHMNZTLbQrQ/hFyxeLanUKrE+/c0tN+gsxJBoJiH5odQlLf
BL0AAy3cVbUwXtvBj3srk6Qbs3GahvLI1MeFIkNdvNmAzg6w7+nkCbP7M1JF/Xsd
vAbumMkBBB/zYZ0u75fs8FKu59QshIorWCrOoV5PcB4uv+wsMDunx1X/hK9QGfDH
7ieO8xRPf164Jlx7GrJVhNzoO9aq8WX6E0Ut1XxSzxvTMAB5cV3zA4zvccWsgz0E
qFDV6r+Azg35N+pz1l2ch5c05UOs1DqOIi3/KUrXXzV7cn0qNX5htSBaiszIPWxW
AoGKZ6699dJRDLXgr79noKf6DhavCXjE/7R62wbGSy9iByWiMrZ7Vn/g726QC1vj
ZuZF5qb0yoDt8tBAbXyVJ6/kcYzl2CACktfLlM9XU95J5zT7gt1C2En8FC6xlMP8
2MYP6jVo7tTuACY2ntGn/VXOsi8t7rV+7rYeFWEL+YP4BmB+tZO6Biv5hEiSWb4m
xGpCCcFulIi7PzjN2FdaF109YwkHDgQFB6jE8G+IJEGcuaIXbgtNpWSaK+mfeW+Q
k9HhSV6c/54cuPhenJKsyqXVYzm6jp41YXhl6+9I/qwaAba+ifZyvN7kDNoLuDP1
9ksZzpF+nB7g1fnelbZbv0Cv4r8YtDGuftxr+Xf1gnFGQlhy/YR9RpLXuY0cLoqo
DsVS8lrukd4D7wosJXEeRpbZDiexhthMaqm7XB6z/khzF/i5Zf4ZLK12h7jHzaPo
PgbzFdESfF15bl15Zx0mcxdpzpOIvwJLT7G2UNWsfj96V83G5NUefX5EcpjKdZEa
JRZtiz86Vrwqx6OMjAjp9tWVLBdCVOqO4flHMHZEFHRsVZIx9x3T5jSPhT4bE7q2
BuQ+oYEDosDkrKichomT2CLMClDEA+FzRqSNUshaWo7fRqOxR45OwVhgtvlTiVDp
FKej88bJmGmZTnO9cidGdAbcTcxBbG9MaI8xLc0qiDnTbR+bPoZG0LskS0BvDhlp
fis7T+jsIG3LN5BdYLSDDAvxWvVMq7YCxA4R5JnNVCkUwVg4I4a6A76btvgze2qn
if84C1t/fQT6Gl+/xO5hsUrbtzibd1F2IinSLU6ZHG6YwD2B+/42gzTmu3izOeOR
5IAcmzxOB5IxzX5DR8suS9VdfQ5E1vIvYIzFgKcQ9+0qCjbYy5gSGAxLQSt0ixCn
2MHz8fSV2AK9lPfnOYf5WneBtIMOtKWZ67BmeoB8jxJ4YQX/iFQjQCL9GJ+4w/Pd
P5EKOg2L4kPtaCqcCyqZ1xJr9/+/q/y9PcbjrfFK8Oqhn0Qf3wQ6huEEe9qtb6PU
0AZvNtbeiub7Wx4TdPJHXEpO93IxIhbiZVHProDO6wz3UY3OehEkkoyZBkLXzbak
/gJSmxRLiJMFBfQbRBzXqpmte9OIT5pYA7LUC2vVAFDSPXdhw/0QNqsWuqSKPr6k
YKy1CqmcsuSf1Axs7oxT7fUarvV8EqzNXOdzbtUjnpo/IOgZ/PhZdsACdr8SQID4
75BqOwqliNv5whOdtg1bXyC6cpeeU88DPjf4JRaxCZSbzhwNalMQhC1mxTsHBZbJ
+cidDGpW2QNsckFFJylG1vYwmxdZva337Ot+LauLsfTRFoOuOAQVDlv27IB13Qvq
DdJAzEzgg7mhlFsX+G+qbxNOXkUvx8D7eP5okydWQbYYsIpfw0R1R/CEZA1BhQAA
T7g3aP3qfZJsF9GituVBCb2Wfk0E9+HnSLp8IQDMhp7TUm1OQSiG4XWgjBFqj6Y5
q2kwUks1ra8nTlWoMQXaM1rSjACANOiBmJP8q0AN396ivnQxE1F0aqdEJxBlg0Gb
yaTBVkhSGUJF/+tv8n/n2ESaHvUE+d3TAgbq6AHSpVSqNpXDZelpTXIpdcR6R2KL
LnDABI24uuxCVcmVH18giQnhDDW/F8ATwZMVN3Qgc2jUJ/WThu5gl5U3zoIwqyYe
Thp1nzbTRy2jcr8oK/QQWWulzF0oYq2aG4OaGDv2VompEu/p+xkRGmQuOj9KQRSd
5leYm7xluzO12VyAFSYeSAdttvMbYW6oPD065g8uMCHjOGxIyVw8iUE/iq1VlCrk
CRZFtEfyAB5aRSs1pjmiuWY9Zqs4T+RIs79GF8HyrSBfqNIUIWCYH362hej75va5
oOf+UBinhXcXs1BpT656zwLmNybmePVBXmko6tZ3gwYiCZwYEZg4E7JMNiarFxY2
Wk3UwDD04SU83CuyESDB5bIAFaedhLE+SjmTHRhKVOl2dJ0fc4CREGY4LOyesica
Tq8EI3x0qQYKTh+RxtJUD6xnoEgfRa5KizUg6lA5kYQIkRSi39XipZ+EIXrOZU57
yKqD+/s6it3Q+M4rB111FJPNTUTnRUDkcul2OtgggmENjph3axMLiazomYqfjgmM
2ITF8IiX+zVfPqxJCQvX7K0hPfRx8eo0d++COzo0gXe3+N+na9IJYBlVQRVqU3Ou
Z7ulasEu3/ZtK8G3aJDeXWE8tmnO07JTxSJVB3d/WiG+yaJzejzvSOVgleHPw19m
k29CCJgLAUhQvvhgtH2ItFcY5C9msTR7UWNq9LuNNh1TgE5NBWZExj+osJmoDExT
RypKDsQPUTKYCQ57VyQ7pvpSjiEU246ujhF9xdyClcsYHL90dzojJc8nmxnAGx+O
h2d0PS6MmdpwxMy8wFAiBS2+z506UqKbOkOtNAdwG9ehAaQmvtIpM3K0xO05PBWT
Eca4KTxCzc6HDOn04tiqE00nTa/5Mt6AFK5JZax/Oo8+AwOUkp66ZPc3T7qQo4nK
SGy4mFAzdrfxE18w8Vp8zhhIWmwjJf9nm245nVrtquucDL0cAdOFZ0idVjbH1FFW
FlLPdcoPislVmW19DBKafTfHUvEnAO3wDpIfO92gDjSrOLhIdLE052sdNFnaMmzT
JYAM7jJ3v+JIFyv29aGLJEVurD/l0K9OKBk7FvudtcR6ldBqvohb10XgqgDim1Zq
QvZXLVAnCWnlVZ97R91zRWidspzvS5nTZpfyh+jscEGXd825ZgVUsrWMKQKVUTq4
cuBzm6DpsDThcnCV2PQMUm5o2B0zQjPFmWfOrGYK9XWaCkWbrhZGA5C2S0k5plIQ
U83peJvyXnF9U6bp5MM89r1yL07TcO56cF7U+tP0P24tfvydy/8+28vC1xlvaYJ8
LYi8s8KMWLaYXWBcWjcZ7hbUrAE9hmetxt2lJDRfetVCCzByFKYLicKaZj3gItS4
/+NVCDXRsYz4VA/j5kCaXOE1kx8mRAPB3ps1nXzuAAPuwglZ/YooEPXjuvkNB1yg
UrXXiCYhMdpGOicBhC9N0Q7bP0eJ0tLZwygCnImB4l7gd/7ugj2+N/LYHLS+5cNF
CMR5OXIPh8TB4h9URTBNJFYJiIXQX5ohmaBFTmG/hVrK9JjJj5mME9ZoaSswsbYG
FGW+YjcGQH+k9TZkZSfBOe2ll+Dz2FhPO+wrEH6UsOQNVYzcJ7m6EKsDwmBA7zCk
zH9v5tD95ZmUTivU0kgFCmAMjxMuFIAmNSZkGTsS2i3pz8AhXuMgf9CYPmctAQ4X
50CnUeK371EKkLa9QuIlVxDnMVPKGvfVNAcLVVc/nrz3x4ceQ3g2aju5ClIw7eQE
kVvENdQOyIWRAhg/CLwDv3DgBEaNwYlK2zRLua6J90XX8NDI0WNyrwEMs6qZ5Jrq
Nm4SJepTLmLG6S2YkXbD8FoPikjT5k/xmpAkMnxL9LyOYgn0ggYPV+xB9yO9Mkt3
Z9nF3wZzkG+mhgiBCGMqK+lLuye0plGshK5NCNGVUv4DZZqyGBuUjqHPCzyVPuac
+MrLaDiYBFqeiawdUBJUj9kOW1m/WbSj7b5U8LuXt9mA2P/MbPJ466H8Wzktx16a
S9oXIubgrNhvkJUwTGDb7Ki4ThMrQGkf2r6DOo1MwZf93yn/632xn0BaXNTiJ1u3
HmVIaEswyIZAvbGLbJY7PQkw2fgfbKYwTexrXH3zw0qfKxa7bvBr6kDlbAzMWqnQ
pOngtBLIXt9mlyjVifBB1H17uEUUvQKz/OHAMRMQmFCvYo6AsMoGjDyym0FRbaVA
KAESTFN5DsPTx+ZMOLSHsEsUponb9BODRh1+KJxSB6zZX3o3hM1KZNL7UQ4klxsy
iFGoM1bq+mitnBrRfu7IPQM1u9Bs1ZHJFvSUKuenlsJ21IkuT1Cjdfd0rllv/IPA
Fj/SkAAAu7YuCSkzXNJfcrgt9QnCFthzHXMDzu7eaFhVHT8IZclf9mPT6cEY9H0M
DF3q3fpFoTuP3bKRnLARufjsvkhe5sWQPFobvOlg0VmS7MbZUJQTJmeA4U6CN21T
FVkXRIJjdj+6/xA9eu2QPofC+KPWkmmY/UGOXCnVaAZq6EJPXaeeQWprsfD2p4ly
uyi7Mwf+4INRHVuQdvpsbgXYk/E0Gj25yWlf6wQNDZPn1NZVq1A8xP59QySLUP0k
4i6RKvUZTqgXvM6R6hUJ8n6lS78QxFU36U9EM0d2SnLg6u/VelZn5A6sz6n6OkTw
0XrujYYIbscdtXTAc4p3CUz++o6qPDaXU+y9ftyeEffOYezKnCtriiVFk/OZzSAF
s8jbiwYpjURePNr054JZ8emWlCW/3/FxEYPeW2+d0EvYyCMo0NaG1iZRFIKJZoE2
eP7XVg7S0zHra0olUN7j+6FoalPVtxIEA5v7qXyCR3qw/IlF7cCA2NCdPrCURYKC
iVxLGsSykOlGzHtOyC35nTOhFDwI+fE+ILTosxqbs+fEQ2KZdfCK3/a0lBjSM2i9
21CQXlenfQLyeYdlKosdRB0uErW0ht8J2BFlve1M7f4nhsz8+LOnkAxAHMzylyHG
tl8fALgCYm5kIoIj4EJPKzuO8POb9T0mssZc/LMpwzJLotEI7uCVdeaBGpOtjVtF
4Ya2rY5EgAKqYaoaEXcYz4TJzeDezOoKGygwxuSLqQPvu0Za7RQH463mNVlke+AU
sDBxRptJHAyl5980Esw9LRnfREl8EnP9D61M/eg9NjT9iGmuEGqa1fd+JBnjzF6K
rZbBta/UZtAi9CZq76V7TM8h4BHRcurr4iFRFKZk1XWGsoVIvQ4My9s9Kz9VLJ5C
bxIj4Q7xA0GKqlcfEPT5QFEqZz6vRldip0RoE3kpvKY6In0/XDHRJl1tVCjCzD2X
ffU1T2AEDYq3T40R0N+NIR6QvGvtb6mYUawPqVywdCXoWsM7wUQpw8Vyda5YKBhr
H04/mRuSyIwl/cJayQx2Jvxkr8eDTkTZ+Ac+lHWPs38WLTp2/ceVb/3KtL1cCYWR
SUafr3Dbr4pVVn7aFTjnneRqndhgZe+GrrFXR5zdj0tkjcwhYJMuh0om+vZdwTRy
iQGGnby6BeL2pT/txGVEC7fqfdwrVSoKgs4JzeOMYTu6BX+X4e/VWAsSpeU//TPJ
6asvV9XmqNU0bqz1GSGgOyNJCqtPgXxMFj9VCdKNH1NkTBEuQ27ZzUG39WcI7R5j
AARx2vQr3K76yV0/LbmzsPHhNATQJQXZ/2ZLbaQ1iZwCYRsIuoXNXS1ge/gi3Kgh
m4flMgOtf6U6NzUkn2JJNmspOETwFPDxPqnCKp5hZx3t7NxDg5n+QSINruFK4azV
QfMZKdihYZhEolw1oJbgE2W+rvJOBNWYZqJo9Hnxido=
`pragma protect end_protected
