// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MXmRFyZdd21ExU1GYy4IFQDJYu2tPcHYOY+MVd9P0ITtRjy+mQKuXhSM4V/ZEj4R
oDJdXxmqZ6JOhoC/GzhvTR4cQsgetCov2TSlDWnUt9D81uhqR+SZfvJr+zf93gSK
uXa43au036UEodzD9b7C+RG3yCGPIHI1kCET9TbcnvU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32816)
PujsahlH5Gn5U0oMzrcxwZ8sT0zNe8+XeT5hYkRHE2doc2UAARbRcXuWEmeftqVJ
T6SIG4YWVBCTFhHuF9g0yGRG1H0CQNtNxYFkkJTePSArTsjFZh8O4ZT7aNgEKXef
od+L8GMNDEsAJO+HM9LMT+t+GamVqTVpHDBqjKHmXlOGbB8bssW8pk0GN4XWOL09
hVd25lrnSDhg8G6p3FAtpprS/4cGZoN7FQS76ZqyvvS8PFdQScuBT0SwJmK3eaLi
qXTEMhS/eB173DeybzGNev1anSAZxdZT0QAhulC4++j/gGAcJZnAQ4h4h0AYdDkI
d7ilW6zbFz4dcPPwitZYFoQbpv+AYyllIdsZ70NW+M2sN/Nl0faaWOjUWA5Nc45B
auZAopN45ltOMldvdz0T6GmrOP4K83wKqrwL93DiWaY9hVlVaqo0vDcr0n2rvLIG
BHsptQZpjSJ17W3n+eU2n5Bl3zySnNUs9lwpLkyMsN+ZyLSR3bFUruWp1SxaxA5l
0M5nFZkTRNubpz1/F5SmnaH0k4nSvINBg0lp9fYGMSHVHTciLl+kO70Qg6DowVGP
mvIVvLbHhe+Jam0Rg4gCRyIZvSt0U1nSY1vsZPWoXTO7xYRMG1r3dvxQymv54Kaz
s0+ttylVOIq6ZZ20wHc23t+EgZBC4siV9WzngATsZpCCeMvVLubNOR2TD0n79gYR
B9cE+Oxs/QkQ+v5oHdAbHCQKAl6Q2AyaBqDCsBLb037XfbIY1Zsg98BhejhZtmMx
dUWVX/BR1U2pjgxrWwGYCUs4cz9OK970e0pyjVexq4xFJc0+Ozn2F/YIlLRuxgAN
2G8XdwYXQ35B/4WDsuzA4qs1qj/8YH/UslJp80ZhbNz7QDxXhFI38fqbJK6ASy/s
FwfxCn3W61e+6vlcZQKeBxtZEc7pwVBXhSpxzd6RRxyzLNIktTsR5c++G3q6C8qW
MYdC6y2+2kZmWO4GGFtJ4NPhLUrg147A9UIKRd3A9VQ7s/We4sSe7QECd49EA4Tm
uiBv5dbG8LJBNdtHLSFQEIsb881nj6zyCzx7OHatl38x/PRcraoPeXVQfZ7kAmAm
tV7PS/ao8JzFh9VwC3NALFNbyqdjY+6XRH4hvVStaeWnVYIpfUO9YIYD7axqwGTJ
DHW+Vmls9UhLaVJ410B3oM0xhbVX3IttqgH3Wg5ks64sZNdu65Ku4J2UFlL8YTfU
CQ7vCREs+x2EFxy1VtVXviCMZk10qytZBJ/7SOtghzZbw+bqyy5hlY71QGOBM1Mo
U6PX64tF7FcQp6F1+IqVJlnG7gOpiV+iT24PDqpFXzj2kZH0QdGT26md77nLHHVw
bhXkavL7CE2SzKWoGZfFjRxxg3Y6GHQ9CtbKXa3QISLFu7igrSxe04ZYGz77xdoL
i81F2hmGEySMSfeLAYbC8AKz3o2tSkZh3Y79iB9bhZz9lAZ94FS5OK8WeWPz9vQc
OQpHoOovKhB+1GqhuR5PrxKj+uE9U725Y3qlYPn0ta+lo/lZbh+etusQpD20zTft
fwEtENi9p6UVRcKxEvPxE/b/s5JrY51j2uNteSGISTVaJUPSCXotxzh00wZEIwFG
dVeeOg198kDqGyjppcnU4QGW8lS7llA0aHC6oP9p65xdnKyxTbMVtcyv3W0NqtL5
FAO56kwFEanMulHY6boQqYUWc3jJNrJzt5SDgAOWS4ZGq0g20YVA9hbUMtueUrM7
iDcT7a7avnmm6qw25U7CIQLub4KtKADsdjItkDCg+sGH27n7Ccnpdxa8RBOtMvNP
PQvsBA1ZVJG+FqisO6j/LkEznhXFvx7zNzl/NJwrAJk8EagZ+GvyparJQR/SF5tf
yN5msZLAWQoVqhIiMWD4NRtkLAjzM2Xeu9YvfomhfyVLJ5fHRjf1etQVsmmqabv7
NoHV94ug//tbmWAFeDXpWty/MYYMedOcOIfqsB7H1HxqxMZ3SsOXQwTAxt1pWI5G
NXp08WAYx6SyZ51zCXn3BKb39RWnOO91ILugDXb/OBFMawl0ItBmKvX7HwMSU+dz
1cNTChVeeWXWJX+VSDaezBuXfPjmLCWY3zIp9GxxRO9aEa1bpbGcksoRKNriuUOU
8zNw0t9MMNDbsrKYx7XFCInnW1oji8VKrwM/AhNKgTy+oUqwhnkrjkN83ORL9slH
P7SbnN0L3q7KHkmO3NV5XcpFHpNsjG+ppDWb1i04BVMnlAGQu2ZctRmkkoGBu0XM
KGQaCTD9zp+kszLDlxaUglie3hI4P2PdFRoLbxtnd/LIeo3zEbdgqacFvWgKzaNn
dV+miH7v0pGzkk7b+waarNnQUfGfZMrSYREq12cdzgVpj35/26RVr0vMn66KGo3u
dJI7MwHdYPP4kFmCxjriD/MRebD0cPbUVghZF1RGCh+WH/7yeOshG5oh+x4ZOx1H
ZPZwtBRJO7IT1+tfWcvT7d/3OPCznupRp+oaNplY6RIrFKTUAMv1eO5Ia0LwwI6D
kHA6eb/IbYMopUhqndR1CriG63ol1WBwfOdIQ/HpTmRk40OS3GPCiv7QQsYio0z5
ECJUhASUaPN/0WUnid0R7ZeE9/SdgZKvoN/ULuI7K/YmNiimfhnmmeJ/mWj1EaM2
+kMAK6VQM+sDo4S/SMzQ858n2rulVy9jrNdyVWF+q8UxKR0cFsvSVaCO6I91hIF2
1425mbNOeBpV/WvUyFnYzU69KtNuxlL+sZ5+pvnk5X50BW+TQlx48e6ptW06tPTY
Qvc8loTQIMb1o+au59EHxSHHUBIHEoU3upblBBRPt5kCAH0BVZH7WJ3NlXbUXKMd
QMYLoI8QUI/A49aFzWzW7rtZ9vVfi4FAMFmw5hVTrXdpVhkSx/OMbd4XttrdfaCA
5ZUFnSrFzT0br85jQ2/uHIprN45Aj4Ep0WFAX3PwczLemh/7leAF541YA/qZ3dqm
gl71o5TFoZbMTrNVq7sUzCuZVCBynbKeuFUI4c5B4duJNOAEskM57zbsJf7EOxuB
3KwBEfUYO1W7n0y/qFENSR90WLDzfy5R49HSgpQabvVlZUzrgftdykeGboZbwEfa
s0CMQ8UvgTIaifwEZ+LmWaWtwwao3/3/3OLc7g/r8HxJzqY5RvBJ1mNYyzPFsYMf
WAyOZ8a8ld412trBcHnY/sSAG/rn/mSvL9PUO6E0n3jl1yN61NIKed8RFJQ//ZFS
N4vqCB1YJYn5dPhVOyXEWGJ1I1vbE+6l69UiKlBQPuAd3zxQ/Jb33X/lziQRk7Ok
FYaKmPDJx1vojwkzRk6KWUrKXUs//M/yoLZyQE3GMoZ0T9tBYOhU0FS8YDRvNsUM
z4RuoaR/R6/OcBN4/bo0D3BWwCGVqCtnVIgiloppJn6X8ztwxFOVkODkHqrXFu31
8i/coTzC4MQcUsrHEIKHnU7onlF4H5FBGYyAPUzMW4ubelmO/9o7IHN7yEECTTL4
nX00Ytk+Q135lvfE9Y8lTKNsZiAf88cxD2zSy5njAvvqIO/qvUFpGKVrnKLCqM6L
N3HksfFwYp5vJD3w36kREBtufBQ19gc2bo0SlH3BPRz/e6Yd+7GmuCQIrU5HRjpy
/V729tbstOG0NwC8fXCm4j9vW8nxjpPNdcmS2f1AHQZ74SxRewPolI896PaBAhEx
Qv53uKcauguLCdbtN5EvCt0W2C3BYD4K6hlaxam1bZCLxobagyUMFMBLfk4MuZpC
HwbEQo2ahjInSpU3RTQGM8jv3VjcrmvGDHpzZwWcMDOwzDGDV/HadooaeIymrwVk
GhoIHxn84OZjZ/1vh+cN6keru1h9dRCaaO3gxBZBQ2AUvcYDyHWzLyX/nMn5oApS
pfaI411dbss88WztUMfoThVIcARkR8afZWfTWLPVZ2NlrlCBY21RucHDNzD9bB08
cmpW0V7iE1rse+9YBgHWVGXI1M/yCUMkC72jfo3L4lqvpONddaPQ2idGMx91T6MZ
fWzh23Hs4LzBtZLik+r0e1dtlifcVZ1ok4iYq4KjmPgucSwF6AEb3qV+Yeehornd
JldXVXq3EF7URwXMP4d2UIEhTBRfVi4HNN8fio55iwiQqVEZFneUFrt2G0FiQOF7
GZ4umOZJ10gDntsDc+zAoQj09qhTUWY1/ItCT6CqJwEqoQPRvlnMm3yZTUDwxomc
l8IG59JsFnySXvdyARq7kDH2o2GqpzEUACHiFEurPOYCKKVwIlTyEYntWFjVjGBk
vMR3ATXiOVJij41Je2p+N/qy9sytqvCvcRiKPUY3gdVbdzMLv0OEswuupzUO3ITW
SJrby0OL715rsRoP9KWtyiE57A+qm646nDTBgYMlQT3CudgmF84Z7zeneIUtp9eK
m7YnDnu57Ii8S3UUcf2OnrdN8YSAD4LegAgpPva8H9yMbhrrSWCCXuprNUgd4uOY
upaTt1dpNFuvUOZs0oHpx7mkQbjoXWQP96lgb15iMFOQefcmAkPur2rjuXZp3Br0
nTCMH/UVQuMbJYLhentw8GC0M5nuq3VPS58K+hE3Ja+kpNby71tZo67AQd5OHzBB
OmEgwA6+Xl3DOHV6Ft+4DY+UoVwVI3Ss16vrJoWpzvfEif5mQWzf0h4I2gvclFEi
qBXQ6ZVGXUqGsPgYHYXeqi3P55KoGWdZrOX8p9P9bIxi9MRbxSXUpLKITSkQ7NQG
Wa8o9lfoZSh8BNXdEM04n2oOLCPdZenxL6cIhHOTsgHo+dPPGKAYli2zFQ9aY/yo
aZ3F8CV95kp+D4GffcAix6+Eezje4XddC0LQG802DJmRgwCpaw2R9Jja3rIecBpD
CF29DFh87+hP6sWqd9v3N9bu6UnJhTpHghP2PqVITjemYNT2nPmOLVtsjPpteni6
kQxVL09k0gucDmqFw3b5YMN6hM/mF2LJWduC27ZU2S/NIm1l3SMRadGqRDeojTK5
iaAHpvNmbmkAYJI7BlUgqq0wRwRI9aiwaw13K8wuYZi516ilW/YU/Vg6qAsxLnGA
ZQ8vC/tQ0zz55KIyhYzc7bWgSWpL/7dV8m7NFwBU4KwACJ11YDzWKfnRp4eAbhLF
Nyq9sfa0ENJkFbf3uYEmYOxSk4zOqk9puGTPo0J5jSD/OgtoBhyBYp72dnYjgZeV
5eW/gAuxdTAScrHkOptezGQC6VvvS2ppaPOB3fVG3MgdnHNi+4//wvWsITVvPxz1
Ist9wDfjugTe0Qq6VMcgEytQlxRYYkpz+/7B1q1rD28DZsq7Ionor2eAmOTU5+cD
VelT84KegkAViFYr1hCV2U8isIIv9WwhWFAuhUBF6OOgvTzICcCuf2EKhr18CCx4
iS+vZaCAWm5rlbhRAtjOhhjyV8WSIZZPquXrW0ATrmIFMKPyV2Vdjj7OXaXUVrGG
OYCEtjSJ1SZTYPnE+qcpO1CoeO9XczREfukiXMsIbBdyjl1ejd8uswLhk6bvxbOU
W8wwbohlqrv33b/mzzgSAlU2Sk7K3PcFdj2T2jE/+qwPxGnrI+gi5tWKoeZqtAUF
03EYvwBrrxnKp+qeR4uvRqPh1M39j5KKiENs+0SYoc2VkkKxuXBX8NGyNDeAIM9L
zqqlRjPLzkrWXtoTE9/Ck5LSof0OlhDv/VDjs56UGX9ADDyqbO1prl3dmXAXYeqA
owCiyiPBIDSmh2gEZggHtpq+QVEQHP5Rj606v7YDzsps763XiRvC/fRt9ImELXyU
SwwLV65ya/6ju84HWaS3pEzLRGHPq1NYa/MHURthRye1nbXg704DyTwhZbCxcsJ6
JLYsnDFK6a7pR5Dr81v3HoqaySFo6Brx0A+1o4i9p3R2n+FGeXoFLLFbHM+TUz6c
X1G65Corn1Uyou0Ua3+ntcVHNDbVsfNJSi40SAF0m35VtnAdJwdW6nS2+pNPTRNj
9OiDBEPMxuWTW0f59L63fQv4Y5C6/glFR+F5Rss6BdTVReqPpaHWHkbMWRhUiYNR
Sn+tByFGm8FCvB8xI+QPiJ8mfrITDtLE4rpON8ilCrIf7tic5luvrnyCnyOkX1sU
RH0XLz+V4lmD5a6t97wMErvfDe1ou0REhRTaD4lOkc3ny4lAkZClnM2li40QcpgK
PpM3YEqcjScx0uv7I0Tz3AtR4gvEpWL+vV5DJUijcUcBVq/CWZlm/QalHCwoqfqL
p8cvT9uWybZLmE29hnvWjFiTjYm56iKG52Wgb9iMP0T5xPHbsR4YJQyW+uXrRfP8
7RM9c/mAjpATKidIOCLkNtvQqTx3EVSt+IPQ6Ydk1khp27UyTniSZq3ofue1Y8L+
URLeB5CRpFSAXZrbyfu5ZEJe9cbsTcRNjJxcFck2jrG7G0RDNlkFotirvANLb3aZ
zcmQuFBbTb2OICJdkxyeR2T/zedggtZfRWk216PKFgtf0CZj2QHvdx+FFohs1hml
/tYP22QOwjmeDwuIsyXNaws6ny8ET1lfy+/rQenULPbWaIH/rXaca4/CspN/TfsQ
GGSDO3Cbasuq4h59Uu7IEv6eFawJFtZR3ZW7pEMV7vwnVQLmRvCHfEwMH7x4VNJN
jHCYPHkWYjhhJp0XenSiB4CJ3OmjgkSAvYCd6r4YpECBmyFe25fwfd60FS4PIT3h
rfmMeZsLnUnyHBGsGnfY6quIsEEGYGuQb+LQQJHyQ5UjHRSzToRl4VWtWpuTmoAm
WHxpgAgzH/bzPly+mBiBR+H5KXPAEVlPkRRnKylYF9WxDUfYsCkbI54SLrRUg8Sz
tc7Vay0fdJiDA5ZwYaEOEG19xAF/SsO0nfeQXKGecB5ueh7eb2e0eq48NF5PiXP1
daf70L5wF52DG7UPrgO85/jWXS03uKOaqrlEMhCNj7h5NwTj0mvGSKXRrqkTU5z8
QCxsFMxPXmxr2FRx5fylnFsAQz2jFXds+yvuJ3LHywnc7oRZ+BisgslBjbzbvB8i
sK5okzlP86n6ylJj8JOrhIocYzvY/lgXkSBPQV9BmeJKr+9DP5xYY5aXj1FWrFJT
aRf5OtR6CI5hNnC0b8Wqoz93TwoOdwe4iZIQbhOullvwUzEDRZLbzLAViXydcx47
nKhrSpZIqDDsmOGO8QKK0+BN5MTp3EnQJv+X5xsgm/LiUfrBfhNNK88EltM36Dsx
ICP+IpHxkgI6rxFcrx1s2InPgSBqNFrobaRL2e7I9WJIOcB+YEFZ7isoTLOM5lpH
rAsu2m+II4cN5TRv4K2omxaGwlyTPHE2u+CEv+X1RCOpIerXQEV3Zyfr98sZOckc
wdYDGUBkjZtqqL3VYviflHJjtlxLZGQO6DrbXt/lb1Cxlp34oppb0faYBHM7c9WZ
ZUeQvfrsVTc+CA1DWGSgPoquKe5NohYYg4TjThQALIZ9wiFlc8SVM9+PM1jLK9By
5HS82robSXWzB4nkLux697/N7e7now1z3puoxdfvPMEn84942Lc/FQojAOYzHJNe
IRrYLLFCDSzhzfL3kG4dLGwRk4dRrorW0+iQ1EY2Yg1EFSzstmQ+7Lx4zXLwbT8O
scOwL+4LjWF72nB4IqKuyZDHjZImv/ZUR19ypfbldF0XGvA1xLOZyGVklBjdXR/U
ZfZdcrfaTJm/4/J/rLGIQ0Z6zzV9nQk+lAhah248A2P6fXcU+JMXbIoS6WxitMva
ALJDUIY1MGpMUb+BfFTgI+Sr1lCYXPv/4J5bagSE2utu1EiVwveo5SKvj9ewBvbQ
hddLMlzU9rR2EBFmhUBECaW1XYWJ2fZVwEWX+/fRUg2GmlnaihYEVN1acxaHxPcC
JAuN3etHzU/a4ZOwJq7fUpe3HMgZD9YmX3KPL5DQRRvVTzvKWF3+WLBMqPdMNSZ9
PkIU1U5i2N4C0NfpGr9F5jXPs3QPN1uwkzojA7GwM8nRUc9zR2+JII7dR6LUmWBr
LRfG9e2zrQbxhu1SK4rxPKBYLZqOIMFXQTwWl1pDCFN/6tRwitsmJvZ+An3WO5MR
4sYwLkUly7zBdBkxQqe1slc/rEaLMYkkC2CcvVqf78hTbgLx4LKqROwlmuRveuXl
G3F7bekmt9QLxOb0Y/qeLOFTfVeFpts1oxwCZgCqfslZs0PzOLB18cWnFP0/1bjT
x9ZqXO+t++cYKyMP+xVBOwbyzu36+SiEUjwSx7hYkd7jSd3lNsSjozGX5YZOKIeD
/gSl2Og/3zLOPCw8s08ea0W3ZhKS8WcpyY19OBl4gHquEkdqXBMahhGfQPI+8aYX
qkam3PDVDCXpQEtGuVfccmVqWu/6x/RB613fOMF64btdvEYg6BZjVYomxelhxOML
JDmXMPLh2z9H0gtm7O8VuIu5eAcTVvq5gbFblTjPkI0Rz7jHY0LaMBaUcy2OXp6f
TLtqCzUB0rbW94s9THN7u+0MBpHwR8tO9xegfsdpu4GURlf0M+KaIMCfrJ+Ya5ws
vLjoZuGpH7rmbZhaZJbS1NP2YaHxG0aO1cevBUrHHxS1R9Huy3nIXbl5KkjfDUiU
xyUz9f2EtL0gmhj8fy5P2Jg6J3IqXbctZZgh0qtUIG00kwe/t5TnM89Mo9Cby5Cx
jh4m9+NkjRw5MOMIEdguf1uosuBod/Y6svDZ2qjUzuT9jk92r5gbA9ubLe2Sv/qH
9Il/VwSXjNzDPkrIk1TKDEDr6IHsdvT3eo2LOx/mGf9ZsjsD25erf8bBUc8kve3t
CqdUoeetaF+EJ1wlQprCm8h6H8oF6CFDz9t7ltHj+5HWlbx/Zw8kkbUHydGomlT/
VNa7EXbGN8CDNgDev+qtYR6UHkA/34NBLH7g0gpYZfVHq4x44hNhMJEf8BMgZdDk
ToKNDLCaAkKzLKX9rhxv1DIu1ZtKV+69fMM/m/03k3GxWIXiqvtMHqitBcO8By4f
z8i7qKCNPHWIm30MBYEQrZeeyyBtDcvBXf6pfZ1Db3O18zBSrtu8egICEoCKeO7C
IfucGS+7HT/Rp+oqqnjdgxPSVrSWVuYWx5Fsczm08deg2P8nuYHIceRBZM7KIDLn
BZbHROMmGaQcRooOfrcrPhPojPO5CHYw8K9tgVdFNcP8Em80mPGvLhyLJe+CN4Fr
Tbx21p4BqVgbYsxv4600KFExD9MAySbfMAB8L2q7+gYgGelCmwzIPzbBYrrjvAHN
LRuUsBH839csazmS9FQgDDAUP24bblbl8VtL5ZN3Fb8PA2XpZp/eo4XwY6hd3r6b
Yb+IZkg+80Awkl9Fzp/lNWLhXL4nCKJSDOCHPsKoV2Hd4a7Bu8uaCR7g+Hvq//B6
bAZKQIeOHQmkKFXhlVOs7/KgfqQvUneWnI3KVFytZptA4FLvBVuywyYejkiMQhBp
IHU8J6gyfWoKDp/jrdAXmgvu7Gf4B7Qx1L4p+roWcRNn8nxV2tYMMQaxGjIJJ416
GVnJq6TQyAslWYJRthiM8sQ7E2J8UZyNeY+IXgaHTSskWzIUjcYgZv3Oy2pVLt0O
5UolCmTThywZzNJjJNFyaCCiGuMPVe6aT/ThLVnieJzOn8sPhRjAvO/TYR4Af5NX
I44nRXZrkbOfOoJg4yuNt/kZrBATavmy1fZUQt77sj9NqcTaDv9eQl6fRcnfxH9F
ke9dMolB/VieOjOEdTE4+/GjGZvYLFYdA4fmm4zbUs4obvqy+f9oebtpgxwDNHAP
nuJK6xZpjoRTuFLdwZA5CevYgvyIN7ywUHQeOn8pI689zzEQHZkUMfgeg7KsTGbG
Gi/E8UET09r5C9qwPFbI5JCvvoSMgJcVPnHJJzkTby6FxLrnZGwxfgY+3NWfvMUJ
UZ4C7vDxlDRgPYDxhTyUCF3mIAvs2WCcFxU7zrD7VvLnyX7kYfIgHQ1pq4eJEKVQ
XwMrEa9va1r4XuXv5+LCWiP8MCfg4fRBnWFONbmAYTGUeZfaZSBMnG+chRLzIs9c
NjvXL4oByvVqBIJnWg7Zf/FgEo3n33NP2FUsduPV4IHFP/cVjqsVB2GMrZFBJ32+
x2z47KB1pbPZF+J8HQf0dntpC74UtT6AHn1L5uKp/aAbQnj+POGAsCkhK0RUOesB
IgTcmCG98+9Lt2teDALlTNW18IswB/fKeyBPjMxDUbur/yAW3aALjQQYhHp+3Jv5
EM5Bnz7jwFtDGfVlWlltRnJwr0vn87kfO05tM9CoDPkFvWO00T+A5+/u8/g6rVyQ
uzRYgnkgt6RFs8EeMrmUI+a1H1ObGRbmDFDXub+9HqJf+Rb6NEMM9kOzEfNEi9O+
DAvlYCu1w734KBqSwQ5oZK7vnhdDytZLWfWv54yLT2Z/a8sktpHwei9td081yvQ5
Qli9CbJI2CqoPEUh5MIQNsiR2w8M6TThuIYx4TjldXToyz9LMydThbfWFF4jmKC6
GSBfS46tbbfrdFFZOTBP5gXyMo6KI8NxJS6KKk9W6CKiUdYdgLB7HG6tvyg8xeP6
4PHi+4jFMUss3e4hRCXxDPScWcJFXJ8CfvFo/2gusjcvkj4MpXbmmsyME3dQc0T8
XrtULhRy+Ay6JswFKL8PPNIZ03t8t+n4FSqDLoRkatajMsyj16a4bLRj9++XP/8E
gvoAyr8iDkut7g3vG3008hiPTvKJLGW3yecKqdTjcVLz0ECSFYMPNN2nExaVaKOi
1hbRQ7XcCObdnm/kn5xBsNCiRpEw2xepzIOLgs3ORZ1JCNjxpGUy6qhTAe7miVnb
YUmvqnUO4vi0sNGUYdd6Iv0NLS6WIDD/UdqU62ObbL4sUWvs/uMkegGgdRGVAtBO
oojOYX6D80WzsuIAQke9tO/FLlDUDAykoB5T/D+ZcJAetjK8+MZQ2lwlXflHTa2T
uOvPOs9TiXG/M1fkgUs7S7WUExT9a44vOIk3kVbyhVOT3mz0uX0HimNca8MmDMxX
CZPHSfzo7cZuEWo1c4M6WlofN/Fg3kKl06rx8f93Sx8C8x1TzEnD+Ju5z6/eETug
syf/qJysULeJT4rDZl6PMNSocvFGHD4pjpASsspLXqK/zvZ+XGVGIGO4FKSBR8f+
rYESRrQ8FRbMeEsKtsC80pj0N8eE8h0mE1QyJh5p/KuevlW9Gp7du4jotjoO2YKA
9fXEykvkEPiuefQPQOkwN+wKRVIJghw/tvRaum2tpVonE/dRBJXTSE8dDwHR94fE
FgxMxC4QrazFPPKBdyw0bo38jckBPg/SFCaH6jI9UKqurShq9USwaRIBwr7dyBRl
tgAYpKxcGVasQG58Qw8Dt9Q4FjW9Sp3Gv1vkioyaoG0rdNECogW9dEccG2VgsxaA
y6Jk50KfDLo+CpLw8x9BzXzxLW1ZiHFjitd3U7q020AA1V/vGljSbSF7a6UTxeZJ
0gzO+ZmCtc35YPT06D0r2lUvhm4LZ892XdDx0E85H5y6wC/58DSLBJqorXDK0qti
28+0qOBD8VmDE3VNrXwZV8UhL3O8xvalA858ujvNkqC/YMYWMjwfaiUhMkP+Rl7o
PMZnl4ox29ceB/HefJMltUSnjdcoahVvWk/MTBb5vU9woXAr5UHGZnGVVl/4lOdk
6k578ltD9jC/ZeZFpDn+zWJwZEua45RqveAubPE2d5FM1NI1NLRozglrpMNEcIh5
fLnSiQtDI9wR58kKkUw973DSLHMx0g3wfTflkXHZqhUzrEpDMqizBWSM3m0LIYnP
+2h9epU6gW10KHSp0vJJ6o0EcW6ckdKMDutH/61iNuEduBM4VkE8rXXvyM6nbcEF
iQkK5GOqYuEeuc3elnU32gitovjj/UxcKMCGJWM9HMfMVss5A/7oXAr+DoxV5Kwv
TXlCgndDsyocxZjfXb251/PtUvzZF2X6yN7v4nmj8osQjPbEMJA0voS1BbgwOnI6
JePyWdaIqR0fiOl/ffsWaHaYa0j2PCBt/dVdwJZcZt3LJP5thwRAiBSGtIkyWbZB
J/LIYur1I4somY3+UiM3fTXSHdUIgjtbygh45ouI3QY1AC8wnPnxgd2D5Q6UcR8Z
PLpdNwELmdBjVX0GkR6po8KyYAY4/dteqFIt9pJyEjxmLfXJRgjM3TM8vUKf3ZQ0
VcDAeUIQyx825d/PyoAsy1x+Kr8JRlnZ0debZQEZ0VYOj+eQz7LjsO+pNz2cjyWf
74EzdaeGHarxSCGMWhNzi626Om2+a1Q039RNMWw+5HvMIKnqq72Tv9yyPu7iz/MJ
gxnSxqOIUZOGGSRBmI+mWHW+dp5QQEU85CsfLwEyr1sY2ZaGOOiEL1+16+7KBqe6
mvs7od63foFYXYXkyitJ2ShWBzNNHTwMtLgAzxCHoxRx52aMXjuTwbYb+nYH1EGa
JzO5j8XjBnisZPv3AfmMaO6DYSnK4fgVnrk0/NGTQaAItk8AK5ZEm2Aki97Kf50e
i933e0QtE5k9bKSgVf4Z7cEnKVkBnVKu56pLufTwbEbFQLkP1mc379UBYQ7lmYUP
0i2RPglgMalQ0G5dQLBd0q3SskXY8hC74aaMAcUFpGrLZUpvL5qrDq94YAPpGrs1
xO1NSNQDA2ZDlJduLjvM3v/4oEaiV3E+b7H//5DkF7u1ny0qmIVmTSVVNTc8qu90
2RA31H3BEzJAe+/W497rQK+EJVz6gnKkZTPwpFOLY3oqubtceAAaDwAzmG7224iO
s9LmAtkriUBQrbKKaTvX48G9zxi377Ul0D6PjFRWi2ADiij7Ba2IWUghi/LNI6UD
t8lNDyJr8JNwNC2kFSCDA5esqjcKtyUdm/QcOR+quCQ65VW7zWuAAA1QYPwbXTMb
YfKAaorZ6pR1dtr/HxwO9JH4givd5MhggTGElsw1Ak/jpmnci2qtofYcHnduBg/b
cqBwOYLnNeyZDZe6vpa/YsRggGX4yvJ/HY1t5xr08cYtEOEYoXfm2dv7WPW/75hk
/ARlhILUeqdy8f7SaomYc55Z03neheK/eNzckgMeFDgTF0GnAIqtib0pQvUGarRt
3vvkeLYvdDBJ2/1zUF7STYri2YCTMS2HXPl3Et8nn65OektvG+v/L/Yrbl1ZRKuM
oBljOcBzJxnjZuT3vo8Vq9/D1GAs1ToT3WoEv13H0FOfMEVweEAE9UHLWiEuOkPi
Q/2TEV56x+DMxcXr7VbrtXX5pqS4UBtxwMt425qcpPTkoTMTvojcPearpF8lOJ7Q
prQ3pB9SPOB9OXfvuIPF4uZyvjj2uMSRxiQi/NSs14/InIaDOt5CJHpyDyfYFAWW
b9GeLgtF0EnQk837AwUctxST/7FGPlifGGEMjoVc0PrkiYefKmglYKMwun91Vzcm
W1G7gfBJIy+dSl+8/OnAtIAX2VpxkeUk6vdfO4Xi8WDp+sAOi+75TGVvi9lBDLmf
et9/J39ZaXK2P2pCYZjaApUNVvkrxjs2V60hE+LgHSKwmio0tJ446kom9cPKZA4p
PVQUutTsQQ73Nk8cHC+BMlkLS6OFvY2lx1M4yx4knT8xptR1V7QZaWP3Co0qZlAz
HCqGcZqkTxkasALPZ3tzez1L3cnhXSEcywkgWs3gJ+4AXntL8FJnG7EKyEwfoGpg
KaPyGYqIgIuwM7DQ0dBxVnrylxv2Ypip9TCMxvpGEAEOgmWXyDXEv7iD1dwEETyK
qnHpQxeui1Zuf3KINXRVV0JFU4OiPyTRLL0bxjVtOersFsVz4bc1VTLSmcq1BvX+
z7YzoRNvL9HDPbofM1r+9+S5uk2SBVBr0fd9lagpIXEVdo9vYPKyqEt05DxI4326
PeSw6DBrKjN245OFXvEvQ/2D97PVKNa3pbwZGOsP3e96m+V7N7SfvpYy8DjwxeO0
wkyGYPgkOCvAe+E2DgW1SrxgsNfJ0Ticx+3wOISWK93eQnF6FOBd5+GgivSYk23n
HZz0SjIoqx8P9GBBaygATWS0QTVLPyHVkHLYMMIKRn66y6X9EyDqODrvBYKvc1EP
hbkDdY3ZxYq4mZHvhHPVR+JLqgEl3cV1zclwaU91fuaq2hlo1PhYjCZAbNUILqqv
Qrkbf3AiCNU0fyeu5XraNPXiFnsJ3SKcnGjf20WjcVSIU3lBtII+WIMryBwBTETK
cxdsYMNolJAy+TXFedpt2f9InL64DbH28GVlAlV39TFaHPPNEvOX1z7jbD7C8lcM
AXA0adfO2u/O/6GIOweShwVKXqhlroT47AR0qlIDEovJGzck0sGs8+vffa4qnd/f
xX3Lb0E4flTgDj2+zDUkKSJo60Dq/DIHGEgB9uSWsjvBBBCO7UQ/nDABOilMfaeK
IYjnv1lVW4sBUoOcUqfdAQxUnemDdfUm8r15uQE9qtCbQX9b0HNrksAJ/n/qV7LF
qY1Qgw76aV7efjDMNFHrXE3yD5ZquEUnXH00ZN3nPwc4Z+mJuir3W6lMBS/LiSs1
4mQhoF/p3PCV6bslwPO7T0pGDAbvuh26wxwPbTnrjWz/V+DN+nkeQMjvDnrOlqEI
z9h1duyJkwD5rwT4Ee1CSE8R3hbu1wCD/Rkvmwfv62u+X471N0ZAXW4VRrgfwLfF
iQF2mM4W0M33Ocom6qVf5jQHb8kgStDqnYqnT63Bt2f8JAUO9vvUmFaiM2hb7j+F
2yIv3O57xghsHxDu2qsw7szJbTJsIwuRXfRUsh4UBDuBPeJF1Cb2tcrRh1VUVWfZ
3jQD8rNS9ak8Vl/MhMQdi9ofNKt5hpkfgq+TT4+eHcOpUM3BN7U7SVHlS5Ya+HGN
d/dpYalBYly9KoXA8xgDcnAh0VSgvOWvpuxwkaOEmhFJXPGANpT8FMb6fV6NacSy
myFzB9Fc0dhIkwXqFsjfQ0COTTb9xB681ngbVSurquV8TU04Ho+L4ZXIc337/d4E
qXu9yrmhg1gbhONUpYSDWN8AuZOqvKHOCBSDeemNu8LCdl33N4Drf1P19YnK50bw
maNshqgcHTpdkAoqU4y47ptWe9paM+ccQN9xNcUl0x4NbfvkRPP7X8TM1W/Dn77n
ClFHQL5ezufpZ9iw8VaWw2I1AU4ASO7xouHSK7PfcW3svvZu3jOvPns3zuyuLYLA
T9wRF0S0iKc4CYrt/BOLVtw1BuTZDRPvSSnmbP0wdp3H/be5g2/+vN2k/b7p2R+b
9zTFLu1UO2ddAobcyXATFflDEvf+O+u7zYDTfxyo11rBHdEQHQ9LkoJQiI7D2rfH
wiRvNlHs8qiBXNAO5aM6y79lRiKLAXU1xPes9cJXbUUZ1fRXecisYeiIohdlF9ke
IktNH/ygXh7CmjQpLrfjPnQspuBLNBUDK5kwfxgSWkD/4m06eN1fkdxehdhlt9Vl
7XcFmqwRnsFw+roWUcHeNvWnjH9gCP3HK7No4ugN0xdcnVcnJOyBndXs7bnfyR8a
RABuw1qtnAWYvcyXH2ViBJlTY+K2w2IJ8aDO5lzbZNLYwMAOKSA+rZWfuLgH7eVB
ynQTk3PHEWvFYi2mmpHiY4TWTtmQSwIIYOtskFZfHEPAvaGyRruVN3s/q0YtwBPu
oN1FdTgggX1CkvWvWIZ2Wj3TQ49Nqf5zBBeY3KgdanZz1anWYyl+Ts6/DH8SmIYq
K0bI9VF5/Bl/2haQSyj3eh1foYTGx5OAlhbtdT+83hxkkhty/QGf7srt5Tj7jSB/
Kr4iK4uK+SLJyCcPK2Rg8e9oCDsfL2qmRM50ZJ4+xeMfJybehtDuGXOrT38BzXnn
dZo2v1YwIbfgSq1oeZcLPiMFCuKPUFHe35N+fcViQw7e05D2hNWtWKBT90ORH8cQ
KuEUpSOKAqLRNwLRbdhjKHthXxjzMoatvJCVapJJrLIUBrWHMnRx/Yj0rcWqjMXJ
1acNu0IGXwP9i53EhysqPpGulI1xPXksnXKwTdIPeMaRAnLhJEr3cIx67dPMHqeD
XZzUa0zbr0bleQrx1ypf2bNybH4aOP0xJ79S5cV0o9h61DgvXadHdECrlxIvGbCE
4x6DRaIaWOaX/8eHT7wh2EHaE0T0Z0wnfRTF0V/lXPvO5MrdOZS8+g8Pqn8/4QRg
oXvqQbmgVb3USbByHrCcauyx7OKjklBvqL07t+ko3ns2pP+ce8Nu5BoQ+DryjiUE
iOw/DGYcJLx0BA5rZPxiUhrExW4xNGTn+sq4TbATj3oal04eFaI7LqZg/EhS2b07
MVdHw1v0K4NW3S2CQ+yAN20pEbBebGlepbficliIgkVn50KMVVzqyHRoWANzKlX8
CcUqVmbIFX1dVYYYSPCPsoRErYcIhwdJzF2qu0T2ZJO2uBdyg05TfDNJo7T0iqTi
Kg6I/6Cz2MG+oOGmF9s4sRyQ4S92XVVxLWfugh50BeBLsk28wYVsJ98uh61Ox1I7
oEbxiRL84OXNfMk4bSAVG8DVmme42SgEhHZC6AgLxC2kKECbUbKxr9sFDzIVxNn4
saVjRyMW/X+3qYgKdH5KMbhDmYgG0CjokI7CDqamvpmF5LBwVZRIrtrnwW1ugqW3
2fA+Y3u/w2Ho+NaT0DsveE5E76RyfD6fAlLTkx26DXs+0T4g6D/L56w950THYkhI
fDpFBVfbE7aw5qOIduPLupAe2T8RRX1it+YMK7PX7Nfw4xKqj79QgbAWPrx006Xc
j7tLUCe7AIKe80BOYhCrWXsv8LYf6AxNhhLChD4DVml/BwwNJvK9wphB4akYHus3
yZ1CXtWEJxWCaWv6kCTsOKBWLJK2yzFM5SN2+9F9UMqXY0vUpXfrh5QmFcYIz9fU
Co3wqkJvu5XyphobwgGuOXA9fEYbU3/gbNSGaxlixB6fwuAUEuaooJBSy5kRJMNQ
RijAdw6P3RK9QvAWp9PnjMZafxvMzWoeEY8e9OVj/FCaPuMT6I1FSQpi7KGcRCC0
KaROT6NgRfEFVhCu1pnvHUazr5ttfqwenIC4MMMSWQR6AK1cslRElbZBiV6qDdrQ
uarlTZaGpxiPvnwHKoyLTaaQ2d9NUg8xYcYCh2FdzVcCD5DTjN43ZjCibV1Ma3ER
hvitGcRW2nU318cVGSzlsBJsUN3rh59Qgbes7eY50Vf+8svJ5veriNp7LpSfEUvI
IVTdqHQwlazXOprCQV1EX5U/8QBdEygSToSviUgb4V2OU7PBEPCOapRjfddSbxNl
ApyOi6Z4WHGgoucVsCdZn6S/1FCx4wxzkTrzzwMwR+9DtSB8m6AgoeSNiQKLSr+n
bEzVp+DbYgyp/EwFakL4a7u7d72ghG698crfUKXURv+8KekGw4muHssE8ZVqIfbq
6TbOpUD0A5R+sT2WJDbfLQCKUWZzVDGyUlrYpGtcLaKxlp6+BHvwA0Bed2+bwJ6F
wRNKohMSTYSoNo73shDMYZiuJUaPdax7Suo924+3WSKniitgKPBab1/RDqc0OXAB
hmYOVLfQAymfhCw7CuiwkJlnLVXQ6vjTk//DAI4yPiqu0odkCGzKuFix/HII6hLZ
52hiFrGW8aY1yxxGavvJ+LdsBUvXwDnBqALs+Duykn8m8p94OgnC5OHiDBWLDKBI
e59p0fd8ot38HYiWnEx+1L3QCuSq1KRfR6ucPvcYs7QoZ7fNQg+4yI4QB9bRrinM
M2Tq07WD+Va9yYl86FzZLNhqKt//r7wdm9bK+a/xDBYfkWCQB72o8zMXVgYQ6rSG
LFF3OpGbKlwit5dHXV/4i4YtvDEkz5bZNGXYF1GheMfh/8S3F4d4Og/VEWjWqKa8
033a4InkjbnZuMVg8fnnsS6d86XhSpLBD6j94JIqPAJQ2oKYvOJJS1rlgQe4G2q+
r88OXhbzqpqRc5iHvqw4iqoxjelByVs6dUv82lT/SckwDiEns3pAa0l3S0U6B7/g
zJrJjAsbFCaSIeo8IWZs7WmP8aoVagsKCIRZjnnt6IXDkl3Q7kN/772aaD8FSkx6
3kmThC7CqEZCFlIcEcqjuLpBRYGbFMR1kXg8HQ5SPnC4qtA2tPvEEs8RoQdqpRaz
Qz59Uw/3sUb73yRILj+hwFRIRY/2F/SIOKS2RUg7EKFq2H4thy+d6DWOV9R9xOv5
fhbIgpfWHGkJgeYPbF/NWH9ir7Wgvqhvaqj80H+OMuCzrjsCjO/Q/PyVts4E4Twd
iNL/Se3DL2skvRESMtVVEk6lRMXFnyhb/2vOjSRRcpWT4iHHljXUyLxWchhSwRMb
nBpU0No7kXJct79x/Tcn1j81DEgVz2rVCh3Ql7HlcvHBM6xZAu1/Xa87SDNjbh+E
jK09ptFdxdeSkRLslZ8+tnaxd+9NtgIN9RQvFLiWLc4T4EJYFky+HwZTmnAJ+CC5
nxHf/9CHojWwiAAyCX8nI5q0XzbNX39VJB5BBDMtB1fDKMbHkMCtlurZBFz7cjOy
3o3NZw2+Nd0RnMMHRfwlZtau6ndczt8f7UWOjehEc5ApLI1+YwsD3oZZiRbcsDNC
C3OAXuK23dEITxgZY+aAfUSs4ki7mE7VKyzjaxZ4H+v/nX/9XdQJfkjmNWRS19WW
NxLXI/gw5I0nORSi7qS6yJHcQYC4mdrX0N9DEo8CGjo8fxDZ/tvsNur9YsPlh5+N
SWomkUju6igHvbayRX8Zt80XPjTfGvubT+b3PSjxDuGWjSs3jdyHLgdgbpxzHsB/
BTTqpEF75buakv4wJQJbZ2SBwliVSxkW1vfB3nj22HQwsI8IDhnWnqWPNMltFbG1
5vR2BJTBrBmoYlPMWizAQ56Dak1ACAyn9Avrogl3Xeguw8m9vkd4GKMS2dSoUqni
3pPTXQMG3jm64D5Gk2G9m1fvbYOBB0QzT8v0p82X3YLINrYDnqZgOAKb8ryCCe0i
ltqEhTMUrSMXhcWTx0bu1ziZ+fB1xwvwj368zZHKVsE6LOB3HZ6PAaDlcm/jqg4u
wknfOcd4yzwGqBwsu6kfndo9/EdUSlndU+irlIFsG560YWXOvK9Oi/nB47B7sfxN
/ftb8+vn0hPuBvKQ4/ipt0jidcsRDz/8ot23Iw7XB6xlHVREemDiZjhklu9WL9Y5
38Dhe6EwZRLib2AdHVPdZ1SkZRF3vHv/L+SWcMqmvPEeCJRMx9IW3a3vX0I6QvTe
DrO5y7Prf1/pz2blsAvdqYAjDGOMhyPGFCq7u9hgeqDloz0hAqlCa3GDaDVrh277
iUv2dKJH0Slx80rR1INKg+95ZSvZUxBRszf/2vWPx9MNbESxI/mJln/o4Q9Myn20
Wpk54lGnGBs43QHWc8VIhuVq3FcaLJ2OdyP1qhf2S8NyfGiqYdcrBA4dqA0p6EM7
P9Oxjt2oH1xHtUYkuKbZ2XAHZYFMWo/yrZIZ+I5Hw93SxIefDUzIxAyBMjgk6PHq
P4tvUhbmGvFz3shdqplqy3HQUKssxQ/Am2vg+HLD+7Ngy0KYDCEU43ROCvqPYMbl
e4hDI+qguF57zAZRYgEizl00y2/HJ+s+4FcnxrPzF1HdXJ6nM2bMXjShugzagssI
Gvkh2r9Urwf3pXMLkjiIOr8RnT2RDk3yp6+9ANDnKYj1QtcHkrAuxTtm5tF2EHtk
iu/y9/vztWpbzoOnJ2sDgntpCR9ICGXn5/MK7zgZEXyGxihrKzJsXXGhbUVXrcmW
tiHZRYGi1+En8T+nVQS3qFwaaUAxmjekRtE5NHOsqNFJZisFbUaw4/+hSSKjIRwz
GJP9gP/GB03AWyp0geTqCqIn7f4U8tVSm7Ct5p7xjOO2gfOe2nlDpPiLF2iDJw7E
ON9IQgAa93WHQrXHAuqsZDuXdKE3QO1FvUGyM8uPlg0OWCAlJRkXoTzlfB54aUDi
IQ6NOTdho2Q9IGXEajAlOrVc2xyNDZC3EBagtvUanYIgwoxVS4jqrqZX0fCfsDV6
MRYvwns10SfhZvjo5rkNDSknTtVNiHAthmKp/otDcTq1+f2SGOO1P0gvof7FR9jN
DAcyJ5VqltkH/uWDXQb2PYT/B0ErGL6dW6+f9ignTCCnl/ilUrQU3tiX1iYdORz5
EvIKDP+gXDA+vrdnJMopsxg0Yv5r4Y87sGAOtdDpph0QgYdNDxEUL6e86ycfnEE4
Q0C2MXhgUBnFB6cCRLWo9ZLEAHecJEjHXAEbRGGo55WBf0CI/QMFG+Chm3ilLPU9
3EJn4anOOpQwKaeYBjePhNYYpQPQnxJnesDus9Gn3sifqk06DTGRj8NHJww4BZy1
Nsxk3zaqUepRAm/65EgMHDXpM3IHIILMn8F5tgf6ywj4vnUWhC7HItYW9i4iOuCA
7eOFTVFd9jb8Ll5U6J/W9dagC75nArwgyw/THlCBHHPWXbEA2oE7Lr3HMI65ltXk
8TAU/H1l5J4qtnV86WNPcWHvvIrrGn7rkF2Izh8vzUibor1+b5wwWe/o7FJZUuOG
pb4YHUU6WG3j5emdGIIxwo93xRn5hIbsVPUqwOSFRfs/q2j0XQutogHh2Z9YJ8rZ
FuwowzbhlAz0W4eWrOQD3SyPBtwjdRuB6FXDrTZTLzwBMC7AcKLrAd+OQeLUF+xg
FJcRUiP7UFr/GRI064de/fslIdT9CZJ1OFtbfyZ3veYr4PUf5SRb5wlfXHYbi/Xb
sWEVC6FwNIcUQvlz/C8o8LOJCWCswVV0g0jcwpcmWiWck43SQGXdcX1Q5MPcxjQ1
0sYnPcrUH5lfPiv24fsN82fGg7/Bjw5HDQIkxcovyAPdOFrn8a+CJgnqs7XV8PT5
zSXJBH6RqDlZNoCmI+CKsCmye27CVNteNSKmwhWBadY+vUj3ARmnUZxRpzxt5o4J
qM4cy630vsjMrKS1pBzjJgOPGh1xuXLIvB/0dzLI24WtOVIEnCNVq0wdRAB/FMpK
gRKGba+f9LTrk8eczDb2wnG9HBBjezXTc57xxPX+ld5hzDK8rf4+mhAxkv4TG4t4
Jv6osYZ2Q6nLHJQ3yMU9w7BcCe/mdOg9nhONnDjpAyBSf3OjkwXXXHTz5K4cJKFX
GIg0vKxHrBHrSklnP/folZyU56l2/bUEOtlhOCAJOtNWNi5/ZlA5AwbozjN7UM56
E/U+0HPvPjQChClcx+oA9u9slPQXaPtaj6CyVQnFF+FWHRohYsbRwp0hunB6dHav
GPgq3Btpo8fxg9uDAyKmQPXsRmiNMGNPh78D5xTbq/hOoBZx372W6p7xSdWkLSLW
yYpI4imWF3xcr1RCnU6ANpjGUV/mdJ0IOxrFBYo6csn7M5nPrcwfsJm19rAN6eFY
Q+/PYOYy4ztnbgbVZuoWeXZY4jQkfYSG5cZBhuVaSMucycQGZdrKfBA1a1Wb2HSG
rPUsoZVxVvqBh5tJURZ4JBqusS5uppj0iydqD2NMQ9H3jRwmu8TupAzXDR5ZmOK0
zJ8e1UU1HXX7ngnihs/3C/pR2kE82vhFl37kQFoMkNsL2g/nAz7X11dWmVrvO6qc
9a6DzhMJucWaBcWd+Cm39ychF8xi2Rx3GFPrhHrVjUOpz2Iq+9K2WKoKO4z/3v/o
gHnaO+UNS8zk5J92Y+wTWEzQ/c0bJhuMLgLtgKjfCZsBmvxDmb2W3qTwjSwrMYcD
1RX48vI1GR0189ETtmuDAIyE2CZVIjamNrup6767cJw+NvyxxDwai7rVc6TlPJWV
A5Nb/jptjw14lJOf406mxn4P1puTHAr6VQI4x0aWezRLkNriV2R/dukrNvyB/4lg
9v4SEmUT0HOkgjpQF+rZqQxTTZ4S02VXgxzSG4DlcNkumBAKCQ0Hm3RjhcWccgCD
kEXsbokTn22UmncCDRFNmMtMP/xpzUWfZqxrDllaAopE2qCdjB8pTYcfBGsZPOW2
0EE/9FxZrnNG/5qpChXDW36ULcfviNpAHF+CuIQFNrgiXrhItPb6PhsJh+bv8pp2
+ZGoz98d1iV7Qim0gEr2TzbU5aH09C5shJpy0IwiB9mkJWIDQ/rGZC+kbUkX0PPt
UuS/FfwR89WEDTdGP/PO0TBYYGLDGJ/aoa3cq5a6/2fdI/Su893OpKmu/xOdfIXE
lWLmHcIrFHa0vWw5poQ2JsnHm66xUm0OWqaZeOz/XLcRF+vjmiCZ9y04EVsDoL01
FpJyg1URpL4Jz5S2nCK42dNULzrJkUUHKs00Ga57Rf0xlFE13fko2MxODpOzB1W1
Mpa3ZlCnJZ0QXXQ3jPcT+RUvst6o3yXxU9Hg5zBbcBr1dOE7YSn3ls4oCwHTr6Yh
8AiSqE0wSqLDoOCfSl29oxiTrriKrcl3FbyD0ChvHbO/LtFt5BfUotwgFm2ABAH1
cWJl9dMKCA4rqXdNyRdCFFEV6fB4iQecJ1kWnW2HA/vwwz0xMdwmFXWN2yBq//40
CGFQlw3pjNaizVzIVewRBp8mU1DZzcXctUTeGP9CevnwbHoYBvLs7yI+q1kJR/v6
CW3LUakI9aNmkE/0MqIfWPyrK2FGKfwXvm+hkko0s/ukdD9KLcL7codE0zhNY7gJ
EfP6yEabUE7RbAxEc2JjdLHmhSRTI6UmZPn8xQYUxu0lt/Kp/C9Gq2gU2NYxRAC4
9sTg7zj+9PzfDwydNbjvm+fap+QzOq8YAYQUZLOVyhH2/zof2RWEY+Q8bzZTQygG
LP4UPu8Q0ULBRDqdr76xjHTlMRCA7Xr02ghi6n9NKXsIo99oVBO5WJbU0fIk0kBo
0oYjeaDziNG8NWIlZyVjcf2lAvPiFDPJdLwcv3jicGTVw3p8oxcOcapYsKVnTKgY
rwmGRhNEp7vB1MQVvLa8Oc62feIsL1d7fv1MPQ0+yHVIeejGsm6g/dN0/LevYH4d
Kw4NYoZQ9wqs+NTY8FN7mtAHrZg7NfwmuiMhnruE6lXD6paUdbhsIc6GhKFwx7gD
JvoY3FX9jKe1j9jboxP7GWiT3YNscHlITHCEERNBU50Vb6gSOk/X/0vqonjdqNxJ
qpMY/ONVQKZg5QmvHnxnJZw0kdEsJw8ONei+C+ph1ElMGHMURHQaUBr0PJhVA7IT
Xeq941BWPT4xfaQ6BTJvA6wQputkyzH41JmuO6mxycf0c+3TffDb3DElSHcYOCHX
ocZavykLD1ShkLcQSh4Bd55iZxjKspqeASRfk99dP0CFzl1LZ3vEd0DVgJSaTdHd
YmxQQG40z6B5p7qxAZBkuTRk/7IYr6qKw1fAFlgP12hhxc0ruWnljd9gjhgudyAf
jPv5F++uvk2hZnS/fjmubksAaGSkbQv/JrrwRtNJ5p9E7aQawnWAf++JUOQl4+HZ
TKUG2iFUtdu3Jt3KFbNoWQRxp8V0EutWhuHrWMWO/8ssY2ddzXwlwGPqbCyB8Fmw
cDCxwulUi7RCxyboz6bQw/xWfzmIr3KiLd//4+riLIJ6YjIRQ+bEYmZcvYwtZHzR
n1UBPBL6GGAsJnZK4bgO3XHXR2xEjLoEUPnFVweDNQds9pcfoyazw2UZ+bIKzKqR
WrZ99igv9rRX4Jgpea5sF2E6o1nGFc+M5WOUHsIafbnir3Z1eJPD82d4AQfqqCSc
/oprcXlSzwR5Jk8VnbEsygZGWTvQPi42OcoofufJZ9VEk/13gqdWuKgwPbSKqvzl
JA4qwOiXwp2QBCno8ZMJz4NAC7r9pqRCnTEZwwKNVlgTTbgDlqxg7ofTfNe/e3rT
yUHi5IXvYujmimvJh8oYptiu76Ih4CzVO/6yyFzCHUNg1ai6J+iM5NeUFR3YaFjQ
oZa2hgrqoBXmTbTvO/ZOG7Jh7+Dy/jZVAur1Ug8fShHg/Rogd7iyL45qw+JHvEzh
Jc/kQfCM601uKY4QTyNqGwvcvOsTbw/aSFDJiUxmj63uBJjn8L/q0a6SfkeXO5cE
oAdg+0f/E6RkP5e0oPHTc0jnMKWby2z3yRvbJqCN+WP/2ghmRnmkw4ylh0DzWhsz
DQwvQfjw0n4PaVEF3C715Pb/LZAsTSnzdiA8I5cAGvzXuRcqL6KKE41aYibmrqIc
roLJkiiq+gizCZEV0mj0VjWH8U7yXljcRIbQzDMma6L9a17N8zspPiOc6cOXzD3V
tAVpIJAE5pqZnUc4tNVwVtxD0iXEkDtsrfxSfj+epVAFEyxYzKMig6oOxLK1ZogG
s+32ziGDvbThszDaA8+xCtZP/f5SHiTa6sUKOus9v/ZaOJGPh0Wsf3YAtnfmICeM
JxEqj3cTqhuBETVKIpxjY2kjDHsc1D4BkWa6gCyNAZzueXZWaf5bqWnoMnUSU1fL
Wphnp5reNlsbu1ND6XBwESlqRHkeMYYZEsM+bVtfAWJ/bM06U8I1gvlI8rXW8Ra5
OrM5Pc7iZZsJrKvqmpgwqfSVu1psbr0ZpfyJBSWAqvNXMOAkkocCkRf4Gf8/Pxvd
EFigUchW4RzmZval6RTJ2niRJMkB94NPjYVKBs63a93jqBrnlwPeGRtLDmv4754O
Hw7W68Nt5sSs7nXIfA3TgGyUQoHW11FwE2LVCVMsiV/fDhUCxzMRZvwzX/Hdz/TI
GiB3FrENlLyctYU4T1AQRwHtZoubapaKlskUNya6oC/kmzqrGzFoT1wLLii/hLTF
meK0pgc60/ilijavjEW7VCjo14fm7Bs0UBW+D0lDHEis2Napz3oBrBqJicLqV0CO
xZuKJK12jpnqW/GKSO2gsw6q3xI82VLAjdmRufZXuOZkgNf/0HBsUCUc0eqcey3w
SnlqJw2a3TJsNCJ+LUkHHvTlnT1+9G6HH7ju5AXP6EttNM1EX53oHwdKuoqjdJj2
cvXTZW72lkkgDk1WNj2ey4kkez15Z/jyKDS8WiTbf5SvT93pKc5a1xfhsLbc235i
qJyaOom/RAUpLUC4OWnEunklmzDwStKLiv9QGWtx17XjgpednyEcVLOrBlsz/Bc6
sFfWyYlnFOlhrpawpbJrYOypeQ7+/bZCR2vt1yRxWzX8cV8yVEKyazwTHVTk4Ej/
z8rlcfxvM2l9THUuQ150xYewVu0DGVpA+IaNwUuapWvGoQ8oJQTcgs+2qSy5W9d8
CxMnIUJITZgnbiD87tu4IKWUt00FAQQBRKj1rECAodHVNFxw/c7dM5fE6RRuztnJ
SazSvcrtxQ6Bu1QAu4A0WZyMY+JL2ppLvMMIyZ8ZZymDnVfTCnzO9aq0k3IAPfsS
0vCnDIUl5dODFcMt85g4/yf4t5Se8ELXDO8LHQk/jRaEmPaISX2LelHLhrllN1Q7
j0VdzLUUGn8yI/sA2c6jjG+eb+lrCV9VSvltInE/5uikqjeAXfRzXWLc9xBXC54O
iP8POixdqXPV2tneL2dKaQZGHyD+Urc9D9KrB+TBm6pKYTy0NEuFMnXLMzbloDxQ
xvi0dHebncKy4KkGRMkyvpWbSQWCX/hrriGyQOx38HA16esUIn0rjZ8vIsaARr8N
f/ussXbTA2Jnqejo3SfkN6GXZPWlO7P3cwz8cBwVEKKJsaoNcaDtv0e9IH7q1LG6
N4KT3lYSfHUpVE/To+y6zuE/lG9rXPz8b4pJAPqob9M4a43BVgMsFccxwW1fJO8q
9fguRAApIRotNahQy0r21tbs1KrAc+gMvGLne1YDyviE9eCf4j5gkK64fyfDcC4q
66wCTm8dnM4DKRy8ICTKcvZGnUs60JsrtxMYxBwOtX81ggN5qhYXVqPh7zUcZtyJ
V97b5ehTkRL0P5XHJJ9VkaFVd6onjIl6/AVTRqvaqzwi1iMosXKMp43UmdYZH1gR
CZydrZdLNmmx4UnWLQHnZ29YRga0sgVat6X6euHO2O7zDsAs16G4QFnMA4nsUM95
/CvepIX+3RnyrBqdSLvCE/Iiubx3RCiRnRnQwwzInhAqi50wXVxUEY/4RJMp/Lkb
3KdI+HPIwndxKDg+6MtVOZEsYN4OdD7kpQogoPBuxrabUkoWZ4kXKexoNGbUuM4U
d7FkAncE/kqbzVioOrNok4YPhI9wZd5wk6X/nRosZ02c+jNDeyu+H73IYJbicJBu
dZd2ZllzRuFWedTX83+apP6MEdbmgz03VkXlSM06YA1NCWpxxT6lO+taTFT+7Ezo
lKqkWRGtAHopjMeZzyBfAxME/kgaBU8+6LCHrnm2cgjr1xQ4BxICsVkAVeYhbs+s
cu8oYB8lgYPOGlqlKSs/hAiKnnCne3WxlQQlxsZc+8nYpR2M8dIaZ+0FqYxR71SC
4DwGf8UosqbM5xJMQOjrt4p2tUz8vTtzlc0fC2TqNokdffRLnmPuTN166K5qNlHx
HRgXzx7Kg4NKDO1RZ8uUOT0a5WOgJNOOUvv/CfAewUb85aPSrI6IrqZ71aXIjrXH
PaBlBQr5lX+L2Kby2BERfrvDkI3hJb3N2tqWuY/E7LRQ9lwUoX8GLI7OTWl0aK5D
DU/4TkjFEmtrUjz81A2YVomGhfS50RGXHbr9zPRQGjAD6U1w/WyZunj1C0WIdQ/z
kMr2mnOzIM7hotSe4AIdG22V0YX+Hyg2aTOxCSssntSmOnw9R9PY/I8gb/nOfoF7
zXwiBNwGMFWtPLKhthGDcd/Ol5BmuwTmVRMLYV2EXoKyah8JP2iYPexLQIQCotvp
I1PjzftJOH/lcSrud99zpPEM06yd2FA4WlcvwkA8p5N4YqxHNY+MDSjQws5uauH/
kd6q2qX/T5tXwoei3XKZCFu+tg/Uf62R64hm7bJ8Eg9MUls8Auzd3Ydae0VPygbq
wTK6hxnmJ0F4RPwww4Q1AeEs8XywWJzOQNMcXzAYltp7Y6xVlNGRXQZGV+5YNCpX
3IpSFoUwLvglXtv+WdrfxCHyL/F229PDOwutYTyWyDPFh4yR0q409HUxEFQhsI2f
cUdPYD92BCLU8P0z+p8JylbPmrWVj9Ah7IzasnPrVuMDlN66daLfWnjKwBKlZ++W
YjdclDPK1TMloGC64Q2Fq8Ay3nVsF9WGuEwgHZAzooi/xl9500zwX5eGuoxCmRx8
+2/Tkq09HXbaZA1XiRFYXwGLYeNkYaBh+83h6KUCOJFhHVyUjwglhkUIU1XpZA5i
7QqBpFPLSaZZ9r03a34xf1+RN7W6rTeNWzkBvwH1gjy9siy/w9w76R1ZqVSgLE58
JK5CNU7l5uA00Dy17zjw7ssIq+JO17GyejbngCnanbQkTEW1qq/Mh+dcoCinnXyZ
ZAi9Tz3cIhr8ZxFoVTAwYxBDH+MkLHnJGgypx0PkX1tFj18iLsIF7yxxZC2RSn0J
q5FuApjR5jQJdL52gE9wefNkSxqskjuiDzGLqlpLwahdBawqW+ydv6qBHAuPIiQK
jOmVU1eg4PJNU/pWtGPnXA59vtCVnkgqbRlrEvPIQI8kRuoecRi01FwkKzDvIGS/
9ojIMsLM7oOCXlha9qT8k9hTOpZguDb3dj7XSrJ1h3F6SEkUUie/ssbCPrhNcHaq
DSegsRTXktmSV5BrKUn/tw6C1sLF1weV7Z4uRL8k8WuF+4TdabMu5lTQ1WYvsPn/
dkfeNv7hlppPt8qhSqh1wl1TjonFagGjvOFwwjq7vvVZvFzv39fU0zsoi4uXp+g0
1k9IzYu/QlOaxdSkrHnGJ9PrqcvCrJoGhKKGLiIButv3Cqb69rJOrq0JaoWLJNYx
okdH3lMx+Hn+hGgava2daIVGMRUXGTzy5OH+2Oi9XClTLRqrZrA5tnEChKAf8CAL
+DsShJITPwVaixSOyjMv+RnkW5d+Rm9StKz1WK5p3RD+clzXQnc1h8xIT8xaFJZl
+4xxAY7OktSgvYK/OSE5fMhGOFPg4HmovL6gM8hrYuMlaXUe9sjFnnp4y7BWJk5y
HqhcU7EwPOzh6AMUEf/ADc+SN+sxHqz2SqWgzhqMBgbBG//02JJriyNbKAiaQNkY
aKc76ig9l0Ap3rVyktb7O8WPrn3b/RHFyFULDiNYe3bpG0t7eDHlu7E8Y/J8WU2y
EzimM1fVPEnLUrgmohZv5R/4/d16uW3VUYk61KiDg3nc8siB57BFeuWZOwPDgLyV
Xr+5cDipa4qqhAmvxIA6ONzmHotthydPsaiHPxCN77Sobf9dNsuPD8zsqMQMhjMx
4Ab3OOcJ/6mn3EsJ06Eq4PIrNp4RXOZKVadJ+jJ3gpHANGEbvExiWL7D3wILHmwN
hyvcurnzteDLXfm5gHjeUXFlZFirceAvnxBi2usMiO7dWmNHQ51QknMF6Sah4U/e
gv9r1r2BYOYNHMXBOCs4u5O8e8tgCx8OC4zM4z9KNxsymRXvrYBRy1wlyPqoEyec
1fNrHaGqnyAr8T12MRPSfFueVQjSoRaB8l/vsCxMEkjZIwctTDibQG3OTkzFIiIn
HXHqev0e1JwvGzPcvAVbnampRCrjXrdbV3CnjOGkALC275biUY4ikO7My8rKtiHR
4yJw4YNRQ4UZarZlOrxXnOIXlA/Ani++f7r0LjFDgKj7o0F/LteDlCvV1iKW2I5R
Tv1xEUpURR2WPB2IppV3xJVbPUjU9w1Ez1CRFg7IUpnJN4OfGVuLjD91xjFFUdGY
PM/3ZAsRxzQE+NCbUKRaRqZyB+41RrQv4On4Yo3R60+9uza77+Gd/R4G0KhuNycA
9uboZjWVPUTO2QTRTHs8wvRFreCOyuTKXE8cqBzylf7i1WuuXagX9ARYXNSZHS7T
ax2rrO4PCtFpyOGV0EQwHnnQqwp3ETwhLyX3ob3q9eYsSiYwsYl6Rq8vNdpayWgY
jBAH/G8J5K7LR0zEFDg4YxQa8gAZArTDcN/VmH5+3vdZvTRvJz7PUYoQjERnSoGC
WTnDvgBTtk76DrNEGR6xzPJO3zELFPo/fWjiPTIvq8mI2NF3Nw6SWMd4lIQcvowJ
UGADI0HzQAwbFLOdy95Bri7tWzo4Loj4njcKNQX/a3pPCHEXN3W6y3tLdx0RN+DN
H6FX0q7gNYY+64OWEhZtbbAivuKxQef8+3FlBYF2LmtLgEQN62bYeswdJ6MNkMBq
5GyWnU51yXKI2OhOeiVvvajsU9fmuUedCzvmuBAsAg9gxBsNgtYT1XXLesOJTvCs
oXesG21kLGPbc+2VyY0p7RO5f3hf6YNIeAHCzw7RGlsTYUU99+AJlO5q4LngpfqX
Xivu+ZUXZzxtNekfFVq8OlxXv+QraAWxbELoHr1tJBEHBX2KUJo9zp6GKpxfCWOi
Ole+iqXp2yVmS/bn05hkNQS1j4SYtEqWh7Bowl6XCLUQSl2jxTk7nNjT3HSZXSch
gYqvlITtaf9+gvVoE2y1R0e/bydGRVDMVCyec19S7AR8j50zZnkilDEgA4NOilKc
NtXDJ/7+AtXY42A8VzeZP8lmtNA1nSB128qNBTKpaM9tGiqNdKnGLPOggUUvcWUb
Fa6aSTsfDwQnHREMyvQqOdseUXK9sfhAqZ1JfnQHCO93dIR/DnxJapIKiChxW3EZ
Al9crTw231HfcO4Dn6eLvEAQjROBDujK/sPaP+RRaf2L598WcgG8BPXQj10Z5wRm
20FKasZRjvgVhOmCp3p13mKvnwHMq5B+9IAlHMUvH6Zl2h6eIHdRbyegXAmrnuR4
pVXMNBsFkrF051eYplxirN5kWHcG6FkQOxXRW6DcQQ9AXzz8/bEXjrxouCV/CuC9
kYG3NA+d5NEFhX3IVZ97XR8n0DAKNjCy8sE4SpQlfN35v85mCHE8pnXK2+lnHc0k
pjd9XlXvueWuohuT1u8XRh5N2cZjwJ9SUgKfc4hEzi1wpID1kXVnFuKPhVv5n2cp
hz9znXWqiGFZO/BDVo+eLjNKxuP/4T2HDkS59eL8f0ImawZnSRUnJqCyxpmpE6rv
oVqk8Pebl8SDVrcuylA7xuaHqqYkvlDhcnKTNUxH+UqF5BEmG6pVVf7v/14t3g6M
7D6nKeflRfjKhXtfcaa/CdWtK4F0gXlY0G/3uuVDxBkHe/cmWOMNuiDR0A13l/Le
PYZwOP+JqzB/JJLNNyCCdSLcgS4/qbU3nyXk9K/9SE5rVHj2N80l1xMpQGHz2Jnk
IwAnoKBZEgIurJNIm90hE+K4F7O42ci1873BtcDLVXizmFHjYsBA04taTcA2n1RS
ZT3K2PLBTJ5znf77rfUksAEOC+3/2s+pisR2HxGqBQRhYabEj6tRxfJU4waBhpMc
NnbmGYIAkpp/ngijCe720JE/ZFDZtPM5ZcEMIB38u+rDqWo7axr7X/X2Gfy1DMJi
GyOhP/b/QSp5nH84oKYY1qPYxM+pDY6eF/Enx/8UGE460PH2QhKrm6yBMypHP3+m
Q3TBD6CGwr6JTvEeZ4ak9PDKsQq0MNskZf3EDdKXCBGbyecrHbKO/sIlWm0Pusdh
kuk8uKhIdasFnTDaRVJltCsIETsMIxNcCpTJAtw3964Wh1eGjXIQijZ3tSWCxpbE
NltphxC00Xxdgqt5lYVO55JN25BygfLpxeM19BFyNDjAOhYpAOWuyaln7GwAnSHf
++CnuX3PcDbw/nQgRCLa5ZpfvMehMAiAG7mEyp4IEKXkLdHW9s5Kkfls+2lWI7ym
oQcCARY6PNuljp0f9pCBBG+Xek9W0hNFjnq3jO+VoZwpE1Cy0b43wmFgLFZl/I9g
otuY/ADc/e4gQD2difhtCLL+Bd9UaqWAmwRlTg+p2rZfEad+bGnuNIt7NFDOzznv
g/wBjfhimInETrOVcf6i/4UwcTEDnsktuYuW1bTQT8W7+jUU4qbjy2Zqo6XFSjIM
OLpMg8wl19YRpXxlhEi9jVW1TpVP2+hNq6HO4vqR790ypXtoVa9eWruvE3laAnf6
GWTnqL4lOj+7apvAXwUwMi/XhHPWmlEcYxH3WVLr+7AE2vmtVPXo6HiqmyLWgBcp
0FhTbRAnXDkQzTLRFO6bi8P2tQfMA4ZEC8qngZkzJIxJKdnrSCKew8VEOHyakMSE
EXMuPbWv3aaodq56Xygt4FaG41aD72GlQ3vJh4pa3VIm59elqr92z8tiEwgMDUXt
6Z2L7d5b2TcMWa0BM+QQcRQ5Dstn7mCEadCBqevFvIPulsRTfAi35QsvjqUBQw6P
jb4LMds0/+q/xv/pw0TyahCqimBBI8Zc31tJMC/TfDxWI2yH86UV4WfeRYdT1CXJ
KxXPYh5AmruWCSRwmAaMFUxULqex9QEXA4xJqzwD088XNXLmX+aHaJ/82Drl0+X7
LIkQjxuAIJ21ijEjKCbAO0meeMhBduYhLbezxOuXzgCNSmR6e08Dh/34nMD+DVhU
OfK9E1+wZJOaIgPh2grw68x6xQyLUHfrGOEfeMBl7VdLauDxYsYyQ+Qj2hOdComz
QH6SUL9fzUdcueZsGWLZRnhn4pymBVBFpAvpJ3v/3cmT4cUtnMJBwcPBR5f/IER9
HuSq1UbEADi65StiaShn71/qNrin1Z2iK946yy7Z6UJo025BEu4ItHhEdQaeFDo4
CCMV+/av5WCNSMWTkiKkqvwPvZcBUA7mYaARQeDeofvu5554vBigAp9A4cqhhXmb
zb0XTh75LrRUBqlpHNeCZYqiL/rjqnpyIhW3iaGRSCB1D3Y5oAUwO7pqDLHUYhOO
AgybXiG0woQ4GyzyGsXljhs28ZVHzrw156Mh0+XcZQ019pZSvMMZL3nGnFGQuxwU
Lcy+wQFX/Ewd2422nNIEUIl0+DUCylfknvbEgFGcbV+jxjZQg96Rv/Y4mFIdDsCh
nvhjW+erd/OouDfWtVdWAkG01/93SEYrAgyw1qgEJLi+ec6rxh90+XkcYcPaWkSU
WMr2RVZ7xayULQ01FjYKbp6yJZDSQt03HcYUMnCAG1KPZ/rR7WWfI7/KmjQukbfi
pe/xap6yw8+ewGT5sHAsgIh46mUPFhMkSUpQT1J4yV4xPfi4mD0AX+3gwG/UwawD
A1QGK70PFcA4d1FKOktKQhFN3ZZ0W/k0tmB3EvNytUyimyFo8qPag3YAaQdGw4uC
njK+GARiuxSTiMMyNXoswcafPUPGGMBlQJislGlNSSNzbiKLxEGRHs9b124qdNHH
RRYz5FdTPuLQFl5/+cMg9G3pio1JbTZQD0vVJrmmLNS0n3OocE/kl8W6oGrCnhO1
aB2m4WzcUKPpdrmoCd5W9FC9xI4xitMRnKOCowiNvS+dnCyHPP5s2kB1PJ4yRE2w
8ERqaKBMoao+UYm+lLpAh32CyFjaEtzkPfaFuDGkA3/spJ2U/0CfCk2WLAbVZIBW
wTaWvZZO5MU2l7O4tsRvtm8Csn00vJwsPCwZzHBmNgDKBw7as4N/hPZElaQ2/knD
D0JkPvtyNxx+oqBptnH024oXM7RULYg+lpo4gWUyF6MAzjERRQQoSzdFCSao1Asq
5svTucnrykeVHPSYRvg1DkJ/r+tXkjTPf0xrtGh0MzEGPEldl0ETNdL47GzWLMbt
2WjnUSy/jwep5I5tceenObRJGXhXVLXpW8xx0hGPnFrJmrIkNIOFzb9Zm1Tr7UJp
YE6DN9Hkza+HEwa4HTJjlVKkcoM5d2O3SImpwhiX/2XvE549vylqSMwwnS7ByNcJ
ovxcqQJAmNWo+z7Oph5yb7o4PV4OD/W7keSR8JuTIua7Ml0hkfYuJb0+VHvn4uGE
lJ4fiVP09qbiFFehXo35+dQg4lHS22ajjzzwB9Ednr7Lnc3+iBG1RNgiU/9jlLOt
4DE8zsWf6OYIt3LeRk7162IXzQDQHmBWn/HaWKxwWSQKrRYZXcuOm5OL+TusUYL+
TMmR3sug7pELfGGSwWlK+coWWfWnRgGkMIUaVlYJKKOY+CCKMVhdMf76hcmKgU8W
FMpUPGbRgzqpXLz9sUukHCSF717j89x7WLWM0a2Kw691WYBm2oXgQgDm8nsPX3hP
wM2IEZb+SV5g17z3wv930ajaN/3pOqOXtoLoBc9j/n2H3/HULyhiKJ5pi4zISk55
0iVPWQ8mjvbUTJ6ia537/8//RwI7nn9A3rJcnqQ4YnYUjFq8KgsIeIPwz8msWwRw
2Tm69T2ta7BbbI9OwZ71CEnKbZP/oEJ8Fn9AMQ32BpuK3Bbefcc9b+e1O02M+MxW
zMKsVDbQdfKmm8YcoiTachCHSp6MPBXqWOquymF6KeFfx+YnI0cYCjtkeBnBUQze
vvtsB73SJNVPKlXdOt5G7Yt9+wfjfSmb+21LWcQRsgoxA1ChpTDCyxCpAhxL6ch5
bdyEyP6baaURjtc2XlfKCCDYE1cFb/B931fkP1LQ1U6g3PCJtHT97Ogl/rGL73mn
8crpbMF04tUg04OeJqcps4ST6lpq9kIQO2gMN1EbzRd1G686x4SwJKL1WrkgKflj
XhVINNmqfwZWHnE67pKk+Trbxwu1VpVVK/BYunyMtNbJfO7r6yY/d1uSa2EvKSiI
gWT/X6tm5+2jpIF0DABjC8+kRlfcpY6CWxWVKCfhYTFi2jS7/tbrxXAkFIzoB9c2
R5yNBrW1Ewf61W63/bRPZEUdtSrh5p/RsHqjMy1/CywaSD+oNnEWZtulwpIJXvMx
j26dXUuKHKfkNG3FDAsmuF2eUhFtLgpCtH1jjXJG3nfTEy4gDuM+wodlJVNkLoC0
jn6DDSAYTSKrbCMuK82MbkBEec91HcsCacfkx277hro/V9y6tEftbCyCRJ9Y5yaU
PnGSumr82urpsAv2cjArsi6XIe2Z8m7D0kdN3Cl+FqEzTX3hxlnzqS55E6MRVXr/
hnbJoxTeGdPxZbNKIYgasUgTF/1hwl1Mzv7U4cpaPzz++UJgut2af4c4ekRIiFCx
D1QDs0xJvUbXuuy4xzt8Tw9x9sG8Cenhod3sn6UWQzUqGMigIRfMq5zVA3c8B22d
EgnPwroAU1gAa7M5/FMCDs3OVNCUnTrSpPCgPfguwVrEDgkquKsbuxdQlgiI4Ggv
SpXZ+mto6RkVR0+clgX4s/rjy1y4o4sLkpFG1ecewTpvZk2mZ7OumSMzh77o/TnD
Dli4A+kXDvP9iWpmRDwxeyQooFpQr8o0wyi+Bi31/zmsyTnvOh4x7njjJzwRAiaK
VGfVAbXx3/3dgxPvtCYd41mlEJQwpVrTgEZjubxWKcFmpqTYagUgQQPsf65QbaOh
wKGbWbib11EjozZIy6t+oymwP2vqV9tvnzh1QATuy5Gi6zyWUqBNYMlzADicUFwG
mloeiNKCBAUH6IKfpDMrrBZuWwno78NhBvRXPail1gnRijmuPjG8/PKiqIWK1oRI
aOPYaUn2NzYLL+U7QCe7mkZk55C4bxR+v0wLvBMp112TRqtDCWd6uIQPQuHChBV4
aQv7LSkXxXhhl3S5LQwhQrYTf+j1c98ms3dVxy7y+SK44oKMW+peedsr70IC+gub
8Z4ZfCPAjfggjxEuXEss0v4RC5H4d5MV71eX4OMHAcv3LY44ttMKdTgv6HdI5icY
YaaHpTmnMrAbdPbMh0MOxvfM3Z3Fv/wSZhz/+vRAoXMqQ9R5bdagdDir/VnnA8Q8
RMFo/n5eRyzvXVxNnYsqMRM/pREDIUACIIm64llaXCHXM/C6zv7JVRk+HEYpW6Fh
cjn0ze/HuOQl49+bdnqXU9qqLY7AT4vD7Y1IxznwqWBViD7NDuVb2hp5Xr36Rbuc
LSnBP58Q0R4Qp8wiTpSJDeJwzkhghGCPwibRSczJbynORBIhUF88eYN4sRCrun+N
XCc1X+no+8hfZWZaCNdjGDgRevpHg2YG0UFj0pJCXGuYmJQfNc1tv+tsWfNhRR1I
ImAY2E1zInURw42xABmptwZD2tDJe2c1YJndn0UZ+N1Vn6wTdJgRV52anNeCEJm8
ygneaF5fjL6RVfyQ7U+P6oMpLdDZmAp5zTatelq7GNVn+yrEGY+vgYXn7qB2Fwsa
+7tU8qSajmukZYtANJ0L+V1lAlOyhRUiQ2n3LrhWpG+1kAzxrX02vJI598LgTkQh
bHnt9qIaOuRL9makNnXvzFLLheFnPszJh1PuEXH+J0ZMopS/hqRLZ5+e1rOq53DP
Ef7fL8/oVzz9OTp6BHK/EafTYQVjf2Ntln105CjLkNB3bMN+8RnMBUQXE3J8VOex
rJwMPvA1YovratD/pqswlCxB0BvOvVP2jz+1IzaNWPRGy6zRz1fFQz3TYGVXZ89j
lthaluYJVgnTRtzpopxuKKJipr+BuQvBy+s9NVBtukYGg2fZB91mKlLECd8UlvmC
0rFD/hfL8urEupRUXUO2yP4q6Pb7hY/rMkq380cxGNHMUF40cl44DAFCIx6AuIT3
JGXIjhh5pICdt8ziqfrZGZeavpku06fGObR+TFdW9jqFYvSITay0lJLFRbPsZjvI
+3p9BJa+dX8DcMhzb8JBUBv9oIG5/d0aVSyTR2juS72BSN3wf1rnl2GSwUdMnxyU
YUtBEJxziM0JX2pYPoS5nRx6eHMPmiYJNh8v/2szEnWacD4yiXZAiJD6RgKsXedB
9j8PKc8JBJ0PiuIQ7lhqsLCgHwDtFMcvH9mxg0sh4Y3cMBKoFjtDncLIRGoFpVmH
gBaercrtw6Nfy250mCSImguZp4D3N+ppg9mzmeuGpb0vcAUyNjrpYfoXf3zLUeHQ
o3I0wPXncbGToa0t2r2SxWDCDaHLIwRpSBX9WCdleJEX5MdNzvkUwT3kGSoLz4sj
tWe0Lkaeud8Rxi0im99DjpzXBKnRVMkQ0pJg61Dv1lS1V8kJOJiA2TQOaJfs2zq9
29BjqucG0KLwU0XDSQ9qklNi9lMQUh0S/KxSZX2JsILXJ5RaEEHnVd3xrXjkwTj2
WD6gNsiByLpKvY1uTPrHk35LZAJ9P5uRzVWSvU560iFNa7sfDBhcXz5j5Itm+C95
4it2DKA0MsrKnfkE8L4r4QC/o9HpL2gDaFhONB1dORgPNU/qKWXC+34e+j8Y35d+
IppwVf9q6BPNO8PvSPlJQ75l0nQcNqB72zBygZ83No3n4/Q8PgIruQIbTa6nFWXr
vscJHtSxwhGZmSLOKoiaCmKfq9FsHgeLQZ3yABhMdnq9nmn+LhdOvZhtccUtZESM
xW5vDTlz7xT8tFR2rimQvfd0ODe4mM8oKoDOeGjiMIfbFRCBEdeN50RRcVWF3rV3
4bEPEqeLYg7YEt1ZJ5Xpuym6gDRRYARCpPWsAM2Jnu7vsRcKan6axzm5od3xljhd
Ey9ZoF3jMaswNuWlggVbyWB0AzYKDHWG+NiyD2KqErD0ep2rgdRyUiPYxd7zDTSs
B80oF2M3FPzd2rMzk26toVqIvZSSiMqLucuRwdIRP+vP02jvZR0fuhPVQvO1sb3d
KXuW6hcI37TESYWEKd4Ry/iN2vva40rFeYXKmRTX99buZZYDSVSvzWEFcTc6hzhc
fnE/MwkHommwkqhkq2nfaWer12heqpl44GHduH2fmwiWJ+N3E7496B0VUfEUWFrG
UZdPkDntPcXTZxlj4tlH+WrfmJGVxo0f7wwRg/GQNUg5BzOO8TXgTftzM2oCxPU1
T//rE+FB/74A2LynTKLzmVZQrPNpHNtM9jjbRcCulGtIG0qZVWzgGk+8Ttk6FxNJ
rXiKf14ApKNW1OLjMIFAyf/kM1tPSBbHGWMBe2/aoWBOy3RfcOwrR61VvSobcs1Y
qAx8jNXsK/TwaDDQCHWWL+Cj9ZTKp4cM4wk0t4kALdWimPByqTLEiJJi+GjWyXj/
TOT16xcvcl/yOHopdfG4KNZX2FFGWlLGiGTbMA2YfGMaicG65n2wUHRPSJEC9Oqj
l89dZCpzaqbqcN6wfkF3YtKIiNCBIrqZfqjZzoWCfaLfDVVXivEm/HRQY9wxdb/u
jf7177RVacDxuT+/g0FfvCUQU5Ka5jIFSgptBUQxMIMhjQSCpV9eajOiqcGsUdua
M5U4Jx96RNvi7rhljUc4St1RsCcok54uWDXShnjztPjM79IP2IxSEdT+HMuZOfNB
W6N8ooEM8jdlRxVAkgBz7Hg4iEO03AkujTfEWe1SW0gmgFzAIJoS0zoZyevDXYOK
+rygw4QQrOpMFGde1i4Ows2qoBfCq5cH/xJ5ZlQmi3tLFbmk/IEuEHULi1X+Woh3
fXu6mYgFp+wmA+khaTiZo9ujEiTIeURUMtQAKZBwKqyBm5dwgQP+RWkbsBPphoiJ
AFA5vQqGNwDo/Bg4U0/cgcs8bbnnwTGai8qhFYCl+eHJS2I9xiiyVYGRyleZS28p
TRzXv0ILT6NS0mPygmv/DJE5JbZP3XaWNlGq2vCOWN8JuzQ3I64hvQVGibAibAhH
gPdFvkYm2lOftW6uEHkI4bUeINeYu3dI4PvM9MWkKN/mGR7NReJKk9VoaQSymnWz
2hMF5cJurLqW6aUjuLHelHeLPlI+MJSnE/CD3fdOVpqglc8SSvk/nz/MpuXqym3h
D1Je84paywxK9cyS9+V2em6jq8da7KuIcUn5Y88qY4ipvYE+5NCCJ1amKtdwtWYg
n5yJA4fcvTN8gawiMdqYMhYqWmSRpJFOdknrrrCjmIexZci3amFV6iQpymwnG/dG
DECt+WyPu34upnjsxC+vQONIuV4ryVKz1wzgh6mtkPJTcOyP78BYEwS7/VPrIqkX
W2a58+zozifH1GWvIu6vj9ahW7hoZmNAvjSc1gQbiqVCYSTV/RUtshFOwNwT4Oyt
tjW4FZFSmbR7nVUh5/9qgi1h4zmgKc4AnN9ennuTKLVWlYEDbHspTMb5xeTS2JeZ
mKwuec2rbbxjJeNL1dEayoIDB+38j8+EHrKZxy+noDyJliPswBV/sVEswe8vHkBi
HzWo+/kIoMAm5NnUKC5NI5XMuYY5FBWFZHlEM5dPls4lBq74zVnEpnM2lKxDC0F7
FFFmqmFRyJBITn5sbH/sxyBmr4ZXhL/rzE/14rK0js15sNqIcdezhtmne6uAV1To
BlfT8/kM30hgfO5ASBtqVXV9GX7T6kyNjpehBEi/WfS+2NDEwGzvp/tJai6YOBNh
StNOYhaH1VaHFdNQHXAXiHBvaAwEObpJRwRQRzlwFcp4pBmodTiv6XHeoEqSQODk
3HY24ytCwUF+0x3hs6BKPDSo0PuU3cdIv2hMlBuH7Q2dF/FfHObMgS69Sm1nDnwU
Ph5UYNgu4c73zsh0iTITdkThPXgXyHMaLDYsaXNPkFsDKZdIjti/Qw4z9di2xe8h
U+3TTXl2QJY9NF3+gZ/6vYEXhssAoGG7EpuAcNTGJwwNcIt6bYBSBYaRtuHv15co
+IIrt4FkPpHElPvqXqQzjnPx1CIqhrssn12F5c3yUB6VxJHNV/iJjX3JqxPLxZq9
aaUxUFwjeVjj9MfPiEsXKh+5/mYaoewm1BrEP8yjJVE7lMPz5nTo09VqBgbzCHKQ
kcQlbCITGKECWI5AxUOUzaeXqhNkj9mQRHraoyxyuO2dVB1EfgaJhRHu8QJvvykK
2Ky2Wk3GALBe0T2lHtmaaGaxdX8muxYdEP2ODQOOW04/0EisHqAqH3JNXq6zeMsz
yYkiG5VKzSwcctqXZNuXvN6FW65U0JIU5Ml79PQE0Sq8HYRbl4FZavfvxhusUQMI
PqTc4nL5u0O569tcZWj6svIBmkEvtXa8QVHNlbywvemiOsVzOUbB0ag8qO9sAiDk
mi4RaGpVsXqAF9Fy4b39jf22zMcLY7bLs68INwp9J/ggRNjGO1TmFaal0gfl1LYs
GUGZJN7Hbl63PxDHgSMP4ljDCU72W6k9nNd047rQjZbI9IiSLtbnmd8k1FnNksI1
W69JvChyisbWt79VAX01qtz6a1tOSrZXWD/NE/Y2opAfGESFeJOTB8hNN79hlAG8
JCcGjEYQC+hCEQyCQ1hasJPuG9LX+1YbUSFB7qR4qNu0Bszeh2EKbNkr/1MBZGhW
K5Mty0om44GjjK7O+/Bn/VaLrIDttKBKWQQPv1spJNofgdQOoD/fRqLUHJtnfsSu
U8evf6KOZmJNbDROd+8W3bXI+kHTCFNqbzV3PtgpUWstNMKDbPdFOddxgn0+LjmW
BTfGqFlNg36vLASZIpgdY38cuLKhBv6IAvQFh1qnv/znkH6Vx9XbeFCEH/VmphID
mdFhxwDCZeLb+8+BzCJSnso8fMUILqEXbLhJckn9UZMscALSqJJfjxTEUxWP63pU
VvpCtxuCp0auZcY+a4wGgQmAuGWB9Db5OI+mH32xuNaDj7/L2ei87tw8VG27TQpo
o/LTBoVukQi5Q9ZHGPtQmiiu7i1NLObtt8HooL/W+7mmxYQqYFH3y1iUbGO7kNdN
5HzCaMUgvCiuX/gm17/PoOxOXUn5hTuQHXRMVBfH0NrFJgokBGHfzW+7OL6gmIPe
kPSwrwu5TEyaxTDhew0BNjBD/taOu7kkQkzIA7EuVI1y1fVgYqaHXJNETJa3F3Lw
R/WICB3RuiOnlcwQHR8YQQwZtITQFm9FyGdaw37H/lcX0NS4KNo9IWyi/Nbt0uzV
mRDwvS3RnRUL5pzDOP+Z0yB3Ufbc4jvY7UOJY37P5fz0hmrRTsPylW9GGgbgCV+C
IT/EnJkjJE0UN08+y8Hv3H2fj5nLaYY+V4xjo7zuvo4J7r/ya5r9gJsTKU7vWA8k
V5j1cWyQBbEpgrlVJa9PBtjwfjWYd0X85INjnWDFxhQbesCop5R+5e/qMxk7z040
QHfJoxhZPuXPHXYMUQDkqLfXeeHC04gUU+gMl+fU87eXgN5BkSnJGYPx70LT1X+/
321cA9bDGNlYdWh+WkD4M+jNG5MNLOo6fin8BbBSO+XI/r41WdAcWBhOCbbfwJmM
xe7rz9AOdGZ6jUm4Cj2e4ompXfwYaTvw/OW25THFWD74Vg9AsEFOEiOUAni97rQV
OHtBZ2P1gKJHo72GPRrdSk1wV/pTvgX/5LwOMKJORGhpxbhcUlLCxyzE3X00gSZa
VFgnkQQs9EJQVERzjneSaihUK72LCsNHoHgsN+dguVUB0UcjvEyHbWqv2B53E5Cd
OQtbK/T614Lpb/kPMjiJVC+ASYwonqBXed/D3uEgf3WhJ7naUYn7sdgEtSM3/ham
VDV03o/o07bhVeRCqtEBzu2eViG3TNKg8q/fYiWihF/QOWieuDOup5syiCnmW5ZW
5hNUG30fMKjkq6TrS6zY9rBec/x5nWDWxapRnp21ZtdRtd1Sxh3MAHvgP92oGdlA
OZhsXGgyDd7sB25lc4A4dq+ygo46anH4wjPcNNH3NBtfU4gfDJaO0bkO4HAibSKW
Rd92Uvh2RSZMKEYubhHNVDuZ5AxePoVI9nraSBz04bVU8F31nlWtnhG1VG2Fkfuk
iWDBr55KQ6OW7cu3rsyqGvhVlYAyMQzowLfRPHd1sfwfzkDZ/fz9uCpjTOXZmIQ0
erG0Nzip04SZ4VoFwxrKmVtU4raujuTCflEkRFjWQd68NdQCxkjSe000YJWqCkPz
FS9/s/6voB5ZqmpyzQorSQvwI8PPsteH8gdkzF1YkUjNKHclxRjBEO59JnOrhDH7
eW/1iISUvAjQOIDFkJXMeNfCqOl+LwGhy4UQiWw1pO999d2rWD2F39WiOxIoVTXY
qEw9JAU3ijXQbGPeu09d3y/Twvc4sfaaspDS2OC4tByaRmBl6gxojOnuJINDJeDB
Zdm5qq6pLyxGqH7fB9G94DeDIcE3fXsXj4qF0YenhRlTK+PRxY2OsDamoyA+LlW/
l+dtLD0g+V3ioXSiKHP4jWnN6UsnP4LMaPUOpLuZwgNDxCukX84f+pzZl3jVxTKc
Wt8lGkzfMKv/OlrnVtIs2Hw1xOF3LhWbvP7c7qBF+r2eiUrcJMv8R9jfo8J2tvv2
Pifw2IJiz4Ziq5/lUdEYypsCzJ5UHxT34wfgTZB0SFdCfd6J8G826mTBeymhjXkw
ynuLEgawhPo5WAuBIBKR9s/nghL6jGXvB8hl9n0H3SbPdiwJ7MQuh9eHJItU2aoS
xG8GZn35PJohIJLQIH7Goi7DvfPBMtDoPES0OVUURgMe9Wbl4RrKNkTfMSyhCOxq
lgc4nZIV9GAx7BQvTv1l70pqorxJh5gWWsOgcR44tCoNKGcwbipH9DGyHX6ntBss
K9jHRT9G90E4yZRynx7ekAUUdjben2G4Nfxl3LwHqUGJh8lM5K18zx9cpf3H218g
aFEnXJOTXwman9wWrdPnaQgRNh/z1rYdmBhDRI+JKADyD5ibredNr+UtbQr7PuUV
E0dLjOq2ovdCWqooQocaPnFACiNxi0FGB4FmulQQG1HDQDeIw6mIRxFENOsNgk8C
wB9MZfueLsdSj4RgESFJVuH+EA4DxT0e4XzdBLwjj7ArfN0VYMN+F7RkGpNjKRue
GA31TAGWM8nCdKKfp2GWil7yNg+xifu4BjQ5X2F9wWjZWPltD3HRGPAa25yjF0NA
WhoNr8Nly8j6+mOKCIHTxrGX5IJ1+6s6tPqW5lxRTY1tCyqDTFPEajWpQNTC5pAj
cGTUn2gixo7PS3TBTcz3QMGDW73dfnjuqT/h+QmWvxQGxQPGDi7NW68YkF6mroJ2
pwWD8gGLwLMHYI7tRZ3Bf9rqIw+SJwAYY/Pa3dd/NOnifYXqEHTFgjoV1psCUoZ4
7tKZ6K7ZR5WlK8HrIk+xcsosjEw1O/dbDjxR99gNpEfGSWZVWQTznOlvyb8Ml5fn
T43dez7wHutvy9g4fb3IgqtKc7EnXPhnHnBfxmbkLsvDkagG6DLUcUtA/oOWMk1Y
EV/djf71AKsa0/B2f0yzZ5Rhln2pxXaKRph6M2Jt5cXlTOHSCYkFhl/Qiv4WiXcU
eEdak3+3uWuoKM8N+2qTXEkOyYh9dYZKuQru1Bquc0np1L8mTIDUUk+36nyjbBS6
y+qoazdmd01Jg2yQYeNS0UGPXhHa4bqTKOYBDvOCXP79kUw/TcLG/6ZzkpopNmIx
GWf/874meWcQDA6rdu09gGkpXQwnsguZbKmVv75GnHqs5RrxYgPcupGZ4+v7Yx7b
+gucOjFDfZDwQbxu1F2te9dbrP8qel/w3IMM/DF08/wN70zqycYdRJEzhzyLjw4k
ZagFvRUOH22tmNe4GZD2GdqI87GgW1BrAR8V7U9oW9aoAwvSJfHZ909yA+mGvXFa
VPcq1eCN7CE2n/vgT184UYos1KOxSZoU6HjTv3V+cWiRUa3ScYqKGOfZG+TOiFrp
VzldSGrGJ6N3FiI5VxfQ/9Tx1IUKPy72WzWB7XtXoNVxtD8EBIlU1FUOlJ3nlQSK
R85ZPA9r368KS+OXtBXG4IYUEdpRSdRYoySMWe+yW5mGRDM9OrrBcx/LKSb3wGbw
sAEFoIgLjIkt83Mor/bYnll6MtCkpZssp3hkFrZn2zVp5gra86Gyl6XmlbKcYg/P
zoHXwzxJm3LEJtJiRsZ0UowPNuuYG9STshHMklilCUpw6bOBnT8y4lpRrgZjGcD4
muYmUh7xLEUBZdjKUtZNIYXz5Whvhi7ZQyc88EmWw7Qrbrw0aRa6sw6skYf2BilE
TxukjR2VzPQBaL05bNanl1TIrqz12TwylSiOAE5kbuP+4elMi8IkS8xqMurVtMdY
8St+YpcI0iTbe63OPZKuBMuA1rvpvNWefpFkXd8/nngOyiV5boBrWBjHYMEBtOVP
tFdaRFaG3ryu9yf5lPhF0LdkBofF22iSZgWr2moWdqufvL+mn9RNopb7dZlZg0B9
k0y57TYmviLPUczRtJwu5JLExZ0PPumu1j00GracWvTlLp6gPXrdhWzOxWVBE2AZ
z1cCusaahLJnd8eoA+yeo6fB7jOWBlwMmH3n9b1D23P8B5dVTK83I91ej4+SDk16
Gfd5M+B3phrKazDRcU4VKD22OIOcze4MtUfF7aV2EeX62vPJN5tBcl/Qo87P97Dp
19qnIZCtUYTeURtUZnP2C7ssvPs7URmveNUx1JsF6Dupi+TTkfV7MMxLsc9oBu0j
mBs5yjufQ/VQqaVUxPawfOpvbkhWKA9zpUsCcNHZPwst3Kly4T/Zw77i16dJO+6z
HIAlu/Rgv6anYjjhzo2cxprrg6ZTDzQbyBJTXOU5KzHZJOljU4Y2N92hcAVfI+/i
augts+pasehV/duwych/uxBPyKGD1+7E7NHpKnr2UKZ1Q39lmNueRmtHjZyMW4xW
GaGzYUyj2DSy6mmbAL4EVzxyzbhHeBxBia6rMoGjOY8pFVGjn6Yj+0B6oedvMoMj
8MZGXHQCzpoPYfr+6DGf+q0DFYJGcYfGCa+7OGekT4c4aEpFDae3SVuKze7yjX9b
w0Ues2c98s1f9RqlRO52s3XGJPx/reOTlLIaGcteHu5q0rVs4AjQpezKsQWgHpQN
mtFdZBZzKVUNDraqLTOZiTQFriNLdjbs08MoVQBsK9YK5Tq3evFkPmC29OtLsKpY
7MF1W2940AzJOdtWv004Gsln0i5se6TYgmtBYHugbw3AZceZwI8TkYXt+xPyEA+2
ukAAA2Hog22WAz+GIrQBSXrVLa/jeRJlF9d0f3c+mAc1jkV7BHzAR1FJt92jsPIw
XtCQH84gREpanvH7W4SVZChyY5hKiHpk4934qWNyfWKCnVxeAOTAM9QoGPSS/l58
0c7HzEH4pALsiMuzeOIL6QFZHTvFhD0XBL2YGuVyPy44unXFxEdUpyWswxELc3cE
ens0+YopD+z8vMb0m1aMoL6Pk9snu5DTDDbDvrnTdSzkMcwiT38u4UPWLQw5qNPJ
YhcdTdBFIM/DogjwRp/xQa16e++uW/pggNGizmntjGmj5p2TV1ud4SvaeKifhQcR
GuJ5Q4yHZXXy37LxBa8jBPPhVeIeJ6GhA42Zs21srlvprHXkcOlgXK/3ABvqDQKh
gSL1Jy2dj5F1wyCmtj6p4JDqCzz+UczJzVwOxOEKsYPN8ZWijsrNZNeioGWrW+e6
0nSev5cjKIqzwN8IUUCkXWPc8SB9G9231eo5wpdxTgSRYC5wuwTPL6d2hi+TMeCR
RkDs4QVCMKtBGV9KnTLSh1gLtgMxwV/HUZLEJoFG2DMDjzcVN3WAILsCbMqs+zNf
nLpkhY002E6hbJsNTCfa70bk7qCUyTzOFF+/kvfzNjdp5nmfZNYc92NezrqJ4Gg8
9fAmWGCs/SJnPfdLIpDlYnEvecb80oPHYSqKrnIXeAcDvy44lWG1lyZZqdeMkrfl
C0s/svCgeSHvrsCOxOTJcp3DFqa8zuUtDViFyrcmCp3eT+Df1V4tpWnVhc4T92KO
aglvSzUwX7aJEkFJq2KETZNH7P7Ok4+dYJvzzU5Oe2s=
`pragma protect end_protected
