// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ge90kmZfWQ+/U0AAlxTCMntLPAxcIesogKvDo7h2Ap4fN6eUmV/XkHjqcNOplQKP
jNVlSgpBblyS9sHA+sVj5mKFPuh8QVm6i8uzA6/2SdaByMOnBJGLbzD+lD931RFl
CDrj3rsd1N8wWf4gntewHbvIAtpm9Z6oZpuJZmJhW5M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71552)
e4OcJCp0NAURLwfVVMgT3n3g8zOCPX3TkfRSKrzGDkBgVp4hVSd7V7GmP2j02Tz6
FOsJs6rPPaJaTboXQU6UhkH6JEu4BmXvntXCvubsgSpMKqh8h+iD56AIFgpDCB13
afRKx9Sm38d4WGwvpctcptip1lLcBGVGY9jLjO86LvWhFtux56jXju8KuU/zqdRF
9JiKG1JMAZ1NPboWvz8RNVmFtFB5nDvXPmzJWFIi8Sw/pfkbCrO5D9go0/OE2Tlz
QpL6za9P3sgpnAnPptvKPFaJ8EtS4KvDj9exJd66YZLcJKfEpuriwOOFudSEiEMW
ICEp4KIW6NCehwpAeUtWLg3th19+eV4eRoWqco4PlYveJdxqLLRCTQ6iG04F5PE/
mVGjMGp88OPxgPLmAZC6uhGDo/zQ7/xNxxRf5VCiaaVg6djQV1mcDKIK/jZ4VjJV
RXMD9xfsoO8ghzIpkL3hFlDgUn/P/yVxfRuJrM2FkT5QjpKX30tKr/tQU++k1chv
GtfzweC/VmgUh+UT1FMKwmS5AgV2tdlFowBoKqSqOhPL0magcUwXO/CYiMnmhyWy
RYqC6yVpHaf6Y8vTLzSYQLm2Ymx/uBc1IRivM5Wje/AaeqEwheng1ccY6uShX8SD
VAFehV68o9S/VGOyE4wMUTspTJ0G91XgRNHrcZhy9VnS4X0w1diWWu83FQNtA2lj
4rV+uz5/c+4zYyCceTT/x/FibDjmip+VVPcVL/LbcRJncCXgV/kHbunRWH/vhf07
zmP1tGiMsb7W7/hT4VaU58C2ke7Z/PwL32neA+HgsCg8TmlgtywdzT8b7or+fs18
0y5N8G0+SficGAcHrHxzki7TdIX12OxLUgsY+1aae6ie8vFAfm5N2RQNkVPXgPdq
6Ub32jqeZ4OPTEqXumDV33ubNv7efZAJcOYOxzNnSrBlX1N6LjwK1XigTQZTa/J9
D1c43MzkOEYuncs1ShsjcrdCCV3rsYUuoWvgxaMsMJe2oCWnlAK/Aa5b5EkTt/7i
v2X/EtU67VbhL3GO8xgTyVz3wBK0eOL/BK6Yu8HFWcj9xALK2M+CdMILpHaO6/DA
JWlVNyd80qqbPLD2Xi4t70vnK+TukQ7KE+kNcgDLO/QkIcORlvRyHP2qeLrxNu+E
BLOocIO7vVfqiKNZdReUeiT5cXq3TYXAtykPFdixwWI1lqCLhE6DGORgNsk1GBsL
rea89oj9+3C871HW41LABfmw9en2reg4NWC0p0UZCkk99RxQ8t2CFuZ2WHGaxjYM
MCkZoxsU19DVm4bIYd5WEaHk8hc/FBRtei3qjwgpraiKK8TFTR6v+IFYn7B0MMJI
enqndkGV81hKLSxvJTi8Pxh8VW8YWY/zqci3kR57UOT4qXU3wsMQVcGNF0KyaoWo
ObJ7EAPCOrlAaYq0qOo2mKyS422qBlbNL/CN9ZAYK5GgzGbxk3TGjnT8oIsqrfsX
dF9tth4jTj82Bemhu0wPqN/UvrFfcv9+AL9bgY5WlJPZUyBFLdbXjSFgyJP5VD+m
C/Y72Y1364T4d91XWMrIsXvaLNzfGxwkq67H59+eHUKVaVxBzZTDOBIpqtWu3yjW
3Xw8/m8g1L/ARteadv4BH+3/bF1cAwdHMJfMlka/FXyLcHaFYn4+mPg+Tb4Jvoil
+Z+gbPQrHpyrg0tD4ATRy1YQl4k3Tse2/ziGO8oQNu7koS/SX3XDJNzob/qf3T/N
U1B2bHMpIXoCDvZhkyIKnZ2xVE0LYRMJg3yMkA/RYtPlDGJFh0bsKmqUyT1jZ2XG
wAtSdCrRfjX9zhfKzdwIPXfrRMztvnE7bmIo2ExXnNPClnIArdLKdHBzcxY/Dbgb
Zh+xci9Ag11pc0gVMtkdObqKJrI4AIWWPEuS1X6YYI9Wibs85ch67RrXacF3nzBL
U77prFIZgGkni4+tC4Ah8HM8DjByTklXFFALlLxh1Tmdlq65iVRXwZHPvRWNM/5L
doTtSKA9iUYLvwvMhM6snOnofFJegPDe6Zg+/5Jwq7mpqvMdaSIzZOQJwGttUVPP
R8ARDLEqH8IsIOxa4VfFMiEt9i6/YPGSiWbG8oUUzytqJ2ytchNw0F4bnro5ouTI
6QCBCNpt2lhTSmItdOvQV4CefdSlM3UdvxAv2v1SeGUEtgF4bSXmQIISPzQK2K+5
sYHu/EyhKLhw2IUN8U2EY29gTT7roKvKKqyNYToGwX5frf0DVxEBXmOz1GgT3WIG
RCF6p/FXkbcxBHksFbp9D9So7k4HaySY4ohJU+IlfFk4Ctarh5UefvY8BTF4vICU
QZwgp4soogSH3GPoqwBABMIPEVjKCHKozgmwRd9o4djL54a5mK2URtNrYIwVG2MU
rAcHuzFPKhi8nW5CFyGJT9jjzy6u35DBQsbo6NGQkZMcdlEUw6MCq+UpzmWXmcuv
1zjiEeXOgc/5c/d0UauVOm4EpBGST3LgrT3YzsdjbVwhXLqfoREoYADNVwefj5dO
L1e169k0Wf6O6x38Nu7o9u6Stb17OXXZ6aRfDPyEi8mOq7c5SvLI8l4mXXdCIbqq
vsknPVAxmunIq3t7k+04UbWzIjP1Y7qBI0CbjwU72JkdUNOcTOzzPdj6l6tTWFuG
2eQ3rgK6u39TDlizJprnj1hEGlRIM2/MIJ6WWpPUUJYBTtkxIBCLKlGVjZVnGbJ8
vuqta/IymPRLX7Yh8VdZmZIpVE1WbtKzjbZ1YX2DmLBXNX/95oYJGW0CyeB5DS5B
/WK3UzHtPes5rmnwBOYBkfpYxw+avQc9BF7ifmJ8zc32i9lDuAJSKHz2kM1WCaye
6IUQ2bmwBu8Lvv+Qmk3cAw0CvVdhZatEgJYrg2a5QnUp7qKzX31ZHXuE/RXisfNj
MT4hn+nCrndISWqs42qm1EkrVQT1rOz2PnJzyFqedP9/F41wn/qXIocBBv/hKBpV
ye79tpIWjDn6Cm3Wxbs2CswpD8kzWHPtoBYp5xpQra08VavC4hYPxvXB6bUnS0Vy
j11wd9XUi0SACN/xuTRNGwsdhr4lMWfL8Y+5T2EnljPGAdxWMvcl9kuDYQdwI9CD
8/5k8/U74e6Q9mPk2lDAPfsnjPqJ0lmDmPgyBVO7TYj4MFSqW6EAjnMuEYi0OdU5
yzP8LTeR8NYWrmEn3DQ70fTT0r/38hB/bAEiv4QryqEhfeVAHMUQrFRwVvCrbdmo
LG0blymGhDPj7DPrnDFeXXErga+36EnIrFH6KDDNrekDJ2uKpUe/9wB6rYijv1HB
yLLOFT658lJ7AJCE5eDi1tE6/dqVnAXgTW07cX3MhkyuW2rNv+2xXrsT6ioXCww3
u6qFbjfmpBeBJZS40hVTw14NuPSI3TplOzhPEI1pouFHXZGR1zwW4/bKrdD+PY4A
xAyxXwjglr0Q/JsLj8KiFabd1NF5d2G08IsNW/J71dntNDwn8Hcpma3gmtPiEKH+
g7ABIcvyoXShUqhGAbS8EQ0+gOy6HnVVtuEnWs2vvqHLGp62lyx8zzHSYPJKxREJ
Rg/puQTVtAcd7KrzDk5AfkV0EWT6cbZHEBm0njA4iexk0WIEfF+ddF3KKtXlkVTn
BtBfusPWppll/Cvgi+vJlUCFyIy/9ZOwsSQB9iCYwLQgUFbT9nvYD6I9vW/nkmsN
lJryxuCjjCojk/gFjIVIU1FeVp/Ir7+sllDnvEKjMLpGMOa4df5fYe3aauDibhTU
dfyAMb4pqh4JD20eKTUqhO/a7AyivUoVQ1Pzi6kUfb9+eF8exlece9MHBnjJjF8D
D2hjVrPKNbudffBmtwgKWehYOkH1t1xmyBDNcwt/7QDMc3Zgo/7eeI43EMX7KwUX
0eAuWRUMpn24Xv+K36M8/VCb3XHqI4vBXhFm9+6kYZQJ1SZLnzRP1YEDvGZG6K78
kO762DSLB+mSNzDDJSFhaZYcj3tIQZ7eAXUPs3zA2npq89e37FRQLaSf8jSGjFuI
iS/HumddxFp6zDCVEd+llx1ARsHQTYKzhNj57UZadUVE/JYceVvxiWqDgdekkL7f
nA0e9AU/kIYODNj6VCvTioGSVQOHRLRvXu60AE9QCnI0zj/dDAHm7xn/u02vUQoJ
/FjdmN3Sc9uoM2YrweAY9UmeLpfLMCqm9jVCA3Ku1+Zk2OEcSjPqbiNsmoEpUJYJ
FUrhBDKs0HSCklot7GlumIKHnnjhNJ+ghs9dF/3ju1RYkH1ajOdxpPqUqvQyTknG
Wa3yGLF7rH8AbtAoDtIGBTm0e6oiakw4LPZTwrLJjsMy1DsBHPg1jooBS9gzoIb3
u5yJoXPTi04BFAmJIK5DVvZkyOGu4DFI+eCjn1LkLsc4LANI6SPxYTvJwvKe71TS
ghZC8/bKAHCjp45Qii2H/wYqeQk2Lp0b9sgEPTxqBhitctGgnMhoHNBuhQT1GQOY
kL/AvyYGcPzZ1v4pdhtzw2YH+V7IEz2U302I4O71EhldzrQaTKbfsB8bR+qOkLYx
Q77+1PJyUxqKHdyOOcUTixCp27dba5R8d/jHAlvOI0Zz5lh8Wm09FysUh69/YobB
lxQ2Vcs+gJw4J9MP9GITGd3an9x1vV5s1VHUy75gtCeoGN8SKn3ERGDn57Sufn/H
qedmC8BGQWftdDpOIoQAeBGbFiAfCNiGAOBDFLHMhrxR06ietNbOKbk2wytEwNe2
rY+XyiPZHmGNaF+IQQuRKZDPmEmFIvl9rG66RBsczRJsWYD0icESNiebivRg4C5m
viKbd2iu5Z/bwitoyYYwhaDVfmsDPbk/muc3HrCysNUa+OeStHj0scOPgw8RbVTx
K3lneZNDsQVehC5NiZqMbq1ecE3wzHtt6P4jNpbHaYA0hNZENcjYHkVN8tTlRwLK
Kfx8UlYq3OXnxkxqkood7P1t/VxVo/jQl8BitgwghiyGYhvgcRoKMDG3GPRkWRgO
VqwAD4YJawsCELBOIRqsmu+pRJhiSn1vmFqf2QpgJVh+06Rnksaw30n8Fj5KkqlJ
EUx2drGiLcko80tk8Q7+y0b36OOEeB8GADbFBSW8JsUsABCqhxbDYctJeqK9nSle
rXJ9v0sJUVBpBNt8kmn929vQOeuFxR5Er6vXdwBlvEUB1Bkw1IaMzulAxF5pTcUm
TmJObLxG5bmkBaPP3+QyBEsVBUGkRzZLDbwfIUsyhw44ao60NaHuUK5RnowaPn0N
Lb8cUy7KDEg1UCR6p5uZm32i/3elXLnEPkcR4dy85riKT3Z+uPezkbwNgQiIoLrZ
VR+UmODgPQYzEWvqcGLePfpqJnf7ufwt7UXJeHHK+kycl2gTQnFkdxAeNBRCy49m
LWRYxSrAP2RS+jFsISU9dEYNUNEc/cdZk/wasDsEqKjZC5fut9NyM1c6BdgsBeqY
m6VnrGocNeTdCx1BnIY6YjJs1u4/oJWECsN6D6BZb/HZtp50u4he1VmxPElNWa8g
bcKXbamILk7OZmQoI1jvx9qPdH+vuO64m23eDjqyHl4T7tlJbjybkkyXeDtzCO2c
i4+Gxm1ApaW+ANMgaKchLaUPrEnNX5PQEYfHKqQ1CrKRKmCjFxOuYc/DgvvQrJ4F
vyV6JN8Hga2217OJXXlI6mPq5CVZieXVUGThbJ13IwMrYQfwe2rPkcFaH3FOYxLW
y5ilfZ52JibW/1ViK86fdAHnKPMctbDzN944GdzzA0vCCQjBPg69Eo0aeA7Dkabf
PXTrcTtqYcMbRZxmBaBXbNSEov5Uw5SscxDuTWr5zkh+hFav8LY/NNVXXlZV+3zX
0NQxARtxkam1CVcwPR0GcDYl6salaMBFEgbAHZw2nczt+TtnyzClZKRx2IqwqbPn
W5ctGXl/PdwS7LBqj5vR04rThKoSZMBhF2raoHtO5DC8PT4W5D3fbc+4/UH/JY48
KuY78uu5GaHzzjwWOdnZVsQ/uevhI+aa5d8e5B3tu7gRWFwM6+boZrR73aemQM/L
dUHKGXwFQSI5HSRnI3bAvy79n6ycz4oJmBLAjKYyoUM38ILEnZA9r/3rD5CcI2Mt
c9G6DULFqphpznOYLRjCRTy9OV2CAMfUw0z7vbdxjGUBz5coWhbUFhgDadlcyQHl
gQ5hA2YaMh29a0eMLwOIfsUBWu+CYhDRL7Wsxms8oRmemi8eXY3PubQGoaAzodZ2
VjIbad+yXpGJtyhb7RlwIfeLun/DLsM52UjqnlJ7RnTCkxFEO2WZHsMm/147ekT5
14cZKewh4SXONW2ltJy/ahu4I+m+4EtBjuocAJI+EWoamq8xUiDpAE2L6j+HG06c
r3dXgQVdZI8gBDR/PbQTwpJImg7rI0nh8DuHKTZO22mFlDYpHU4uEeGyQuXvLkag
i46dMI0RnkScMpzB/1AGJgs2zcnnyvyPsgTl6k4jc/1owi4vNL56ljDEM5hSLZV+
F8n5g8jcQe4NWPnt/6ZwxJxjO9wI9xEEgifAWa6O6yDnZATzWslpdb1wYPCgzxhK
zZKnPkZgsmEjo/WFMp6k5k21eKgSHrqWHACTSAWRZ/S2AVlv9KAq926G2qzTELPG
o1WrOTtuqhwuhtlsgJeha5pBkz65EXoxcnOlVMe8EC7TgC2WtNNtxn/5RA/BBtJo
JrnC2F77Uquj+8eih+qQoqE1j+ChC10dY3M//IvPoCPOsRLh8DOyI8gaKDg3fZ3t
iIxafFOiapjgYb/bYF83ANmJDvjy4Q2Pb/JSH9FaRzcUelrolXH4mXayC6d9kchB
ZNeJ5OJ60vnsGgdQEHqhgVHRWuRGT6xw7J3ydmu/KqPdhVjRLQ4QYXz1A5QRQ9XK
bEBLqF+C+Cg2ncXRGN0B9hpjTvITdys4NdDWOlQ5I71n3TJL+DdMrueqNDEuQ5BD
oOYYYry83WOpBPjM++LyYxwUDas99vflObonYYVBW9V9hLoQz3Wy/SdsovQ25cuP
C6vn6MM97urf9Gp17v4JK0e1agw8ik8J8SgMrrw5kzwcjLjn7tTHZSdIYWvFWI1o
ZvdMqzjWtaw/7dZy6H/GnQ0zPoJLWHhd385MFXV9wPWjo0dnVIP9SbMxGe2hsZ0g
t+8t9fKP/7Ow2d3rC5Hackd9XBK0G1oW2gTHEX6CVuu5fYGrRdyBki9hz7quDx98
mvvniJtRiqKWhCLv+sLT+EJj2veNeZAvpOjgrPrI5XTiOoPdRrQxQ/YseB73jH0u
fEsy2aqF1N40EyzLXIjtNtiXEjFSIcWsYgmFrSSbvdq98qqv/zxPWRtKbYDhGEMi
ZGxH/bw3ZzpTNj842PLYgnIrcy8K3Y9XPVoy0ZwTnKNKbXQb7AYLG40h/hWYWvOo
eynRH/g5paX0i35mrBftD0nlPFeoLjyGY27W9y7JnOSfBMXeGNTClQsLXGfq3W0e
lytv3gMSl+tNrgwAVyC3jepP2Pg6xgoTpFYfwRSxib8gewIOF1lfDD/lMO263unm
HZZpK2QVF9EjDOryh9OI5PBQx40jTiJH93boVYFUJQsyd1vm5jkv+JvtXBrU/FeR
dJ5J5jzsP40CFWqvj31vfYnXZz2NMsKqIhOc/cfJcORKLQraqp7hGvzBTivqYIOD
RMosT9XEOgwUYGBwfpPIuCLEiiCV8K1uP74j/Pn73SwgmuHvbIVxrcfoD/bPLOwT
OjyQG40ZLQSvh0C9uNTJVoTcxS5tZj66Xc0TsyUtai+nEsmsEx2FqZqN2FVxdkja
mEaG4VgqmMWqGLbhiwQFxahN0jsYqrsZdg8VzIIsTpvT7w41mWn09NYt0vEJcHoA
kbxYbjgJWOpskcF/eMw1vEpyk0xZ8r9D2lB88Uxy9mj0tbvZs2RURayVp9t7OGEc
tsWZMsWCQoCR2O02V7xwZdSOAsPoIlhxD8He8yHEVSmqqCQZQawBtQUOh8UKinqP
3rXuf/ixaB6dZMi3c3ztbQ9n6eN6NlcChcjfB6wUHI6hbIUQm7RKIyAt7/6Z+8ZO
4M+EWW1h6NsZrbkogF76z6XySS5POh8YEELVLjhJ8j+MtKh3YCdRmkhd+02jIpe4
T903AvB27tlwxREpCNvuDrx8Vo3oUfkHPCdl4NFoCJl0UbClm/3sWMYMNqUgZOV1
JwCUnWU7vBc0pF9slntgW1LVDTiF0l8ArpDrYA3gwJone0IHSFYdI/o3hz7koWjp
LEWD8iVmL0H8UUyPBtGRVxoTYAalR8mKLEQDiZu9N9cUJqigakM4wh4twOWdOhxU
EAWOeduJd/vQ1xQb2Y8/vGeEDDtaXEnSxm3NPo29uZIWGiDzpKLGWKhUitzCmDLd
UFXRBxcgVkZHs2Velik20W9AZsDjv+Fqx0S+PMlqurnlwCkLPB4NkriUjF7AyjUT
OWaaL6Axuc0FIlsN4NY/KyjDKY1k0XtJ20AWPCTMmirnRywN+ptfAMPddSxulWQ0
/v4dM6hvl1v76pcO1psKNOQwqBBooAIXlgrybqEPwcz8vbpq5YimjO+0SPRpyTO2
ybydVuISC15PdfFbtYI9VcTzt/iaszDKJhufCLY4FPXLW7UTACy6Cy8BAxTcDTwh
XPj4U96tApHJ/6XEV7+37DMh+1+F7vpHaiyv3J0FhxgAxTrTwyvJBOUcD3sGThdc
QHczRYvmRBiEstkCXRBQFaGY9m3zhfUFmiOv848t2cYg6QDtjft/91tXShOvl7U7
QTHfroW5TDkgJopITYzbGhd05BgIGmAoHYPvWgloM+1s3yIuCx3FU8D14Ijgsh6q
z5iNBoKmFGcAa4zTvvkNmzWyHcYeoKniSrqIB1jK3nFoYiGPEBhG37YoJwKlbFS4
m3eJvpLqPncYNp12ypprGk2D0Lel9KkBMQOTQjaeUiCc1TsOelm3RxnLA2n5J+E1
wV4Xs/6svhMaM982uwy2qeJMQPPXVdVqYiV94384zKnbEDFs/kbKT7Dy8KppyAFA
IXqa/G+vvRXotOTIiXRKs3v4ZfAzSQWVmaj5Q/x7aTVK88/Oh0wC/panv496wQYo
6Xr2/iY5kWwbVePaFUTzQ/xyFURfAbriXzZlvtwnc7VGwn2cFDKNSOlnJy63q5V1
mFBWnPCbUX8JiGZy33HDrA3rYZHFBS77NISPR66kQXXSfjZl7cXyE9HWbQ182IgK
hbUdgkdqdvzXRIlHlwk4ElH0IHw4SmRn5BdMKI/NpTFef25+ebTgGYZYkDaGbu0K
8VOZUIj3UQ+mY9HIjBZ8Ss6VYMvvOpw+pint6c0zaBDiX2S9tqY/nbzjgQi0fdDF
pJm+JrpAnscXpojq/cywmZIKjPdul5ryCYx5N6UZgKbs+3iVKnBQ70Y51LRV8/4c
cHrA9TqRrn1DdkeVcEeud1iQfQ4MxYuQZ2symvtKk9OHGq8Ehi3eweDGfU6/8GEL
8rMK/uaX1kb9nF/+3e2bOwIqu6Ow7vjCQv3hiHsHt8NJo/xxd5TGLZMaKLwwWOG9
7ljaYc2amCJSb6XoFDgsgV0qEF17CUa6wNUGuBnjnqJViiqzdTH/PMiHaHHUkr5x
wkhBBul3xVPuCa3DHmQKNqc+85xOkWheuA7SWQbLByzMv1YESm13f4DY9dfaiZaL
/PXXHdhx+EhHsgXFsnf9CR40gJzgKpDbkRviUBPBOVgJESb7PmPujSDod3YCULRy
yra3tZ5h5xJhqMEdpdj9RzKBvmBT1qbwiM2YkD3EIc2NDxtPtohvF80dnnHsZ/Q+
A0z80RTBaaWdwsxq8XO9zYGfQwUAN/XqwhKw+9Y9ARLm8DYLwggD2uEILocyhzXr
HM4uApijEdjdtHGNdbJtDulU6B3nK8qdKCHErMzU4cE3HTL1k0xqwebeXunD3ejb
yFm0WrDhAz39Sog22OCB99VTdXjGrlHScpUMQ57N6h1RHNuthNDSWpcuSzWMJ/n1
k/zMdohXaIRdS6Uc25p52KSspDqiK1mloBuotX0mucYLXTX3BAB7C+LV3Y4g1Dr5
eTzna14fb+L2lZjarIb0UTJpR7yeoLT5iJjOeTdb2QEojeBpBRbvMIuSnizjlK+H
Xmn+XiWr90qAZOnXiwPrWQJBwnfTY80eAgJ1084hYNnIjxcf7As2oM66MpJKp/iz
Nspw/SEBbbQiP4BfmH0Lf6Ot8vjJqWXL8BrhnJedxhkkGMOfBsswRt94ZEcBbKu7
mtn3gb2GFOHQaNOnbbDzjJEgyyRLlCfe/MjCSiQftmk6+4cALn1xRdj/h2tiyBS2
GV+BcuRaonw73pamXJuV2YdZaw/3SEhy/K2L/RLDE4jfDDQOt8QyrGjur15DwUXg
g2/x0kIewBzsk7BKZQM2aWZHriEwoUxf5X2iJeIC3DHbCBLf66ULOZwxvp4BdHAp
us834cBp4VtgNLrczANnU/MQyqyo+KqMEW1PAlelQSbOX5XjSLDYdep4epfmeSa+
9IKoQ12Z3ZLP9IuKnoX2iw+I9P94g0+2bsn00VdaMbSvUl2S589k0CkZ6CyKn+EZ
tk+XIhyAzTqS/AbOGeKZmrk93s0YUx6H4liUnanyhBDR4kbr5nesjQzK4qB6Y6rC
4X6WiGXy8+9p4pcMGS1HOEyffR/kIzTn8VVRVkGhkITUJc7Nfq5qatjHRQUV0ARC
jU8HepvVWNGlzXfALvojg/sHl1b2LT6QTGcijo3cFSUJ0TMtAq3eeQQ2OQNXjYVX
mZX3an2p73zFiza/ntGKNx87I0Z+qOcwmSsL/3HvuwznsPyvZVEyzusc1I9vo9n6
kqmpCNXTf7j2ARCy8NOUJiPyiH3696zNTfPyuosy7fCkav4fPs5MZffD/Dsb0Grd
WKwe4f6YLM59P7FewoOrdDFjBcEZDO9zKAEQDQFGYAVdP1XnzKM8QX76TLlkZLl7
FQ9EHvTdU/8MejESvuuntNNmvIPXXpwIvTYaOHJ60Akk7OSZlFQ9Najulb+EhNfq
51YeKxzuD7HBdA9VDLptsc4Y+yV9WZG0yrVww1o4Jrs/9AChdm9GLCnxa+H3cBxS
bDq4oDhcJFtQ0kAy3fBs2oIFrsQKprQ7vPzoMX0mWQwjCCovFfUD1Z9XiltrwiA5
qRUlicfwGw434zwgeoTuWuKOcWoVjQk8vtp1aIYhm3G8wD7IrdjBRvnKas2V0KJ7
TLsMqGhy9Cae0iOFsi9Ro1n7RTKuiFxpGQv0vD3kdg2y7nmMWKktIh9VcutGfIch
lFCFzugl2F4bI8JZlOysufm9HHJmf714Xq2z23nDPl2FcZ9LPP9iiL1JCkXes+yX
NbS52lOs6hRN5QYCqOFq4Jf6buo7DhVTVq3tXYhtanrqvgdc5h2bNiVaYX5m0BnG
phmwhwvR++vD/xUfPC2hHX2eCcQLDnz8+jYLb1bKV2qY/dqlPawhgtrm1N/V7w9j
xdeouOFNVte1Fni7I20uIlGPBP/uWeLfqV0qPagwoEaXZWeYJRev7YbPkDeTGE6p
owRdBvzPEelSulILL4yyVh/NsuIr9Sx6iaHyJFfuK53tNjMC4YtRJIw+fe8+sp1g
p39CXj3l+wKuE/wRoQmaSvsG4LI4OO2CNNrNLeKRzVPq6ECnSJfTA+ltn9oFbCep
YZBUbC4ZEns6JKvJzWMLh8x9+KqDqUX8yGNpwLt7zxLDhfCH/3EJyZRb2Pr/vIiW
Rvch9mZFI1W1WRJ/IS2l5tpqY3qFzWqc0UrEdJly4YeD+vihq4WsExPPTRUvwJJ4
fMpndZ3Uye6w9YQFEQ0+7VNNk7n82HZMB4C1UX5FJVBxeOd6MFXeTgu3UA6jEQU2
CChLr8uT/GRvpuBRoY2ZDyTge25qvr/bYTmcRX2zT0Ch0XezyHnr86hFPNthdI6J
d8HcLOfqPggf2CpD/DTeCtQM0OFbhjEzHsUWuqQUHoz0Yvmy++siOSL2+XLqhyrB
jd7PYMtJTOYc8ZUg2CE0PUZBcw3Udw5Fmdnxv9j1DTtGddUF/6gxQqTZ72ISFOm8
0uEBO54HCJngIC/6MyJi21BnVbuqxj9Bhzc05OQgmHgKdlh9dc2Kt4w+nh3uZbIX
5RHN6gGGO8ZYcGFa7hl/A3H2iz0CALjgtLKT+FrFLT/V0zYvQOTr6IY7pQOw6bSh
+He3r2DKoQVrNZh8GMEIzUKqrSwU5VaeGOedjebhReSqcVGlMsjeuhIcdFNvumn/
8hYm+AcNYqlZanaqtGrWn6P7svSYEKVE23fql55vrVeebxplfbsDpcUpQ55LWtpK
nthepm4DlhBJSuk5leUASpjTcYm9VYYotfdNL3qxiUbxTQUYxp+PZ7wevxlPGzGn
2X+uDSmQkwnA0mb8o+LGEUkfKVoZHmpihYOZDtmGZfKSBXIxzcbvZ+74aUPNyOcP
H/wvkl5CeU2Uh8sh+7+D4aQqCsEzINudIeMbXzR4C6p9aw4LO7c7SmXDdr3QIDQR
IiNj9kTgV10BMEUPnUsJnbfVoq/ZiYoxKm0ssafv9VnGCMe4I664/Zg7HoK3Zf/Y
JRzEhZo20JMwYwvpBD6+9i1nDDvPacca5s9cBU+JysgIikja1yZwVgVVHcztBhoy
V7MRaxwuqhX75m8U5WORZiCdlwkpOkW05EtC18TWX1n4yu0hJEUoCOeqZ30022/U
9nd5GL4zBwjgVDa6S0wQVYkc3FPqPj06BM6Z/5gBwip2HzSMCVS+sSavsQWwX99v
kM3k0DEe8/6EOzvoRMSJY4zdfhZtiZVq1Eii2n69lf+1qVMGz/eL+LU6Q8IU+5Gr
Pw/s+kyEBNClLICKNHwZF7pLQsmNaHE4O5a7DgWdDyDS0oB3koOewaOij6glniax
QLvHmT64DirEsDYEC6uKmp90fRbiounaArgEWBlWTcGPlKP7K/p0WAQLb+KvEAg+
X6nEgtop1RKBcPr+CT/9C8t9oOZTSpEIejrGX3cY/dVRV1TejcZZaX+jSdu4DRtR
Z5ffEWRo/kIeJHLhHz1RDhYsCEqMQjMfLugfEcqU+CmW+ihMnPu1wZubigj2Lamf
W9hcaunhacppHeG82C51ruFvyo/uqL85TyYY10/QNvXkbHO7IeYmfqH9nBO03vbL
n1gS4pAHwRKkBu54cfmaaPSfH5g0XumyJrg8Nv5O/++m3NN8UmnQ9cPVcmq/ZPl8
mZsZv+B487hVRM+pYSuVtKvkDEW/gH/aP9F/hJCb+3oTL8sPYZ/aOT2MFf5vd0+2
tslLHzstJE1dwh5PrFFQcDuudua5EEwjGWesDckE/hCxZbaGWkf//4eUTGNfENFk
CfBKhdcP679y75cOlQBDp5jFoQKoBzRtenkjsleWXyPW79cKNeWVFHIJxNh9OBiA
k/WkV5dylOzrO4tUMR5WRBDnNfh5jDrbtzQU03F1rERNMenEDSDadP38Gr/qKi5x
q5iBm6aijz/vDvO5m+P6b/R0Pqqjyi02/i8eRkbAOsdKY6/CMTLLJAWOjSP/Eq8r
GqgGrkGOxTYHXFzIoWfUB82ycW+c3zOSa7gC010Ww3RLbAg9XhZ4OCeC7kqgzIAd
4NivF8s27kE+0Ciqujldygto87PqLSVCWBpZtavWGzFSTfu4bR6HpXVznfc/dU9f
t4i2kXXyhswYMfyvBhLqQy/OpqXnHnQNyCz8+FBr9FNDKfZDfCim3cDksZkU0/2v
lS7e0JT9ynU9+m4oAKlsqfi+xJEq43fJLA+OlsxFsjyq2KN0Jm8Cw8ryCT4Lk0CV
ue4M7v4XoEtubLVgNNaMohIdXsLProIBtBj7+xXRfuV/BayiQdn7TzIF5kDHOfkz
fuWRlGQc9ETcRATYP6b+17piqVUf3KKdp3DiBt5vWMUpJddLBWZ/qEWJ25DomkSn
+c1SVSGPjcu5o7XLTYTzE6nLv1cx/ZLutJxgdbnGAuX8ubgnbAsBiKSizyU5JlYO
Yt1WYy1bwNhZ1/7+GEI9aLQMTeUF7TXeXVS8LZ1FyUA11f06ibrk0sEXkILLh6/G
uoIqjDTip8V5Oj8DUbfBgQawHEEP8JhH2M365hNSPSAg+kAupywvlm6TJf49s62S
mmo7QB/61L+i2KWA290EKgoxKDhUTt5KVyqq9oE2M8czTRXB2MAQrAUhCjlRE7Yb
4wtHH0Q6tiDmDrQYc/0zuemcpuO17gzZ6GNEGUeb+cyNNnYL5Zz1s/G4208ldmvO
eZU3RVtZyYY3kRUVGeXlRSnb8PccNkQ99SGNVPKjiEvfiHktPXp66/xsZOdoGQOA
rpVklFng0VrIHijVj8mjbrb1uyd1Bjtkb9dCV5jZZtwKoFwHbb1hYrN7ggsK60sf
BD4reoJMUijxb8hSTwYkqt4mFww90bSyJRjcqI6qtYV+7EbpLnMHsJRRjZILh6AL
c9RyYK7+TXXVh5i2mu2KY21tldVJlWl2+I81XEnHHtuLFRgiDgCPDSvEdZv+gehX
HKpNvufR4f+rVmdt6GMcW0Qz+AKcRE2xIrVtKT7vxu8XrX/Mr57XrJ0mw1JPFVTJ
l7rAiuNdXywhN4y32gs9VgFdojmciJKlJt0XV0PIEa34hICenPRqrB0Al4Ay2Oc9
rPQlJBi2BtmHdNeC4fupA7PpBm01t0HtMPPPKNl/+BOu8sOG0RDtyV0J4X2dEVdf
CuPkocY+rYGqkpvdrCxC0ju7BBLf+uhYJGCHcVPW8qLFlLAbync2it40B64hQ3U1
nZScPC7D1KWiVqu8QLABvYLH3GmL2DH4XEEzYFH6gD6+4oLvW+NZoWPNcoYwADG6
URZsDCU+/tN4F22/Xb75aai0fsQouq2OU4Ayq2HfrIJfpcPRpOYy7ZkbCoJg9DTk
0l9LH3tYvIt/4opwL2ZxDSC/F5lJ22Tf15xc5Ec9tmSQiXQO5uTNQaNdspDUfO1O
VxzDmVaTiz6mKpEkXZPbcqvV3Kqan9w/si1CAZuB6KqhpyfcbSuO56pVFHhHoT1Q
ZDg1ZFYJpEtAcHF7KNchv/fl+8gUvaX/VHUnev0MMtpc2GhQKLeeB3CfDCBTB5Lc
UIINftASE7pxVtAeGcQHcaFok9ugRxuIKhVahcATA5tjOfGub2u+tzUmDCJl+fl1
O0enEEzBeZGoBbwEeZ994pMM2HE2Pkh6T/QfIj0ejrhoLo0hfg38EEMYADZaYp65
5aEXx8GBNsD0V5bGocFxxcZpf2XHbGGWhMtydrSVHUuoI1k+JFwW0BY0r4RDENrJ
/FUZzBvIy0ym5wEaKK7Q6RHXvrdrm1nXr7QTPq9uasEoJ4L62KiZldEMh5Bmiyqz
tTbL5t7pjKeKvZeO4ucsWWZMNzcqWiVJJZXATgj0TNpJwRgar8Q7mrUmeLL/2EDx
LBFZ02vfeEfq2z88oAbswtJtB+ltLEK+3/ML4MDkctqiWMpiKapiSVACsnfAQHgT
NcydyOC0aGW6rsOlRND8Sk9BD+QqjQ84gFwP+V6Aijgl/MZE5jBhTavCK557W/Gp
jrAOmLnUsn1+01zCD4EjySgR83l8bWrsYKRuxw9kzo9sWohHVbdAISm2+qfPur+y
zAtKJMeqp8219so6EukJmPENUj5ajTRrq2kkwEGG9LQJTomE+MM4GNc89kSbUXAs
WPoir16R8s27vdCaKticIX1t2z4GEdBpgdn6DQoA6IsUw3S2IRSGgxwmaiW1XLWP
12PT+40PinSmvkldwvlr2014j+AeSlqRI2WNvYv4o57f7dWiQqu1TaWl7k85LJwo
fVSQtLjJJW9xLwNqRzyjIcQHel30gmkayGLZtHhr4R+pswKmF4HnnG//iilYlVva
uX71pCVXBSCruBcet2jx/o9oY55ccaTRqyCHk1IvzmTDLgAKP9RhUmDLiSyWXWm7
IZPek67o0e3G/a82UGxvRYxklka0DXlK69qUmpa+0l8aeczik2nnXVOLJXENA2cu
VdKEFfOPlgKHBr7Of7LX1d3wHvOxHpHEyF2MBZn53gCp2BIh9djMcXw4HYbFiUrM
Lum+EHs7aPlxIwvBZ8ZoT0YTbCzWb8XLF9D3Vz4ycKnJkTuQwcdEavhQ2RYtdgnc
jRZcJSSXR2x9F6gLjhp8ylvBWN6egrpnqS2uQzn0lUAdebtZU7MaFG7s5Kv/uNSi
kQHLGNIGbLxkLagkWcQry+UrQByB1TAg5rrRtjpQIWEwns7fQ3YNDLrjRh9QvdVU
UroY0eKJ0ydq/J50OVOVnMjg68SCQpw7nI72AQI8QoAbOuDjfqNX98CIwcZRv95q
Gilf4NkXAcnmIhJ+D3EFfHeyeSRrTo4sQTGOYwrSZn9abjcv1mMKCmJ5sAGpZrD7
hRAJ4fmmiTV7+LjkX+jN3mPOBX/evEnJuGGyBY90FQ4IfA1BpzcrDjqWvb+S6rT5
D8MbR+lSEd8pvpoTZY4rTUwTMBW0MGLwmVAsKR/MgebIIDGyFFQPhq7bv/mZKGxx
u7vd16EWkTtT8AJ2d8o2UKa4CF/lrqIKJ3IE2YZoLwVAZ3fB9EAYXjet/tXNMhH7
g0i2cObUoYM8jWDo0hFsu6dGSv4quHhgmNMbY99FNp87uW8C+r6pfMV4VLJPTKES
BBiARZxh6Yf8/D9QWNhplluqxwqKFJ/oLCOJrFlXjcQJRdn9p5PxOPNcQhFGEXwu
Vn9/hBB5R02KFNdvGjsMrUjdsIy/0HaXV4NB7xyQLczi7pwqdbx8v6OoiBIedz36
PxXrLMQd+bDBpfDJc4/wVHyMMZnmKrZtnUkKAgqPtJMTTLO3gUCatcWrfolOM1W/
45tizEwbzRRVWPuECQJ+vhQj3ETxO3/trirPADxZJqFMysIx3l9L2QDScRgX5pmV
N/RxJ4EE7CvIMIOOR/Cveeydy6UV8+Di83DPT4LW80MzI68zJYgVnW5OBk6qGrpJ
iclBlkLKFCAhx3MtrLS12s5ZODEo4+Vbba5qcDqrBTb48AACVpHJ48K0Ua+1Umuk
ydp8j+jgPuAfeCkz6uBVHJkWbdc1Fkgz9KYsAKEXpUWXgzjEuSFjqQjJ0kR7mTlh
yTQw0Xe6vZVBox8BCjI7DKx64TLGNbBR8op8fDLesVn3Du2jFW1PUT7brVKiXPrB
Ci87ZWh33diTQw1PGnNCx34JkzysCqUgDpFLBdVcxd73jX3l1gy/naYoiQSHeF4d
UHmSWV3OcBCzFmUa7l6OdwP/3bevzMmeTsnq41vDvG5On7qIhiIVH8SSQmYSae9W
i75/CHyvnwUYoUlM6nFJNUi/pieGXzAcWPwqcxXC3oc8N7QoRPSk69XxTs4IfJOB
roLI4wY4VfCO8fLk0jAE9I1mRo6A3oaO8qXDMvrdMbgEkOkOfmd7oOjR0Q5+V5Rd
H906QHEixdY+tdaGwMoD4I/rVxg94vOseAjwegtE7XFu3fBfN44Ls+jHefBXGELx
jr7VOoMgDRMxl+lqUZ9jI0ErNbYSgJPZ8ldYJbZRRaL8BbI7uOjw59S4ObOH+MQo
2QsAKy+21W5anivyF1LAQ2/qUSBsLB61XnEF/udix8rIHsC9uVf3JYYYY//st+pT
jEQsQD/fyPIMlBtGCB3mFfjepBEw1Q3C8l4kfni7kxwZuDF1a9ZkIXsGJM5gGfVB
yoaTXOyC22QBHNg8oJWOKOdWyNPCyU2XhP0/YOSwOEXkGMXU/2Um6mGvh6DHwj4h
bG9AGyJO1xKsUZmTzkrtjSYRwP6VnKfgwk4KxKxPRKq08UfmcT2WRlkna/4mx6YC
QxEBAhEKpA26Y9RRagobhXGTyP/XpiQFOLqM3pz0Nrfib1Gd2F05VI+jQFzMZ4Cn
T19nK2PrcGnLUDpEYJv4Nd01uPAiGUSnXZLEGvbWijitUblFV2W+C1n4S46mpEYZ
UcxkeIN/4S8ZYS/NowgkZfC401KYLqOptCWya/RzWdk+ZusGn5HcIuyzuv/ppRqq
oKO0Ll3ak77EKnmPqtLkULl5zgQ1egIRC9BEzynRFjSXwGCUVLFy3RlmZulVYak3
Xs1E1vo7rH3/AWVXbm3dwdWNbmP7lH0XmYZ5haP3aJFC0syNHqkJGYZYjyY9cTWJ
mqh6xqdUld678bndAOuqTLtuu6UAuubB++EIS/zeSIohbfCyNBDka3AWJpHavDHN
opwJ7m9XskouDtqT935bgmjH5oTbrXUGCuEvwFRQmukaFiTzV/kpZgpBIidzc0Me
ppocVtZj1lfNmdfC+bqFojozKHwagS2Czm0gP8D9CIqRVezT2KiewT+osc5zvhQL
siOrEsRZkXKEY8T3T7P/ul7tntJKgwZz20h1x7Bhr3PbKU/RSLyZ3vvM7OTayE2g
9Bw/UuNKthrTZbqzM54Cx1DRVqTZRi/+/xq5nySfnkNpWIhDMdhkfseUFn4xZLJ5
7U4Gvb6rLESlf+vFXaKbENmclc0DjSQbzOTs5fS7s00Qq4yhf64IrFNLOHQW107J
RtnOJWHYUjBFIljciHm5Ek5OeAwrjWhEuK12WL4ywfJRXyHmYrdrvYtnaYffBUdL
fFMlQquj6btbnLoKERM6Gz/87jq/2PJGGkVF7dx/KoNxOJO5Z0H9pbthOqNrc3ZX
0qwaHw7wtIzzLreRxhbeqU2MVR/NuMKfDsFNp2+uGQ+60XZVLnWWAp9PARgTO7vr
7TCA94Ju6cVasrhuqV37gmNrqIzapSZbeXC867A8CK2Lc5XqZtCsEsNp2FdwHw/3
qhLXB6xZ2uMqHqYVtdd1bSvrvJ4b13TYyuBJEDqDcFherUeGGVG4iy4mlaX/+a+5
iT1vL95mFkQM5k4zuOZHC/S0GUVNFHIcDt0WBjP6v5iZob61sGLCbpP2UbykeUEz
C/xH4exUuW1DtVjRK0CDKFqzirvNvNb23oMWwNtRdsJTGJ5VU/4j5chOtXab9H1H
vLT+/XgFeru2y/y9cCKJYhOcqsQ6P+eqnIoHBUtQUXMH3gqa5IgXggc3YfW/zlP0
6njVmrzD5dPfMh7sZ6ggutDBWavL4gxzHaqIYlCc+BarN7eDEAijONGVXrEvWFzJ
7HMCj0HKfJgkXcHbfwdQtPWscP5cJDZkkdSwcHIedUwKKr6tpsBnkufUB4kAIpG+
tevhWbjwuLWHoLjO12kcW4nXj/eq+RDHPz0VPrpvVncCdlUh96m1A/mQC4eyg409
g4I2lPmPxTy9guPNJsm9hTxTNJMUpGT/Ak/fhDOnHX5eCql0QLfood5EUoMkTl+o
+8/PLosgPekSmzQiBpLYxFWRY8mzgTbUWH0doo57Eu81GF32UJfmr+Sc0SMrjto0
y0CXkDo8S/vDqHWToiFQf+MNMQ91NyDAWILNR41U+at0gblx0TMY88sUEIJ5a0fv
vxAndSLlCvBrtg2+oHdLLVVzRgUbIcAN1QP2+ddZ08I/O66fTKlRdJI6y2Yc9VBC
cmTGfxJX1zqVlzYKjKCvkI88z2ruf62V6VfSFQ1axjPApIKuZT6FX5z55LdPRScf
La48tWrMA2XkEgPs4k+FuIjKu4dgb82IYDqec58W71PVzleJEdq6sjHAqvaqpyMm
pNJwCQoeF7qSRXIJ5tqX5pmE3Vwcb16HWVB5/MlSe3J79VkhFGkgJfww85bukooj
yXtvUyUwgDwHGApZ7o03Uh/9LWI2OBx82vIlnwpT77h9iKHVYIeoaCTHD5sdopE8
XiqPqvo4q/2tMmzdzcBGcwNE9Y5ePzUXnlVCm1zGE1mkeW/kOm0W7/db0wg7dj5P
Makq6TsX5/4+18W5199jxIrTV/6C7rnpuF+fksdDE5LiTx+JnuVlKPvhLB92qrfq
OR1Jy+4isZiL5seh0P3BQHaMOv4Q0EsS2XQY7CgoaBk2LdYLLULgEXToqSk2yGmt
snbRN8r84/IcTQYYOjpCKhZTj9EXoMEQtXq9TDEnGEGuD10Pjn97JDepL61jfYkD
UfH+slTZysgSV2G3yRrHiuEGxh7OEM0SUEJMAQkQ9J62D/zPZ7I+lZFHHDmBIudH
gB6mC9itJ3WtxghQV+t7y0YEOtJbFBfLMqJIZxCvEUKPyoyBXITaI73BA0fLyQdT
O7cseTd7KLky+9xPp9duadvyy/njieQwevHtQs/IsW4x9EgnURpZW2mKy+syH/iU
HLDWkNglrbXV7yq428Gk2islo3Ou7ZLvLZDvmftlwxsEox/PjG2P578WifpCiRMH
Gpbiqy+C/ITD7GP69bW53ZfAtp1waQwtrYip+InpvOg54Ev/YHcl+4YiWsdFfBeD
YuZ6tRWgxZotvBV+A8MCju+mDAkR7md+5qgVxejCHxPmm1dGMr2iqZ0Ptg8bQSD/
2v0i7S4EHQw7fOx11Xjj/Ge9dwc6W0oscHhDiTOO5qmVeEUJMELPdwDuM80lItEx
cYKqZf1BVtoAsoF8f7Mmd6zu2Ob9tm92s7BTl2zkrec03k7yb3aEYXD8LIkbhzt+
E/c+rIbjWDdqH+nAUBfzH0QHFeaOKJzm412RrcaurANHFj9D7gZga5xl60roPFLh
PYdQt7F7NUs7rIVzO7rwmWalM/NH5rKMZzM/9EXx3H0PLDum1Q+rp8wY5T3686SN
f15qICRvCtmXEA/oxUksbWh8e3zLFH07YseCFeB1Fp6qC02QRDyIho7jnJLIhi4f
S1WkImgsVciR2GaejOaR1NGrswJa5mTuyQND8qQADw+8fsUYx2w/tUA2vMex+qBH
fOevxpnlW4hgymHlbTAXJ5QQS1mrm5PkVZ+grcdYdAay4wXUzYcpsIS2E1LS4Ikm
SQvyb5Wb2DnFK9AtmGGmKJfI13n3Hmk/iuGNh1eoDdiRugvooRtNYCGxe0Sjiqfc
LmGth1EtSI99CeNY03VqPH2B6UeJByWQhUv6ZTqGs7Zh6X7ply0PiJaYZ/QOXzPG
xh1JB05eNodMHPY0fl8Bi0Xs+8F0QBzwiO5H6grWe2ajr0FB68MiknBF6whY7KxG
yOM1mh4wAp0w6Zzh0PdhlyhuSJjJCJPewPEuqp8Ox8ck30COBBtrSPsh7unFHFdj
fXL9GIHJXneczNpaT5dcJzX1cBMCNpHSo0XtzMXkL/mYoPk29Zb8kABlyMb2poxx
b51OOghd9t1nL6xrVxUUCgFxMIsZcd5i19byWakI4gHrPcu0lV0jFZH1H+dz4RnR
QqTAOB5cUVXn1p5YiJl9iSNzjSYRSfTiOZ+nAFkaHXb80BCcLKl7YFw/kOl9KTE/
3CT/U/CBeG4daJR4oMZMwqgB6oIHXOPKC4wko+VZAc5mCZrgeJYgJLWfpHVXJX22
dysO6gAcU8LZsdivKHDu94TZGVIkzEJk0fMseFaQrU6HzCXSyTfnsoj5W4YeQtFT
u7tA/XZC2V467c6mmF/t9w4fwlUv/M5KDrBWIyjoJQHKGbHxY4avkC69e5RW9ZhX
5D18vK5WkJgbRMcZvB7qV2PFoDoNB/VwSRo8mCvObaIERZv31eBx3DfYJFLsyAPP
BMIBsVudIPw7NfBRi86c19T7GN3aSLbNeqo0+5Rx6x6/7PdEHphzDVABaG67QxHU
OYd7Nf2XxPqkQ1CxzIV+msDqPRwYzq18NwIVGxGBYXQbIJSsaGKQV9Zvd0JLiVmA
vuE6t2kXqCll/bzs6L4qKJGqJT0kpG/UGM6YYOlsU5HGvqRv9GGLfFjDX344unNX
O1T7KPEcSsryEqKaCq5N758nkrE56LzkqP02N8bN50228DIrogLPPTF3I5Mr4UE7
2BU9V4/3udrnE42a3DqwF519TkgM02yI9O+ZG0Iaz3XORGpMcY4KlzHOxdbWAop+
ocAtRjbE/mUsu6QNuzfd3wCJSY+zyhY7stqHDsYvgYmIXndTy1kp/IArHQTy2XFP
xuGFXYzQsfHNharUy9Yr+hQyg/ByZePGuCmQzUizjqlX9rihQEJfx+tUsvxdCvag
t2pZT8Sf1Us1D0sHvF1pTyc0eMxe96IT3W03iMguY9C9zeFbk6WrYr/Y9NqI3qHC
j1KaWms/cy+5hxAO2OtGltZ3lvCZPU/SaCdXhP/1eDqXphPk4g927LsKtHK2ctxt
/JVDfL3WEZ0OSxLGEeD7BlaAjZ+zqpALj3X+FjVO2qwmSORboKzkB5liTDf8dg3X
3v6GPI590y+gWvebSTgp3YI2x4SEg9+nJIxvmJVy9tg61dj8sNXX7sWTzIxrcr5/
Lp+7CH8q9eRv0aSpA9+HEtYtURUNldn+G7SgVGJrjPulzGwkHgr+lmK4QG/I46ww
VfRt/Jg4TkQHGSKWFEz04lVI5n7dcQ2WpJbAXMTfDTFwqW3Ks92hmEDqUPmn/9JP
+WuBab+of2CG5QpDTJEBzNnCekhofnd8TCyJJ0VHduwKH9YCo0qnsrtZOHWbKs/K
JPegZBG6YbpNOkQ6zk/rSP/W1LlIVo3HES8wuj5RWbX3bDNFoXox9gE7OcMvDEoT
j+ivl0INI9GMvBfGJcE9r2DgVGegqXKeIDy8GERPOPkISVxhCCAyLDfJE6wBtmvr
dWLwKeLnbALdkJwNq3vofpZhAGZN6NSAtGTF3jYGecwSEh60ai1R4yTJwSt1HYoH
rpks3U5FCDuFaPhdZKTQR2O3f8Vnds7j96VCiS+CEGyqtsL3Vg1+MqzaDS7D9m7Q
k8aZNV4sTlX+M9fW4wEysQPxBxyS3/yjhtce7aidXawYmweMJqvwouO2chVNOwyO
lB2Y3Gx55LTyg5iUQrjIWX7+Ac1+McOfQprtU+Nu2s2zj1ifhf5C0eChvD8be74r
91Y7VkuzF+C6479E1ruIqMF7K1sEfr9txcEHyzA8T7+By+j30cqQDFdkg6W6EKfE
ZR0xuL8Ww31GcyCMUiff8LU3pIPb1mf4v17rji4HwcLQesT08uaRPAGvuMPplU7y
wAOak0ZWiSxC7iJhqIImOumh5J2n2IoqqEwnz8QjEbbFOQvibSVKH35LzeMbe6Jl
clmszMoTOgqP62jO9MjWRY8cVGCBJbvMMFko8RmYT9hh+IIFFa1idQEpwGtqosDL
pid9LzHDzSRYQfw+rQRa9ID/e2PEyF8LXyuYjWPDuJlkLQ+QNAhQFpR0kfXdBmDK
gdkWFF7OC5HBUz1/UlPFH3lEbVUCwGM7+9pj/Kp3Iw2V2INIi5PRbEBDZ0ijVO4k
ZQqhrMj1bneKK27nYW9CRY7gpKIHMgKUCKF/UHUU7NzKsaFTBiltABp4FBEHo55m
zNkiLRB7X3fU1ztfJUs44qIYC8X5LLdBqLX0a9Kf6N3ERKSZ3bHkY5pshMm/nfKu
+uCaaV/6yuI/vzL5tKxwg7rXEs5vbtIz7RhAQcA0scOZXEDu+5Fsxxqgf/++7Ilb
+ddaJ/e8UFMugkgPuGKxqRJ3ZJdTX2NoK0B0rQiHYxDJ5kVbOH3q78ecusrVun6l
GQwAYIT/Z/gBSw0MomlV6VbmPjnHIN8b7kxJAgxZwW69apS7EGEvS1j+7hxyKbqD
w8ztkyAulNc64yaw8RjE+uv/pkNG6TIOlbKqvTUlrv8HiIQieg2BRZEqlEveT6JI
SlV8JMlUfoYBQo9gIbfb5d1Yp8cY3o6Z3DLM9A8kG+AOZSukKzwqFwtQsrb0qitP
1ZImlSFrG2zbnr6oWFs37X5YFcEaIYUk0aZLIViz7prI67wGEblm//6pNVXMWJXS
bl0LwVDVJFu9LBsICQdbMwG1uU40iRcHb5zNdNRXBm/ABbJaVWaTiboQtmgjbRg0
zR9aGQMIjaXQCKa/FM5CQ1wtmVaYZjgv0HmX9Sef4akIz8BHCBcJ8k6FH8kwF0lh
FUG5u3UnDe4HKgMxNn6li2/sPjmM9ibU6DSiWhxxcFJHOEI5uH7DtDq+7b5Pf9LH
TSNKsCvYgozIpTB5MkpN3XFHvR1foCI6gxNqBnNf41jnbflcAACzgcgHk5xKwg3M
A5fyywU5SBB1dcAgd23xLWNxtHRz87rmZkIHbvH0ALgDnXTwXGTf0x9u437hSRfy
cZMVBoiskMpzh5rE2PIVV4bhLrnc3Nho0YZEd9Oy95VjV9luaFwCSsJybqNgdlvQ
laarD6fIttuy68jAgcRPfMnE8Hz1ws7mxLWpk6y5bnL47J/lpGhir0Bi9PLdocCh
e2FMVBSf71iI28/JrjWCHaGyB4i1KcEIvnxjZIKfSz/fHe7StnIA6povWK9AhGgR
iX6j/D1xMFcqE+BIgAEgDrM2/1z/GT+JAss1q6WlFD7HU/nZS0If7LA5rK5lP1hQ
jl7o5GmLJey14InB10aEC/Yp7mPhQXzD4xFOJgPwgieTuWzPs2mQ6IoShgeKDWFH
iDhTWz0X9Oi/UAJHSCvDqu2tDn62Zh2exyGJzdF5dlTyv9sawzeMt0QX+vmo+LoW
/AGYb+JqF87U1eZsqZAbjLzeePV27KK0jCh19oVPzIfcyzlwJMBck4WrotDPnfP9
1pS61fQ4X3pYUgbNHAgPMOMENFZ5tNWezljWp8X2vvmRmf6PBZpOtYso3Jwv0zFk
1w/s3dRNaxrkWGBarR8lCeby6oBosSCJHGNqtPnKmv5QcQ2Em3HdQdocpRCXnHYi
yzhZlamrvgcYCIHP0m2POyovhuA+QcRmofMkmu7j1YkmQJU3FBGJ8X2RoNTXKKBU
RLEWX/AFhtZqeOPiWw/FHgmjzHK3VLSKgQJIunRVvHc4pg/LxJFnpDz8xJw+kbsA
T267zo1hocg8Uo2F6ZdT40xpvwi0nGsfpWITqSQ1ZemGhZNG4xWBJPyweDE2SZHX
YVvZ75DO+bHOxXKLaovS4+v4qZi5dpxaCCQF9F7bnnN6kxmN3kX9tiPWstI18QPI
fJqYxf375dbFK3o78JXv5Zfh++5fNclzgyRvWc8Wxzctbe30XlcFByAu6zLsnwDW
N0ZrRmP9urAaQ05RJ/wwdOhW4j0Hyib5pf85KEB7DvwdXGrpd0W6A644DlgPEoDu
y/ax3Na7b8Fno+0c8qABDJGES0maTMHJBylDIq4/fRDJEwuq/vh3Bg0W79q9aC9v
xFALTdDvYXOFFnISeILyGWV+N+98g/0UEpZIkmKHRiFEVhHpl9vngdhrAnBVqXcE
5DeRVveenJXFS27xsitTO54gNYifFLWJg/So2t7xX+OiXEoNUZSgOn/OzTydH/tK
Zsz47feNPCSWmJrqsNhEbAdT6gg/Ski6m7Wx4m/u3F8Jd66JObkgZo4ElJJHpLmC
I5DKiWhmfpUWLggd+fsIYUTwTv7QLP0sXbNDZVp1+laEMzpCl2OmsX/F4l7V3C0I
2VkUaxN1GuecSQjd2HxaHkRAcmmkRC0pOr3ZvRzCvuviGL3w4szAtrWjIDU5tzYc
VaZOt0jjK7/y3d8DTGvwBs7b6kzi4Gg9Wq8Rg/MroulFoAO09qUJkoqAeIn7lpmt
HPNCGfu4aaQzZshHLwJZlhvkbsIzABiiLyWy7YejbsHPexw08iOjJgImoHKalA6W
ofkpmDRnb9+PZTo3CtNhZ+QRIW5QGitfWL9DmDY8MSH6StpFNi7jBEPJXXPStZP+
6RJPpJ1dWvH2WWIbrG1F4WW6jARsfa9s/f1y00/lboj8/ugqYTXzYgZuQw4niE7B
xNNmdZIsAy6mVxqJAtz0XJpeQ5wgdZtuS8+dG0u/39OLduSMznvV4tyqqntZhz3u
aDq9/izPUM4TIwe5R/LRrkvC+REwBbyVZPjKkFuCSvydaQkBdyArFiU3ARPHYmVV
VjQ9uqRU6x9B2chOEZtAS3SX/u3YBb4NNS93VXLORFtraCTWmjngpMwTV2eQyaJx
bvnFwYXFbhPHk86pYeS1GfFyAXBc3z1K/ZCGRKoep8VytVv7V5O5ySGQSlfA88lv
5xqwhXBd+4oJdSZDAeSJoQL8INDqECFH0XEfdBfs9rRL/iFt/usWwiOe8XlXxVZB
7l7Ypnd2raMA2zvd2o5OxDOcQKrFznLJ7couyYyfdsRWB4igQYq1H7Fz+1I3INiq
2lOfAv+L/6udvYrYM44UChuwWZ4v/RKssPeU86jwyCjDwhOsFcNpekFYuPKVZzCw
S7LP9lDOc3jSeMpY2zhTwIZzERE2SE+S35HpmOHzDgC/1MIqrkbmvvLEA7EKzv6n
Ga4GNW7IR6yiZgHqY6O3iEuE2SrRnuZFSdAsx2yCtIrCxna+w7M8tdHyJo+yHlKl
kgdpAE+zTX/8euEECoU9u+kLyjGN6BexyEJm1mcjYF8IbdyPWbZbuoSjJ9lDGn0g
Z2eMEgPQG12B21dUqYjfc4BZVJqgRUoFTr5Lku+Wb7j1EMGOmxGI+bsO7mU/MBvH
kIbK13ziaLpmLs4lCSu7gE1OiG9v6MBIi6BSorGBuie/yTHo3X/hs4tCGjSJYHQr
WuLGoMDWKB7fL4AeBLKQEbwbqvCVsWQXndUcAWQVqcv/zrUitWKr5MBrIzdnQY5C
fyjOU1NkuIjzuIOnPiMXyTkSSrTg0TCby9ha8kUmzQc5LNy4cEATx4WOXemffw/m
nARVEZlGqem0fg1gLVaGa6U/mI6/RNJ+oiNyyho6Y0fFsMR9uX/ji4l2z7VDvOyt
f/7MW1rdfKnEnLzHL/2Jve+H4VZrA1ipyPX9PWwZJMQTif8E1muPOJIIJZKx51L3
wwXfD5YTmlHeiJhpB1Ow9FnCZnZ1SwdMEi4GvReIWEBBc49cvuW/agDDcL0oIs19
JWdyz2yyZb2Yb47jl2Uhc/Ua/94PNtnLHLMqG3I5RndPP/4DJx3XzoAyp0DflRfk
4V7mcucoYKX+6Yh3cxORG8PgHz88owYOuonkZsM/TpqgiFrwji4VpXgyRSoySZdd
8lzBYiexgNZoGLF/Ca+FWcb5MKv5tDPNMVqFnu40lONRw5AmyAUVH1hjab1Rvqku
bfWwYEMD9gDeNTAe19E72sGOmpucwk1qKhTe6IbpTcAzAtMiDKK+fuwpjvCnBleV
YSyqoQgwXBDsVVKPaWebkiBZkyf7rMet2Eb45oZPD8lLhiZbiOlGwlev+oe7hAAp
Vxs3vxGnZXpYK4YHUqMFdC3F/i6kWKM8WOwARVDpCh4S+3/xFFZ1tAh6vhT9PRQf
TRlz9PDeL/PnmZo9Og9ud+n5kSsdn1KvEGSxI0G8urDBFBwazR37MvKpswySSXXn
ESA55sYa2gm41JPfu7o/m3NT9wm/Z4elr8MjBfBp+JNAM4BRkT8mskrnF7dct1IR
GIgv1wDrozCj/ySqXaA6ED1P0NS7DAAKbpiXn66nKuuOOPYaiBYBImJkt8A5g+hE
J019nkNvEh/MexNWqNJTZuHSbG7yYR8hhfqe1SVb5AcxIOHlUqa3BDsnzIedSMep
jG+ZZqm5dwG4UIlMy6556m9IZ9mRV3IXStOGp665Wi29/cgLDPxeyL51Zg5I9QqF
KtUwn2HlCIRgBw5RWt+Jb3E3JTL13DSTz/9C+UN5HLccxoUQC8zpZs6LyN3tC8KF
T5ZnAvY8DWfNJyRL0S9TCClRrMvqtY8poNUkabAevD7HavOOETPhC2VD+wZNUK3u
nzgV0YFa0KaF9mmb3qpDeuBpTqonAX4Vd+82eeu/w7GUqQzGQY+STAKnc+JWLbu2
5tyiV+S+RNJHJuEnLO4G6H8lS52zcl24lekOBBcAwd3tnJX/1wTER8tdBh1TmdLe
Ui/k7ZS1oU6YoAFJhEis1zvCz1ZmQY7vgekiSNxcv4dUJCZlQh4CIoxCMZy4m6JN
OEWp+igkrw9gg+fxJMrxnw3ZSIsH/mQfNQi7xvoPaoWfF5SphJneO6SNsEiJWGql
B2xu6jDVditZY1MEeWM7Avzh6vbNYQThRK6Yq3lv5oxIxPHfBL2Sac6RuHCOs0w+
7TZJKypp22w19gqYb2Lj9nJEzlkVKmJjL/afQrl9UeXK9ddvXrdCmIrwO6BWSMPe
UQwk27jRYYaMMWV4zhpSXFCMWoT68I5wZsBYCalVUIN3EeQfjdAxp75pZfa7sQaq
PcCrJegAgADp48d2SNjPOfLUbgx9q7DTEkFpPFMiyLl3ZxzSuhkOTUuTNoQqWBVa
1qCEv4I9hlAUCg2U2g8rWpGAKp4n4evQ7Ate3wW76M0Uw7xQBLCa2ck+fDYB/vKa
CKV+OYKHN9hZXP6iuHTNuc9alLl8P1T4OiNDVPAru2x8ts8aoaf09zSfbsKJoWW9
qqg+kVxCz/81t//X8tAJcoVU84K3xIpxTPPGaTNmIjdIS2uL+lAp4/qz44Usr+FO
1C3gI0x5tf4hXgdYhRpJcceM7ZYNJBAE34IkTPQVeqHYs20W1KTtg6GHPaa0ZI87
jIWTy2kCASlMYZzBtxbdjIECIkazdRIqGTT5kR5onqlw0YNnPNdJ5Wy08pl9beao
DA18secfxpXIQO4BobpNJllQ5e2uUMMQVWAWTY6NeAuJKZ4Jyp37SZI6ibuR7zub
f3tMpH2aEGLpex0XwfwJcBMUynLqS0K0Do4PWB2A0ogIFSGuXv4A6NYrBiVEtfMd
1jGKCCc3xmVjuYsjHc1ZEFggE0qgKIaJd1MAIit2O7O8pJkK5+mCHgQvwxlkKW0j
0iQ9i7kAZFVGhSMcHpYOvhbQUlnnPv68sncyZAwYIU+PTg1zaPEw7FfyWValDAiH
98QkPRRmiK0SkV1x8VcRrkr1jdZr/hhiviibqz7QAuX9W4SAYpbrwHa0UoVwk0Ev
ZuAfRLBM2NOPF+Z/+8er6Tzm9xCTI4O9Kly8wOT7arffQfbgXEsea8CpdhoAlED5
bDpBKimWkN8fZXvB37zgX9AimF0Mv9zaaeQXzaGjdExVnMhPOY5j7ginkvh7h2TW
JI2NLjs7ke9lnd2QR5+FuaK13+yUKAqtOpcK6PNi7v7Owm/pMy5Nawc+3YMu+hSt
iuZ2MizKRiQ6d/kmyuIRr38A0VteGsh/cklM8OflXltg41Lc7+h6T/NpqdmigwBF
iI+2JEhfm26AZriZTxpHaYjfo6FW684UfaTsaF5Xal3YIydTx/W3uCRiumMaOWAr
SqME0j1p1co6u6BywBifuZChwWsH4wloH82/oeKy6Vgyi/7qdzL6FKl9TXJQE3tG
Gjx6HT9mBCQtg/aWbgXPKAFWpL+PRI1xIQXwnGWcyRVX6qx/MTVG7MrK+BBQcXSO
IHgiH5Swsb3sb5WQzEe2wB2KeXNsGNlG0uNH50aOBwJg/VyuCrHV+wNquDKPUnSz
OvgrMPsRD6shBUkzqmCho5BxJ8lSp70I/MFNMsAyt8Q4+FQWYngvrJC444oAYc7x
mmJfooDoeOS1G9QI0COHmFTn5aY3Q0QkUU17bumsJuwdwiurFXJzbwBJ/4LuL0d5
fbjq0IeRDfnnHsaN84EW1AuY1R3wlEpPV4ujZHrZESA2yIhbm0aNiIgbD1AiiotH
PCgFXahP29Cg3OjDw0etl/6NH64pQpq+srZo595xCJY/2/3irWe/CAMZt+5HX/gT
5x0ktO/tZ42iu9zTt28EjVOhJHqFWQdk2V/GRDbusBXuD7Aqo1qYC70DqUo07LLF
zP8kv7nrOyR+RpVSTpx+rysCDRZ1OslN3++JJ0DUbY/u9EWkA60e83WfpgJwRANj
FIhXFFHt4ENlUWYWxpInoiLprLWilaGujGsClP0v3L0IsSQQ3e+ywGwV4deKyAHk
5bE+/dbE3lnfAJNWoEUer4CUl0C7OoeYpphPp3qIkO5CcuGbBTejBk4dxaPoZw1R
DdXO7z3080E3nN7A58f5/lSRL6SkpxnWduytrRQ4rf69aHEAk2Wtfu9cLu57POwk
uS8+VevH6ebUBRYVdJ+MsaSC0KzBdHRT0g5xDhtkG0JL9r7bECCTR+d9CAIiI4/E
IQei/VGIvGHu5iXQGU5hXarx40tRiX+xQ09fslrqSr0wV0hyc8MGoWsJFsMDSGnW
W4OvPRRCmCCFA+NyJRKVOGFkkl7sRx3UEFTgP+e5jgU+Lf4Wb/1TMagib7QXDgyk
plRe9dHduEO9K/mwXKJ2i42Rq0liBL0lupWpQCF8TegunGFgDjQ4jAPNQ1O5a2sh
Ymwc1A89inb0tXBiImhbXEdEhLlJao355CrI69XHbbSsNeRR+kh23ht4o9h6bqU3
mRS786bIDyIh0ZRoFAJHACyBoQgMXj7c1I6MwgRJpQQzQIsLWLWVccePOHhvGP7t
fF46byfKpIRfwxX/R5UtbLiJ60NdUWdoPwSp8JpihKnlQRnNvKglbRNaLFcCCv6z
9uXUIsKwi+oZdmha/NPrI1VGffmj40vIRY8H7Mu5dzWpcovi74tm43R9fYrvV0+Q
3RkZv0HWLPueHz5kq24OTTVFT5er7F/RM+Ns83ryygWNSrTPzA05AjEO7IW5kzoa
2Z0y5LUA7U9605bAyCQ3UOmT//dJMw1ls8hLsAymj8G2zYsUpz1W/5EHbvS8YvSg
irpwu0LsS2zlVEUrZYj2m7OHhf7I1rhMiogVStgWLq/emI3IYIwm0O9MR3/sx/2r
EQWZIk4OuJRFvsHG/Ypcv7KxqpWoccLWlJgAxR/Pbw37JGTTkJDH91+BdaOlJ/Y4
JzZ5LyO7FHevjggxZmL6fJbb+Pw7kcKccmtPCLu3dgjGz3zk5nbj1uJZAM01DovG
NdmSpNJiWpRWbcJCSpoof7HOAW9m6H1NhZrAmsWpIBDCO2G1ffmb1qu2j9u6pIWa
AFY5869k2qudHhrsEf5fIcpwn2dM4ng6eWH1FTOpFBauR3+ctpa8FYrcJjNo7wqZ
GAjRQlNiEk/eaN8ojGd21tlvFstpTVT/KZ/+iWN3vXCYfC5NVHN4UwFTsorbn9Ui
5nGiH1mGwnv0AXSgjdLN6xGEak9294lenzhu0ncsjYhB/PxsO1XI2TEUftNCvUIV
uG/R1ogtWWsj8cnkhdYRuMn+JdIGzhcxUpZjJaPTctvMSZZtwA6MpZFqb9m6AD6f
+SYeEAofSyxaMCLwj89+quROM8Z9RoilFmWaCh3agR9SktDGNdynzDAa1osZv9pe
KlupURj6UG5oeAY1LMBMOkdFtA5lFzRom/2xafXwb37h/sCtT244qMp4Py8Dl17m
KQSR2wlvZIBXpdyJtiFg3V7jwZWfRBCJIi2VQ5mC0ymxx2w9CVE54op6lJIFYbyy
7vrhKouiwMxL1xys3fE58ytepR6ri9FBp5gBRbqAcZywiELcre9BEsFmmDubVQSA
f0IdUnTObMqEh7z6I+WilRR25TYR+j2Q0bHAOC7Of0gVuLXfN7nqn5Hg9Ze+ECpX
pRZ8ZtIKjS6i7/Z50Xx7QIxBe0MsJ9/6JN5wbrpe49q/dwlFnBmHWDtd+KOd5pHc
1ntB/BBu/97PYsp88n/l8hHabBuCEkbgHaNJqTK4CfkebTB7xnK+e9vki6LgqNlz
jMiXy8LZjiuV7uNKXNISomZ7FeVsQyqtKfxYYb9zIfNR9HMyRUIXiJsIko7O3IkF
XXYeuQgIU1Fc+O7/cZh+KFFaSpgWEAayiuAdKWbq1/9Dh2Gth9mBz48E4tZDAs+h
w1iikqqQbb/tBA7f4oE+wBM/1W2CwVmL1B/5CHHluFOOgQpQ5o92ncOXEk0PtSiv
Jzcew3OYB4tsJ/ckUNqLfNFG8A2r7PM+ujgFXrzVdGIMrCT6izgUHOm+KYS9n/Mt
6GC9Uoww+udVON5Ns4V4nWw5n+0QfajVMWPrpTLeFIi7v08qamubDbuW8tdMFlr3
SEhsHVkw261oQGTuZlZXrUvkzKbmEFxHCrSfJacwGic77s/pqz2VqrXPe85lczmZ
Aw7qcJVXKgVt2aG+3Qoh36hluTK6UVTcbARW9hVSTiMMUFCmVtMSqjA767JP44PV
r5k5kRJwkx6kZEGPxXggz60gEwqWo39hn3yvuEIAoeWbVv9dCkrJEPb3QrSfgp4D
Limlwb3czGghN+f6qpPDmnmKgxSGfVW3sT0TZxwBhB5XYfBk7y9TthgVfmMdj8V7
wjQncvvgLiJkq33IZWKm290QXwHGLSjXXTPQgp2ciGvzsURQO79rJSnzNedd3GHR
0dfb/T0yv5aK8B79YfXZHB303ZLfoqx8Pbfy3uhgJrUnPnBj6S0EqexEKnx+iwhJ
802RfLzuUm3dbThZc8/ERP8e9710ushBP219+5UTtI5lbkH0SrPndXbKZ2TQb5DF
r3w23THEHPR8YDxz8MxBRYjdUlRgkM2sFbcU6McbSoiiVYgwzVWaPO449xhym0Ua
eIOPJ7ItcSH6f7pmMeyRHtVyVpzYQyDuJxJApGGEkQ9uG7eMbDlrKDIFKvcxWrRM
teZkMc5t8YjKlT28fksFeOdE9lERFS5MBvkz2G9xy43GFQrCyARG9h1ppbVOG1qA
tYoeJeq567S4L8By5sdyno+VT0b1Vq344wDuFKGrdu1fv4XaS2VKruzwkoIeMhLF
QtPvrw90HCix5juykadpXDh+Zg5p3fMjzo56SaDonD3KqiKy/XZUpxVubE3HXaZp
xmSpae57KmldavsUZju/BC0+5TDM/lnjFKZxcWSM74O7Jur6EpPMTjLiXfrdYKVp
0IHabdun1+eIscX9+J8uu+dzC8/U44OD9qay8gU7xKpvlSGceP7g+vSmYxV2LCW3
KykjWeoTIR3o63NvDFCggXN+Vo01wBz7/x378qzc6miwTmI1Z3E0Ks2n6opUHLwh
nqsgL9qbX8+vqAas6HSxGJzgKo9AjON28j9oRDM6TA/vBEHpTfs8YpPv3RBmV8gO
ulvQBYuKaovTbBoOS66p3r0lSMgKOy4wwgV6LkaYLWz/6S8UKDioQGduZLg0ZPIq
+w7SenH3QswH9y3CXM7mtbRxTRb823UmBfijqGtMlznwN7N5tuKhW0ZmKsItflE6
0d4khH98xHrNrGq/FIsJgF70bXER7hKMyZ2hpDhXi+zPL50zSM8qnht9KuWjRqZY
7xJDz3rO2QYd1UtYOoMf/W0ikF5pRRRxnwQ5IJuoy8AaeZh5k7ilPtn6B8/CNA2P
fFgUM2EcMiRsR4H8BVENSORTUEOnDAC9CMMuBI67+WZTEW3OpNJs8X1WHkIAb/Uy
2pND84h0tNdDUIVUpG6rcA4GtYRFeyCaW5UH5Pa0vRxtdO1ucrvdMva+Rhp0bvEo
YXPKAONp0QfgFpRCLkaSCSUdxWtRaD6iYUyL1Mwfzxb3fDhLgMtFDsCbfMKgEjvD
aM2WIqi1KaPaq75GxI/Ue8oc6rRbQznal2dh09S6OBPR9BKVDK9rwW2yMI6zL4F8
UGsZGhLz/pTd6RHPYty3xnJDrQHbOpt1ELYFFbaxI+f/q4e6X5oxdk3b4YBTKUE6
HEB9183uAqZZYcvrMlj0mtx0wBdB9rk5tJKqn7FcNOEL9nhJNJDUW3Jyn3FhrYlg
iKqGVNNrB6kAOq6RSb3sbl85DU4HTtZuZxSk6rBd27RQBj/T6otlbkcCG1JnGaO0
eMB6QfQ8XMWIyyJXXyITmsKFd7GMZK2ilWP1aUm80nWsZ6uzieWW6eSoVOmI8vnc
ZtWHMBa/3eKOS4KaVEhDYksHLtVbx4HMeqfBpAmnm5K79Yfze21LFol27Yev/fPy
h1c8d3P4+guioout7+eLUdvtwIqtloWdsPF8c++6nyiBMQMSzETBVLa+UrdBEB5F
I8lHbeAADOUZ63blEislH+T5Jg21VHWqp8MV47BU7PRY6qnCZRDOwOF+lHG7rGyp
MstqMeigQNeWyOcr3E7lYrUyLrAfgYJshdIyKapxNcjZt8NJXNkbLbzzlHTOmvx3
sjS3KGqrG0xBvno73n6IGG1oEimF4lFWN/gtz4sLqeuIOvRC2+NCyRo1hWY9s3yZ
uDivycVuHXZIgVSm/bxOYKRDAtrd7SUZrf5aLSz/LeZjDzD7pkLW4Ddj9z6T6GF9
ypZ/7wdk3P/77bxd7tmgblofMa2aIX3FCKM9VXmlVjbs/VGzz4MQzqyvRtmJTX5a
Y9YSvpN3IdwUkPmUgpdr5hKhBRXKXhyg+n9rPjHsr75DLHRh1/+TLiZobgCT6N62
qaZlb6fnjJMA1YH3aWPqs4cCo25nqcIDcq8uFTzfRcaxjHF+ev3JKKOW97XPotTz
OAbpfG8pWKolw5strmWLL33uiVn39D+w7OtzOM64iLN9ayGhemmvo8sS7gm4nyg2
wMzyegSRmKtUAnDoABrtz4EHg25jOnm5eDRL5k0/3hfa5+qH4RILFJtNcidUx297
Wi5/mdnzUOsWzzYY15syAmBFepNIsj+30gtwxODEuTooR+l8NsK9ZbmGKngfz204
lkpHvU1nZThp5+bkUeleMHDbdDRzXlFRN9LDAL9Uy3geDfYkDrMu9ankysyeh17B
lXRkjYy36iK1C5sFfKhuC6aqw6GWYeUPCg5q1n4TFKnsbZQDbR+17vG7JpQV2vZx
4PYTw//iVeYXOg5i310fOY9IFI3bqfJfO8ADaxbUdNqm9qUZNlnZYfAGlXaYBWo1
6W6BWlTPgr6L5tujXFJiHUZpgMMWXAgEJC4l7CdiOdwbZnYLoNpzVbqn9fGqVoEo
K2hI3iM1sw/pAIsp8ZhOu8aSnnXqPMYU1Xd9Cfa4Ek2wVbEFEQ+QaA9WRk8aH3CP
sfjt0Ew/pfkE0qEvq7qTl/5LR+t6ly2QJGuPlINfdkaSfaR6eBdtBM6rjcmL7naU
YSLTCxQ5jgrK1i/9gpetgnEKD6YVbR9lMWTv/AAhXmSu0HRwQLHLZn29iQApe9vN
mum8bGJz0EBW6S8QyUUSDdl0/Bk2tiVBmiu8Q9oVqbBlO/amdh2nZTVlXCaFaIC5
iZ4Q9X46Q1fyoBdQDAl4TxKF4Y3IsBtUM/vExNN8nayNJSAx4rSipfv8pv/qqTfY
i/uL8NU6zt9Jmp9dJYQ15XhuX5dVJaHE3BEujQJfz8wWCp+/Hfao08FuQj87Miiz
XOiBj7RO1RytyZZGY3eVPVFkkzHI9Y10W6ADb2EGkak6ifSZW6cG8kizO89V9Hbp
4ddd7VR8hJxmFgy7qVQqPGjuTT4M+2TJVCECbsBWZqg4Vw8UAGDMsBBlOIZctXvt
UI0lvCmCTE9i7uXtxULb1qB2UEpUCyCHb6G3we+OhhNMGM2Y0zGX+w8WiVd5r0Yr
C3DeaSsvOBtXR6OCuZMT4FYMFmcTo1gQjt/yr7u6eVJKhrY8jLNkNH58sA/K7QLQ
Ykmylul3728Vgp3c8j72tb0ytXhu5zL0ux65lA8I1MZskr6DhPJ2ruNWWAeJtera
fK4+jqQmExw7hCzseHF/l1wRn++BKeieudFMndudjS7LqIbbozYzdmUx6aNxW8qm
nVtDTiG88srmm9qknxBGyev797uUIVY9tUfPKzE5uUUJe76CgP+3Xkg1/sWWxBxK
NOsUYFjekjEwXdTKhaPm1NiLA2JEo7uvFk2n325qJl57nKCprq5caQVWkqgIt8J2
izXoUkK9vK4QYPf4jjk2+WRGugGPW15MCEdjHs4dfyQ+8AzSfmqLuB18MSlvkiGW
PJy79JlvxHNrc84mNz++Psz+wR8O4I3HsOXp+JlUaRQmEgeAK2NqrpjTM6QZLxgN
iQf6Sn6dzZvYnT02IBIKO9UeCQLq2H8WmQ5B9srRVixWyAEhbKnB5/LgCFu+a1L2
xoKVIA86KWFK17/2KIskd0kqJ4JhbQu5hW/ZPo0Pbrc5D863uhSZ5QZur2hhE6Qk
+JX8Z/Eu3vPRxv3biNGEsb1vWcbjlG7tyRdSTbZNM6JG/nonhgIZzqqBsABoRhAM
/hWmzMw6toobthuguRbRkB4nY9qAMAV290D0MFrjGxBm2XqzWEN0cWsi+KSRXI1K
fzb6kkrALWTa8gXjL34Amgik0rknmOwAEDloOyji1fq5XnOLzRkGlHUvZ9tJrktX
2F3mOZUVZ4fY1Cw+KuJFJrfBUT+wa8tuSchBhKkAu3MxuiDBLzRZr9LDSumrg0Fn
6UaZJxO/tpD/4hl9Tu4FGkHg8Lk/EC2v8HlFpqG+uwv9Cf/g8U0ni4pwRhf9Kd3O
ToDo3EAdrZBy7+I4hA4EWab6XZLKKKUrKag9YWDmbH+s72MI+XF1V4SRR2Pqo8DD
tgZwGaypKJXmFTdHrHF/naYUhONXp3dsxNk5LDrCltNWKBnc4ivPS3TKdZVyko2u
vzbjP9XERB74vUTMUISFExmE7VaxETFMrziR1rJDApYq6R16o7nIEFY5e8RudUtc
HlJNi4s1geZCE4po1ehWIjcLSZLh2viE2B3oeUlOI5PwGNSICdUhuar80hPGbET3
5zUHHGiFxzT2En3s9LhVvzXziJ4+3Q2zxippDNN10h5q/ICOz0i8J2FHI1wVf79n
VlHYAuInuSJ+IvYmgwrjwf4woNt6EPhiwGBvnj2sREhtCM6lt4OwvZtu7qF+whhN
OFyC7b/6mx4lMOS61nBGbXXfIipumfECTE8bE06osLlQCk5Qach5Bei4IYS7HKGU
7GHZ7oKjqrM6dxwHatlcyxz2vXx7M/OZwPPautHO3WiFR0gS8hjqmANGxVX+O3f1
nH3MAFXdxMP8KLqVkOERxFflStWc/txyYzNqRzBokmBDTz7IBRpLg3AIDOFI+Yt5
aoSGhExB0GAQzbKMh0PhnVEBjW2jpAjpqjtrOMZF1rs+otaFmGscGr6t0Hkxq4bW
laFs/0rMdIMVGLMd8gq6shhAaV5XAL0koaP1oevhvbpgVmVNx3SG8Fbqpfv4iI6g
VnvUx9c68rcNIi5k+fz8xPtUYxPrDe1JZ6CQc/euKLkswhio9W7YsWBUIwWGg+S4
/5hhBQyg8KCfwBaxCBAaB7tsOyHisMCsoEtCIH9PXQvWyerdXMBWVBQIAZ+syULJ
0TpEgo+acPPIMoHILRuSFKDBM0t/vpi44xj74Oz3X8D/HZRS0JTKnPbIaFwjk38W
cfwLSTLcN6poMrEq59LT8ZgvEMdp1p71ETDd2pKhuLDDdjjuU3jMRSh/pOqnr9S9
L/BrbgChlSORGXoJnoVZt2QBFSbsbWJ3GuFByEt8Jov5PQlpL0jQ7sefwQSx6qFX
v0Z7iGMIg3yXafk0uG0lV7hGa5cPXjujlNbCWUmfUfAVTBx6JqesHmWE+9p9QhB3
atv0ivLHmM1g4dCoN5bqPAv6WYcdZa55/sLDCZV+ss1VE0alot4j+7nOKyacKMNB
P1IhIl75yGho4itWQUNu4M47V5TYn0sDF/e7h2x/E919nimN7k509n5ISv7cVcjv
YUk7zpRYmHcJo1RLzo155ea1NluMw28q07dZuHIUubQqvedy0yA7RyuFx4gXzMLr
YYNwG9T3g3M4gijk04dtWqaaxaSl4HHYapE/SO1ZvcKz7+dzturHxpr02M38Tc3K
47zIYFFOj3gEQvOpuItg1+t43aGZ89qEGAStXFBHsIxV9h6dk8iLskMC9jpMkcQk
pIexagpdeT/kuWEYmb1aRcAjDgwk5syzpluRjSi8YYCohraDmioIvxKTTvC0lzd6
oWsNdeAArlauRfRtyc4x/QIsVnlx6Of5QYa/APDxJ3JyiXzF07DRe8RIQTWYwNxZ
QQr15d+puUO4x9O3dNlOh+fAzZAZBgVVp5ZzbxzwULS/oGZ/s1gwZuZhQJ6LMuO8
tkmVOkqsNr1Dt6sJgbJRPtZGCrOFAs0NoTpOg5kEG8v2z/EPb6aEj65OE9c5UQ4w
KLGECOrZZLAMbNwlv3mgOfS3DDWNy2Sw3IZl07b8bLQyjJHLZZhpdhGPbEUa0Dkx
Rq0CtO9WUyj6Vc4Pzy+2YefTVVt59sHivAKr+/2ZABvEExaASI3uHP7Y41Qn4j54
H2LBZ7FVVfvjggrSA3gYnrmMZj5CegiV7zDlOjSy/mAz/XvRSz0Gj9YdeIvkdogO
Mh4VXRelhwGn3SE3hqu4ulu+tmu7BOq1mxEJiQXw5QD4oLrV/8JhRYXwSFI3iZRg
2rMH+W9v/aZ5PIHOkNfnJlVdKNe+18+yVIpJ112MrqURXIRA2+frs1rM4wPGchYV
Bw38JFPsuVQfosCP0OW/+e9szXMbgn/fTzZMnAXBEel8mUy7vXu1bHwaa5EiT9EM
h9Ah7O6teCFAGO6G6BPmUuEiBhu27mbbHmxMyYqHm7Z9I+g5bm6ewXcgTb17yH/j
2LHvNH8IyPGAFNnvKLmVj+dY/orvFzKib/zX/NGqeMEJmCJ3QHxrI+eUafT40aKu
QxQFxiiRa0r+qhdkMOHxEAWYG9KUVNoDrcpAP4Q63BCZCo/rIMmgiokzFF4Iy6R+
U95z4gzkqE15t7GyLguaimis7dwcrFw+nUY+G2PTEIzrQrhI0YJgbCVb6er5DYpu
v4GFeEoAtTN5w4Wbv0b4G0heaDbhHkjK/WlVgvTinq+ldmnYJHotA+w9iJ2X8Vvk
+CtNwW1on23Chs6TpwUG3+kQLkemfzGipylWxd8vr3r4gQngZv/lX3Jj8MAoY3sE
PIrk3kDkaQVBlVc7ZddnYt9LUD81C0TmX++ZMWJW2BJ/HDgrfPaBax8HZ8cAD36X
O4DyBc0qgIloIF6FMdnuKDv/ckji6UaRZESHco9/fkRYKmTBkxKavaXwVeW/gMNk
IqjUFSMJgzIIBaXSzCYM2ZXcZJlOchhJ6lZ67H8pV8YAbqOCe2eeRYXRfH5X113M
QSGHgrb9/26kjbxmzwC+ensaBsKF+qUWA7ZL+zcGw6p/Jr+tgGJzwQFAPaH34o6E
VriRZAlmcIVEAIrtx5CPWqCQVNut3LKOrXz82RGH+0lyvjh/bu/2cqTk6C4ocRMJ
nRIkkzAmMIgVVG6dlchLL7M0Y7st3nUBEHK5Oe013e7vkDx/kowTfRlz7CCPekmM
8vJg6OUcPYrTX5M0h6RhT1KCpBkdVzKHrRyaetVZZJZaVHAK6PYuGI/jEa5fTZSm
y+/nkJr2XiPWV40Zt7yTbS6qx0r9CxqVp5FwQtX+m+JHNmWaSEcM5FLg6VuOMRdo
9Q8z4muTNdw+nJH6wYdykRBf+40qIvesK+d/TI1uuGPdzgFucGvmb4LXztvoeZOw
pTUGb6cjnCe2hsa18MpL5mn1CzA9YigWWuu6Mm0SFNDveZQ+y38wpKprryU4EC4R
Ha6wwcLUNliJwiEkIrXv2xTT8+NHktnWr7SVnI5U9ISM/B54F2eo68zga7/WSfLR
uOU802k+Hr60St1mjUOPWWdFLvOaBmVLTebbbqjfnSgG2bDXWRTUS9qAOLaQvgtM
iaFoTIUTdQjUQtsHPr5iqRFyNh4RXKHFum3bu+6YeCnPCiPUZaL2GxJVdE/aLDuz
vCH3byIbGUHU3xA1Nos38VBVTJA65U533qZT8rKJSqCCrODePgyR4t2lsaoi81yS
DFZHruhVYBbC9slEA0jV2PBCA3WdUPfmXXdLkDgmhIqcFwoggPa3LcJHO6JuWnp5
DPVt313JdM3E8vYeuyGyukzX4CeIX5faVXQnDj1+35B4sCiU/D7CG6zsE0+qBKCo
+CyntCXiwB0Yqe0sW08S/r6Bck8nq/Lct/Dg+u17gB8nScMhljeqOkma5AzW7w2N
5vq3Sg1smL0S+EmErZppGAvYFiPm0SWn6cU1NAVo5dfzqpClzzURkkR60I4S4X5i
6WiImqwTWK8qeSCJFh+YAJWmApWGhDAtBERRJ24UgKB/yqBPrQk0B35KF+5vtKTh
R3Rs6HXZZtte3mc+v+UH0wF5DxKZzGVwZwSCXxBGdKX2rA+5dBgJTOnxgXjCyGcR
2EwN3CDwg2hZJg2skVzmU0nAfP4lf/q9dEVwFHFR6DemT4UzCXn33hWDBgHQtjxe
8OyNSSFNVQu56FCYtCoNlOK24Z4XmF0jUl8DgVeTcpPZuUXY56XtfEUnQwJpqmx3
kHpiM3mx/74blj0thss3abzTBeai8tryTR2Ut45W8oek/uq38isoQILWqkguqeUl
oTOwvQMU2lhQkW7iCPDEuhp/2jhWMIcSQ/cNEzTtt2M8CfAe2L2hs/Llqm2H88B6
FZ4D4yjqBHBjufXjliAxXqC/66vQ5f0iAofMh98xASTtBLBWcprKA8/mg6/aHd5l
3cMY92VrzbdDKoUp6AJMNuLc275uYrcbL9kXzjPNtcjc/UtdbZxSeJxT2SGwH6qr
E11UZEohxEt0+ipEFIWmlK5TUSRulcAKebLr2kD1Sb2PIzfjRikQSsStzIjZZEB3
qAtianZNN9iMOknwAMeOEB0Zjurm/1ZSA8FnsNxitIz+sKd8vjBgfb2ZOQuTNmbj
ooTpwhYbtOBjvP6QTl6TSI5TyRtunvzxH7GxAjYTTsVALGGZ7hkQ/r4lKrOXdVW0
SaW6yiLwGVHisUFxinyPcCABkrStxY2K5mNQcbvTdiY5R3Sp/XTAwtr11ZEh8Bmn
m67/NOkeA2pSlCzuBXVXKDo1/ldnD00GY8zWuyXHRTMm14YfC62h+K1SkgBy0ExQ
ZSz0SaFZXjvU2xIiuqldxqOpcTNmJDQPOrJW/DYUlwCbrrLK4q9U5OTYcPJASy2j
gOpf2bt7ngY4Fo1o2FkyHaEnQDm/npNM6CXDpN6kov4lSilc0VP5Ghal0vF3yxZk
iyUPOxJBijusgYbKScLV42zNNUKNWp9DCeNjlLWni6A0uPpaJRWZiXJEbEdYDcGv
zRYn8PvJ01XynK6QHmntJK2AuL4wJZ0OsJRs9b4kLWH97yfTBc+Q1tZ7DrB+IHu5
0YFCRwFf9Vwp55RxVgMLoSix16Yv+dlaNLoNOxOYuTic5QiEL+jVY77c93E/l0Em
crcXCyMbJNmA4G87QmsN5Z+QnuYUDSwY/ekAGlOyxeP7sKwZ3gVGlavYero6Px39
qu2kXP5H5K9yZIhrcyYhLkriflxT2biyQvcgbg58xh2gXafQX+EI4CFGKbM3ECUN
lR7o3pFQ3dwaZgMZK/9+botKJVxfTpL1jcY54bJbiasIWLEaFGODQ/fo9FZDDsgW
GdqjqlKRHRm6T3m/yHUKU2mhkLAYIOypWJcsRCMi5HVbg8cVSFXPP6qp1aDByRAu
KlhQ8zkozneIlaAswnfbIgWUFczezTbvKdqrWRpe3w7ecD7hdYj/B9+3j2g05jHa
XbCzMPqfuE3od+QHRCplnaxYJjr5EjKq/eNno8yFc6CwO9iJ6YZGtWiop58jliBf
KrCJ/NFdhjseEdaT0OlpnGJDYe0JdsIKDQBLioyGSCp1Z9+tx9XXeXAjR2u8ZJ46
ZsHnaOhMV40aJu8J4IJzFJRQD83maXOwBaGb55s0bFGK/BnmyaeG3fGk/95TtX+X
MPrEduY360Pc4Nc/z/d0EhypCS8LLkedtjSplKj1ZE4KsBO3VvHuGanVMFYE0Gv3
dw7ZukI56WipKznGiSHhnowXMyhrlZ4ucMcS/me4d1VMRy0Ymau3TB+5jAkQaSe1
PXV2TCWnwgcdmmqxRQnEOkuS0rzUG+z967x8U5oNQbQbN+B6qmqxtTdoKG6LvyQo
EpPt9f2DhgEKJ4AbUUjvh2oRDgFcAbSZDbgvOPQKQ1Mbthifgk9G7LBpkxbTMqFz
XWy37D8PaWAzbk32N8Kh79JGOCNMwCn/R3tymPBSswxjB6AaferqmKPQ61UwHBIN
/KVzbScmzjR+iHq2jgvuvwK4FRUKOM57LmXXk1DzkQ3m4mwDRgIWY8D6fazWMnTX
FZ9dIUffuy/cDPwwicwvr/9AKoNEtIBnUrK9sjftL7ZZZRoDZoNU00QviIRNBRzL
7b1apCHJQC/2jf5iL0I5jHe5Hq4TnK3Em2FHS+E4WImcjqH9AmU9NE7qQzr2cBqk
6f98hmiTgBxLy7iCwKPV4LuPutU5oR/5UzGtui/tpokgOj1Ya1j2I9BuHzXgJuC/
oUrkB78wX3//TH2dX6xPKEgsnNtjuvtNR9WsEEnn4RqWcOpVz4ZPpodeicOlZBZE
QIzjMcn/4l6hKfAbmT4CxEQIyIKOM5Yk57maVYsy0fLjnieifCcPHVbQ3Xt2cfSt
quLxzSYSGQfChoRHoUYM+0P72r0OzGRKWBzKbUjnmeQJCt3mDVbIRnIE9bgRs+Sw
WyWz4l9ItD0U8Fp4aXi2Tjwu5LyMAxLwIoTpMN66dJWtDdwfSCJM1b4HckYj79Oq
BYWLVSnthhPRW3tsxTWgl/Ve8iy23lbe3LUXdmqXWFOJxxafu8gracAzyxuqQ6ir
Xe30urjUq7orPuqciB4icgiLg9hBCccYYVne5XKUDH1t6Z0jihfIpvfy1Oy+YZQE
R8DENJuFryAs9TJxWU/bS86RLfMzDKDGwKhx6+8rFQXgT7rW59UAL2UXaz3h0Ule
bFGPK/FgFdy29e8Mz0xqZiU2BZocEsM2fs4eukHH0Il9eV6IS0OBXCZACh+vxnTK
2DSroo8bgEpN0JjKnYYwYSIJC1q4eFkOLSqBIs9uzphTtzyCrkPf61HW1H67EYb/
3WJlhZsXnIzERghqZEEexwTqcq27CtliNuo/HiCPVClEc7fxBQawGBdCzKxrEkR8
aGNA9iPBK1GeHWzGxOgZ5+Q3R3wc8pvTsCRc7s2dDJEm2z9K8IZaNppg58fW3+Dk
osmjJxSqchjiTQ1JtrftlZYX8ekGq7x/60puA3vg732Fbk/7KvQRQZhDyRyk7CqF
18aXrMA0KhavY/FZOVXpg7Dvwica9KrTSTut0Bioa1JXc3YpF+02exmViutMdyq7
7byOALhljnNpE0bDGxzOHpLihWPOPdD1i75wrlN8lldiki/OTzPWQYQs/vR7o+US
p4tHHXyK5TCmRZ8bcEkrvHqNyfwnHX9JYYWKTNZCTC7xlNSF2v5qnZZLsd4sYl71
CYqcYoJl9GJ8Z4QsNoTTbjblPCiVHLzWuQH1Kk76Z0hjQDTce/qnPZf1KAiwp/2N
thI1FzI5o66WzI4g8lnfJwpm7jNksqnCUduRrS7IgUKqI+sR0znALitsNujGpXja
P555tUeyO1muOoUoGHaTw/9Pv/PSvfw7Gvi4c/htm7oMtXp9VJsrqApqEFRdEsVF
M81MkzuVq5qZlUv5zQB+NrzGyxqD87r49FCiFvtMXYEimnA2aKTPXflrI5cJrbYw
hf0/M7KSi4x1YzDaiOeVWTq5qG7fVONL6Wg4swGPtHRCIpMWR06osKFoAzXzRAL1
mhZf+VupguMGHnDwPuDvL5wrtCHj/YoruLILVutWqhuIg/wsyt1sEXSh0aoMTnOh
HDLknxWKHLSGTwNrW3W6Tp7ONEJ8dnigzfSmrAaup7wWDbJmlS/KO28gxhJgEaqu
VigqYGSAcFiL4alsJnPWGoXiZ1SV+MGmPXUZqgtRgIpcZ2tyXKsvioYz9UQ7bquw
kqmD3SXP5odGopzio/EMR6sl7o2Hpb7UkPc3emwhbvWaZspWWh8AyQXEckjcRjkl
184r0G1d/3nRxyag2m4BOIuvzdQ2Jc5TK5Rwa27Nn0D+ARJq0PCOW2mhKoyddJg7
4xoSfYgBHsBXVuA46XN81oalMAOTfmXkHjZQIdkZ2WNCijLnzsXRimq7PilyofhD
J9hM31vziUvCORz4SusswvQnrcr7pBvmFgRCUxfCQrJmVTQz1vMsVX9+zc43n+uN
VsYNYL3vwi8cUy0xEzIYX8CvlJSzwtKD9q0Mrlc6wmNOZdxWYBCTLUwVND6A6ta4
6HWMG+dgnqbmVxefc5sQNYm8yvSMCh1yyfOwGifzKXZUltgFPqaN9dTZsda20MK0
rVH8erwEljsYJ6vQQiyqUVjBif1bkev/sdZmjb2dAh719Nc3+dlpoa2vSj4BI4yv
EF4rG0lqvkLT5f3K6uY7avnfrHs8bSG/e1DodECNvH/99Fj/3CQOwPLwPoq2xYOJ
4KUH8WXkjIjTMd1EQaUUjl/rjMH0RfQ/q45Obf45pwW7my8JI3r5CZbDSefi7bcl
9faYpKAW5toXK9b+9YtPvNGgMPB25Zn8/2xbsT+705l6SCdEPg7JeaXa5rWNht3O
UgzqJP5ksmS6glLskX9V9hnUro8SlaeKMxedkoMiX4vVGj69vjl5jebj50e9Ropz
hbB4Hm4JUjO2FRwGIyxevLThYndvcTDOzmF/wnR3Rx2CeOresAtq49ONXmgVXBPb
0tqM2vqYCa2TLQwOs48XTPV6DPWfmB6xyHHC9C7aeTiIQ+FOR4ZxYqRjPVqul6/N
zjXzu9NToi54bEKyMXpGAbW4iZVDwsgGQ8eqiANI+RexojxETo4uOVecN4A/Jgb/
OPzG0imVWfq9/GZki+awHGAOV4CZYuwTPxfFUrnfLVJRgCoiQzleccEMoYUDWeNv
5Lxt90ZFzBzHitrodnIkSQuEayUbBpAAXklvw8ZzE5jyfm9p5+LYplkSWfiAjOJ6
+70aGsXi7Cl7hbn+0Nv4TZl7MhjThp0ocNQjXzXujrqmArNEAtmVcKvVwXd8HwsO
pEkYlQNdCqBG96X8P4JMlIgcMd6S3wewr2KdYQpkxUhx0ztnkGBlWcgvljgh1kh5
1qOh6K0PVVKZ1CHzinEpGqkpzlvj/JA0y3u/Dej/i2UjMWlq7JSMDvI0b3DwdFts
sxUxwu9vAjGaYdwiMzdnEHz8HX1FZu2nLihq4GY0L958nEQ97ZuYQIZLg/ZvCHJI
oAJbw1r5z6A0xMHnT4/Ilhf7bQggxFU2+XCu5zrWkcUfUv0lK9MhVdQMQjSM5TLk
FpNkhUeKj6tKVEQKWu7zeLI++6F6rgnUU8Pgsm9hYZKb2xrB/ZY9vtdjrELDzqRm
IuYyfockXT0lUTINSvokUWKrwsXDRZz9MlmP3hBI2T+j9Ga/GFcKCH/O6Z+HuwQi
zVoZgrmdgc++0CXHDMOnKT9a2o01J1HRc9GP0pasMWxpT3igcOKnpTvx0Gm0dtCa
hSYEXAMIK4po+hgU+JE8xBZ/QzIuL7oaanfSKiLPQVROu59xPiWcvndRWO7SKB4K
Yn6s2WTvt3TIWfHxMPgqgwhyaWq1LxC/rDl97S+AzlMdn/bk+28+CwxGTbiR+Qi5
GBRiX0EvJAbk7Aw7/Am2K9Tok5PLBt9q87ZOElZ43s6r0AZs+u4AxDKqsyCQ0FJV
roKFL3cZRrenvYk6KGY2APSvEp/JCtwggrctKO54YP7NpDoT3XVNLqCTVTXlr1wG
tg1PmXol887N0T2tJB7Ju8Drrdn9ooLH/bJHX1CbO2surm3ZOzNX+N6WhpKjCQB/
LhQYCo1pIM1mCOFjoCnvI9SIercEgQNP0Axy7J4zxZW96XuH3YqRto8aAJZyPKNc
UkQvogUvt5sDx3at89hxZs0hIzqexkxe9FxVSYH/3WgJB1Q7rPIpmvceWDWd8T3H
FGALkZzH7gxD4k9r4JLtsGxrmBXbLjMO1KHVuLDJx2B63yAA2+TbYqxC/CUs9Ltt
z93oD82RB8T2vURUPmFu/QBhiEdQhXqwM2wqX9xZWcrt+C1iCf3/JQ6uTg4yhjeF
lS11r4RJgCHaUDMm3YrxYDY/eDpYfSy7PxItvB++Dp+KWGQ1PS3CN8C1GC8Wyg53
ay78ttuJzb9bNXvIOe+qX2GHxPccHyVmCgNnnSE0qsEYRYGp/R4o6KATDY89/V/R
drEiDxgnQj/rWLADeO9fqSVCrXZ5fUOlSOfqOyuYr6ShM3zTH7xIwcYSk5N5xnGi
t1VCj+f5WMv6QkDJi+X4aMTAvaMoOgI1EOnsuGSfHz21RDjaaCpbOo+RkgWIXCXS
9ZGKa0+iwTDo2ndU9EZIUgzeQw2rimFMorfJ8CUafzjYqxZ5G5ILLLCM6cbN3fzC
ZF8snYnkbylAAQNwkKQ0e9sZlwIcKhCzFszeLJBoL8H5c9UCzDCpKfUE8H+8suqm
/yYTUOgcRI3qUKlzOz+IQ0YodPV+t8v/YxyCrIL8sSvFu3lsSOGSH+Qj5P6huPgC
zXjKdLwTiKZHJzCpadBXDa5QblHfjo0Cbarbx478J9SpFueWBU6j5QkzSaMAOsNo
m3gDtU0AdtIx2yaWggduI632imMUE8H/DfSnZHiFFwfpdkF3MR/hTp5hB0hxmdD/
0jRx84j7174VPVmRpz6lttMmylFxrhOP+ZoP0jbw6PfkhKAyp5U5vHBqGBCFwujB
GUsiSKaFlQk+t2XDZK3mkhv0xeXL795eG+hznwHF3/0ES5pbhmU6Pu3nFouvzeEl
KyQiJ4xMLu3ch/pxq0+F89EL0UfxZKxlCLwHBY9UGG2DE3zFUnlc5T8vCFDB5J0h
fMn7cTJGjnQCb/H8U4IaGipuQS3Be1yrgGk//JjCO8hUT0KsXYHLEV1NGtqHLIc9
Q5LIiiWlRFaYTunokSgiFoRi7OzcZa4RwH4F5XFTW0TcTNUfYgeWEunnGlH6fXmP
9uXGPbr9ruIGjJd21M3E82SLV8lOgBs6AHwllUl8HkpD5SBj4rqv9Y48SrpIKFso
9EfQOipXlgqDOi7mNOmY5Lo2Y0PBSy04/qY55ZwZU+xL0fy34xWk+9YXZUr52+kz
8my8TbuRHNATM5BWYevtm6+y29xYSmqSE3FJkjFkUz2mpwWHohlS4ljT+ziFWazh
kx3YZh+jFmmDcpIMy7UkzKMWJx6Ujyjjxejaqmi2/LxQqsqC6IuHEL1z1v3H33T4
sERqrGj+8kUTb3mWG68cZYPGS6VQDONn0cxPTwoE/fmXMbIroYe+ph/P33/CqT3l
iQFLClg43XB7syByNlRMOmrE+dAo7D0aGA0CPToEorDw82vmpCAxMmXXfDOcvYmV
UO5TIpvtT58KYlENNStItapJ0qCHTGnUsYQWeDnwBMUPxmE0pz7SbVdN1ash4wDx
VZ9yr7B/yWQHsXbHxwhm6Yt+DHnBOlc1GgYV3X+mjMIewR19FewCu/Ehkb7nv0xX
DZ08G2TuWspuA8EVysrCg8MkMnPcO5D75BJh/x2bkgxjV7+oRGZa9VQSsXYKSfQH
RpOGpsighPxznlskVk7pHhFWW4tzMkwB4N+UT2nLU7Y8hhJqnEjY84zleFRQJFAF
RzwXAJzRmJ6MOKpXdT4lEUmP+dRpz4IBaiiy20CbUp8QoduhDEcCQFzbd56triBr
MJktqryPtsVMdPqst1NB9MpFFqaYbciXCXYPObiY4dw2pDGUHWVtZBAHUDiVgrjS
1b1mE6ZE3CIqAOSIr2TjwHdO4ViSqVs7N9JOWhBRyVFoXkK9cG9qk4t764H2y+zv
9jmq8qwkNQJ+XTxxNn47MYHz67Clhcz/aVWu68HZdPZ+7mD0hlSxBaRT3uCTYzcJ
RutHwPtNMmFgistrJGXra/sAYWr/6hpqt3MdmC0yLA5JRUEo72RA0INw+/Dy1OAM
AAbjoMJYMx+EvSVWFQroZkx7OUJmsgZkC4Aztc4d9Kr4ijwRDqEFRGPZRVu298Rf
yrRG2Owfn6+jmBWhs0qujRu+pJqYaB0zyWdMWfUxnPA87/2Y9wpC9sGmt/jsPR/C
UD2tiBtBq5Yzaav5Wc6Y4PxijGMrWYKrUy0BKmPq3stk2hl/CRPRAEnbXTRpGCBF
WT1Ie+EWTWygnJc46CccS5eviySCKH/F+WM/UMtrgeDUB6jJcg/Kwbgt/CBMogoa
XyQvgLy56/ZBX4eg9pUuh8NzwKyY412/jo6OkJd7nVYrDlqIy9hKfwvHluIxwYJd
zfd67gosZTwr15sX7ZQdnBMk6YZ+cKob9Ljbr3rwj2FMrw+9+sfDbzIc/mYg3L6v
FinRQQbZD0L6IF9itP/Z1MAmIDbJz3oY0WhdKcL+CCT+RVtIJBCiDsPAxFTg0cS3
TZSaxit+fZODkAcJ91ZwrPKF32s5laN8B+vJCYD1Od9q5bEouGARcpi7tyyjkvkW
8yigLjoTnYICBHqLdCOcfF9BaFq4e6t8UAWu26pyl5GEiVvg304YJvEcH03BcWfQ
cO8BdUZnzIbxjjBsGdkMx/HHZ3tdxoa9iVMmBGcDgSeci5LeuoMp33IZm7vCrE+/
VXvOREnj63s4+0Gig+oCifCFCTtcf0ku5QfvndQI2axhuTouI46x3az9uMLF0Za8
DjnEFUleHJRfWon14Bx3w4XjXZmqyD2VFcTF4/OiySwSapdTNULdP8RWKhkc1u97
kOXLIIez2sHZAUpu83p1mks0C5G8dXQ45lmcdvKFj3FEn38/IPGeGoTBCOQpjKRo
grx0jmq9LBWLLdNO/+G5YzOUsdIYOivbDlZGpP0oi+gxMVvnFnqF1W5PJfGZq1GV
m/iW8TqC3Dxdp3qpnqC+IVC+7AZRhMuaVbwfqv3wQ1PRyYUO3iGD7axdzbCM3Tfv
SWyOr3SnwkG2e9tuBHlPU0wRqyLOb5hZ3h0thzD5dLAzt0TmJy3FAnNJQRHdlouA
9dHC4tSk3CX/T5MhV1gCnW0LP/PEoXpX4E8F893Dbi5qS2U3f/x+6NQvb3hfJXpP
Gd4vE1JvimMStHVdkqiqv8WNK6vDDlZ4y0a4iWPeTpIAsB+gkW0FWm6fp2bCQFg6
KatsAFUqfKlrv+Tt5ni86G5q2NufhlPhnrCpkugeBrj0lh92Eb2ZDJrGOnJzCwUz
odXeLZJabUGriNNi8BOQGT5feOVyykRYsnhoVo0zqL2qQRExCa+OZYRrjmpF746d
qQVDZY0wAvj/q8I3Pttd6RvP+647YhjCXdR8Y3RwwNEBVsP/qwGdWU753C/Vafop
FrdPeIOhXE/V5FwX1GZIQ39lFWnZeZHYIIKZ+PP/vNPTbqLUwkoCWhw7Rdentu2L
CmiDSAaGFktzaTrZwPSlXkemHrdoF21mpJAn1o5UuOl+D2zQ8HylmuHAftjOhPzL
zFwMPW+EjWAdu76imhD2FybA/33771yBuT0p2mHn1G7Utm3VJ3GLm/rhOxYMOuak
XMAjZT0ahTlvvzj9zEvPykNUERLeeYlD71BAk9EXAOAhi2YKgtji6dN3UHtP5Fg0
relKET2X9lLvjYrOsk2b1Ajd2f+HYFZn+u0mhyKRDaDV4pnJepARVhedRuf1pCMZ
rexXce3qbm/TJAG86wlQp0hgMmx2ZOo7Jy+2GaQoq+Yq0qz4uh1kPlODDU5oS/3s
2cU2pB+7Ks0Z7EHOXTcIOykQcmtGo/c2QEVGZvwUuI4u04Iy6JZ6u+caRPGQe/Wl
Q6zgno9jZ/SROjXj+PPCzWsajd7tD0UOzmWduhI4fiWHJR6dNhqR+7DOm3OWOpwl
GQaD+e+NkzUC1gP6OnXucBSDUG/2AB3V0A8iznfXHvEc1meCyFjkKkPZx7IJRbiw
pi9/tj7kTQP2vQ8zSelrZgB1gU1MtC5TerH/recKkakkKXuerKWEY/DqGhG+/E5+
Vfm+L1q0cjpQEyD1q2CL2E5bn/mDPhr0AzxB1Mjis5w+plouCdTMmEtKf44DIknz
7JVwf91G2pMQVr2Zpe5yI4p4oEqNkIyejXkNBCPHCZk2CP/MfYWb2x7Rlq65sLfY
gy2zw+JwjU4s1M32xwHRRrDPuk1+zrOvQd6KrPZ9KFcp6hRnF9fAA2em2XLooHQR
cZC+ZWHUaYzAt9g9WJXBaGDrDRMTe6C3hnO7WZbCmHGZ1V1qJyFunrpWTaBvvi68
XmD0UQz7ZTQDWq8X2a4zLzetqwlVzBUQUNm+xnXTwFwWh80iIq/s2us8IpinixAO
2YEXdWtzoPMHTnX7mjGtJ2ipRU8Rm/TIUqN1vHTsmjlpDhM1+FtECsHChUozUQpZ
/naxtjj3uIvfs+4TUfDy9M7RFL+W6Ut/p+42C0NjadEKiZ39bu4BSL7ooTeKWLJz
Eqtl2sKvYwxFf+HKw2/xM3bl8PFd/DwapHY2D0gSklLfnF7MNXhKicMxa9GFevDj
x1ByoI/WaJSQ4hy3Y9sQOteUIex6qzcJkaBX3YWzBhwvmD3qjiIZ4pCW80xPdmZv
ootTx1hMHPBF37sy98BoNzFWclYhr4AGrHMgHnMYH17jpu7qbwJp7/jgG5Z/dQ2y
Wy9kG4chXlRuN6WVi54xq2ONwUC3dPcenl2HLyL8Y7rxDe0t98fgGrU6R3bYHcag
0XUSbmAa1iuMRdRIFkf1OWPMapFkl8P8HMISMzDi/JjrLy9ZMUfVIpHrPi/AMUbu
Vq4sfkblsnoQKPsNqMGaBt28YW/RLrfcI05TxJ5TblBbRLHkTOkDPwc/b20exU5G
RPpVNZufMcxmVUDs73NQdaEOt5y4qB2NPTPCaUDZEYfZwIw1UCuDejl3NNlVxr71
qk0YXfDqYPOfgXmZPK4bp/Bdou283dOpVU34y1EsH4+iQB2Z8mndIeXKRtPjLtvD
O2rgCRI8Y5nQ2U37vBVZio6wZI5+0vIkF8VUdem+c2Cyu1CJAQ0CsIQGT0afy8mQ
6tAAx4HYDhY+koH1Sr5MRBSimC3l4Fyjx5PJCJY3G218r5q9Q5sd51Hzj9hhjL0/
FiKQtL9d7GKQwRnptylpPbwJxVAekUqnFRRTwtOvpYcXqug2jOLNjnY7m6mAnhK1
3lkExR3MazpOZ4V6dCB2khPVMbEfWRetTvlJaMZ7zWDY4bsZGb7SRp7vfY9fiPm/
C6VYySN3F0pBMA+u/yv68yUJl99EvCzcDRBGPFosYBp7r7WO6fHup0+g8au2Xi6H
FBzdYSCU7vfZRNcW9pd0K5PC7xf2IMBXr/qo0xjKuJjEhPd6jQoLZriDRHNtvKPH
2YTFXkbh3bhARuxwhnZgUQFclYBkIBxlHoT2hqpUzu6GZSzNPN9cNmoqqCc2bJWV
D1Ss/iICFOyckDIfAfctg6g47rwd8KFUTH1mvgyV5derKintRmkRWyE7RbikxS+8
Z7/XqfDXHe5vqkR9zP8qjo+T7LRsEprDfica70AdW6/k0mztUx/5ga3mOVf+1Qk0
G9ieiFMt8Is74CMklVQQAMwgqLUYXc97eVp4eiq7HdMd1tAU909oCUleBhbL+7s4
erQwHvF9XKbl58qES/WDQy6cQb+ZlcbG71nJArVtARiXtqJlzgVUZSrbimmO5QLa
9Pk+3rH4LH3fQX+DkgzhDawzqt++xS2WRN9uIvXOyZd+TH1rv3xZ4d9OoF52hhnC
OBPYZkWSn5k3k64cYu9AAkB06evpzF8FkrE30twSLEYoGDlvNv6FEpZAioVJpZDF
yqUxCUKG05yQg5Vm+e+gK6RlwleDvWyTE69dBfZt9TsjCbz7B0DKyxavNsbkAwkH
e7LHOXxQjcUUEsLuuDtZR3PPt38hFUmpYO/DeAQ6BgK9Y1KRSqKtE0T5tt2Vhnuk
a4O0ZT/WY3v+iocRFPiHfWeniAZqgAZiuxUl91kZQ5ta7JtnGijeRV4ZJT0ZJ+fC
UoIheLmJtYqmBft+r9a33Dpa6gwhNfyWAK3pEq8c7phFXpuvwJk46MnwluFxC00p
p71BpnyneoP7GzSzV7ie472X6EqjHMdWvgCsJaYuh56bQBEK4+DsVz0kOSyUAmWE
OHyfXXoaCqWL5lHvIzPxN2aR5xS5E0nN6rtxKOrcB7uqzKMpOsg0j/+/o+ffXxqo
Jbf/Pza6ZxpzYPkjb4HCzReDumahNdmIxMQ2zKNpMr+NkyV48pkvv/GewuYG7I5h
rsP2bE1ecRphuK2A9oixEEbZRcTK5wnEbOTln+bZUHtUACkNQh92R0AIO0ylVOfE
U5R5xR9cOKhSC8xhOdYldxLx9mlPN9BZiw8vdH16hQC0peU+/3yGaWbApm3rbFdd
XcRio2ZCUxrENbyWjQR5f/ogpGukKEkOSrB3Jy6uBUD3gpf3AfsyoNEKIF9cAZeq
aviNxlrnlG6OSeWhEoi6EVMWyIZ3soqavXoiec/gGdLfgQY0cVp0aanGond+WnpZ
yczZy/oWc5zumgB3vp7Ij8XjARSHVjL6cwG2fAw+4FHjUtqmHaB6BgnKMwH2xuBa
0G1uXL3/SXZYmwsqiJuUF4eUPzxpykHk6e/XlWe56+ab5ekN0E67+KnWhZZl/yBx
HrNQS6OVkx8XrGGNWyfaicy/SYsfjWa8l4T6iKQEMfu2Q0sWQ2pt5zR4+loMBBQ+
MSNOyqhcDJjfqIvX9IflnbeSK4qFOYdfDb1OntBIEmySAy0rz6OecLI/OR/HiDMF
Nflqe7IBDjvssqHwa19dFdJ6fUbd8OnRPwmznUtip04/pHEmpJS1zhJYOon5BuBx
+R6XjH8ZEDdhmCg7PmJzziF9qE8DqzUypw3W5Gdv5k/UVJbZ0V+Trzx6vPOEqg1z
VOGtqYwbPTd3kiRgom7B5LIc3xuzn/gi2G8sldwZNapVO3I/7PSMHk7g3hdhPc9X
N1qBoRHbL7O3hVU/HnE/FjmTfIyUEmBAQUhdtEV+/FcWUstmXfxLoxPLhDtsZT1Q
uDQSnLCwcAD49RFEwgXi5fi82QwUcMB9OFErx2DxBn90jO1s3pw56l1UodfZT5DZ
D/B5uSa0zVBMLbMr6fxmE++6MnNZ0GRbSKHrlOgCCIUnU0oLno7HBs2jZ0pRYkp5
T1uN0jKlKCJk7iHkOVXqeRs8QkG46XouDcP1/41ksq/S9hmnaQxz63kWWNO1Rnej
MnQhqpUFfjHerw6NTCL6rz/FDWP6dHRLfZ2XIpXybGQKbCZd207stbRZhLv54mZp
JxxMR/1VVCgRgcLvIhHnSJvJGR3xcJ4g0QR6TfRZYQMKZS35y20aQY5uCHLXSOTm
ZlZpYryiQxHJOmxt0nwCKSPX2QEROPkmeYbGw92Ld7Wf1QE+kaXbmiVLfcUJxyEd
Hvk+l4Z4pKwQ1swccibxePQjInXI8XzkrOKFo2dxY07jU0XJhZanUfM0RLHLmmaQ
HLSr2Qk/kXV9je3JuilOnMy16Kz2N4Nn+fMHmnsxhDQVWGcgSa7aTCsxyFIXS/fw
zrOpvEtLfuVrAGfuonCusJemMvJLRgT46coELPwUvQv01yxnHqv3bFMh04GYy0LO
jWoq/IW2EOerm+ACgrKgQjoxQVMg0V0GAAk8NV/XHQvi5+qwWIflsVOIPbo9GMNd
HHWqVAR6tuGV4OZv2wB4ECJvW17+ieMmc43mNIDyZNsqy6Ce2PNHp3laIQP548TJ
2Db7GQZkt808ynwk0a4UZhKINiAaZ62ydWP6HhTbsW5TNIWTupQM3A72m4jyARow
8+CFWcpDIqqRduteT32/JRlxRyLBAyO38V2PfTeXleLp7sTi//tHnyqG8gw4xIQj
SRclgYyjr+969mwK9tgV7FODJMWy6Zh+UDTnMqlbgyeYtXD7NGpIL4YNPOn60qK5
Hp/Qjtpjr7mszdhonv/8O71qgNvFH7WA9PG3V8aCaR5/CoArb92F0flqzlc/Fs8y
TX1pFn2ZpqyWZqy16FSPHl6A4sbmIfdRjGgpie1Q/Z5JnottcJUuNpe984fg+K1F
XcgR/Ezs/gFV7BTeQf/wijEMbyp6TTZOUmMK96C61hmMCvKffvPx63r5gIS9GjD4
rH7ozr6a/MEAc9+sLNdGk90Nloj9wWX3v6hVJMTRCUnSpIZsPQfp8AYNV+dtwiDF
dd4g5io0HYuM7X/0bQHKujKY/tMijJpXy4fxxtTFdVqsw8OynMpQrWrxv5HhMAfy
b0FF8uig0fNDFV/sdJHwk1DOXIxAE53/eTtgp4/4INeZf3kHHLoSsLZP4SGlN/rO
VfNzJnKdzLGG93rhiaqe9d5dn9wACphGxBAVFpF5iD1dEYHdCjylkKjcusfdeP+t
h/O9OCy9fQ+Gll0mDgy8rlYEROaFPaGbiYkQ2rL8xEuBcyrJpQslPfE5t08u0T1g
/L7Qgvbaj2FKBukS/JfUw4WC7zfzmPSzV4Zpxdn7m84NvqEUS94jja4B2fQq8xVA
SS2EEf+2b+4qdRDX8umGezihtu9I9vnbvblve6+we5HaADeiDhydfUmgNaEPNY/Y
WWEoeS/9Dbc+G4CcpumXiRVOLyQLJluVrWXCUF8V3B95ENiHMWqCgEvmpVSKuRE/
5jKaajP7wkv6m+Ckum5Vh31Fk4JEvZtaHzmCC+R41BK+CHjm7bqczBsYOWLW7wP9
qfuNJUB9zNWry82IW6kIDmae/6N6fDNJ74HbaeIt2fdsGwUnvTWpQ4ehacK7oRfa
kcHQompMjQbqTQN+Au0ap7gq2EFqhUEgtB48eRT82a6RUOYf571jvnV7NRwleIC4
i+IDKAsW4kpYJLvjNLODV/mktS5C03VePcOC9CTydwFJAWQu7GRqgLi4N9eegSKw
p2koG2caE/w3KXBpe2HH+7PUCMxnWfP0mjvUds2lUI/a1t45/2b1+0+XxhNv5oOX
CCxU+GORebYMCo9wcY+f0i0QSl1BW/9R1uT2PUl0wFW5+YMMsWnhl2r471hYgTrB
sBE9u2KA0SyjkKTfkc7s/khtpaP4GJbYiaHW7iUCF0SLg/QoerbwVgwZvI1y/XOw
7OVg1pl6x4NmML89txI6lbKWMxoqMoSng/x5eG4V/pqr4Mz2hRP7SV3foJjqq0Pr
EIVCltrdzWmGslWNW0GMKKappC9hoSXGEqZ/Rlg8ZHQySunIRw2y+2v8SHti4Eao
1fcNXBVW+x9figZrJg49YW2j0Cv71Zjos5ui9LiCHfdfmYBtkAuBjVllYDUQ7EWI
DEsqYxsRPEerbmyB6rECj/mtRQ4GiyCb1Qk96iGU+FO0N2UyqQFF9AW/y4OeKGSZ
lwjsMAH9MrxnUYpu7Xu/9rVp4HG2aP/dQBclYaBopLxcTjJpJeRV6JbcsZClb5mj
8Tj0lMFmc+mEu5ji/DNfPP6u6IOT2GwVVJNEQ4JkvPjDXMivfZPCTu6Hen1gq+Sl
83WTzA0/2HmIUKD89he2Jn3AlSBy1vajelF9RSYY5EvsZW3MxDnneiRrEppBKSTL
qBxAoVHSco3Z0mPV9Oh4AQzm2lTrd+was+//dn/g4ct1I2aeBGkKp2kFFGlqec41
7f+abICaCsKK2RmtULBGziHj1bX4xOrcK1x0ncbftpmOTL6dYBo94ZCOxpfPq4RJ
Y162t7FaIFQ8mC2mTj5tWfUA0glsSGRntRZS33FdSO476B7ywJnGjrZvUFRRHAm9
ycQ8XHLyMPUeNk9mgUUNfkU82V/lokq4SXmU6bD5/5UrzkbbUIRjZjcyPwnrfKkt
pyZY/sbIyoxpBtLYdCeJWHzTrgtSyYReIAVl2TgXHjqMyPvbnPPdApj1WB9pj30M
fBn6fl3g4ObystewDg5LHf/oAWgWLBCGCSbfAbh7RhYMLyxq3nKgLOBj8B04WoOz
m9jujgZjx4n6kRzE38XNDxcQ4OLUDvn4jLD+RYnkMFus/qfCZfgq0qqsMBC6cxNq
xCa1je96nWEhNtDE7vcWhJwA1/DH9G2yx4PyDW/w5FKjYUG+IZhyXKzkEn5BWDPb
NSUxurvka8EBfoHTtTHtR8GW/2ljhdauo+4s1F1mqaexL9vDmVxq7X+t5EdQU7Jr
hgbNDhTDXVnFc7quq8whdQb0+zYazJg7fc9OH/k5xeDKjNMFEeXVXb7oCEkwk35q
rYqrwUxwDX4pKF8Mj6TLRXdTkDM4Ma34f2Z1gnwLQKR5u88p/eDFOoXGKnRhhYCj
JLTv1g75V6IKEJYQRByPwqjExRiX0yJMWpNQN2smBZnSDnNOrpo1XVxwDYmhxueS
CyTc0K6WTpGP+7lZmz/YZlpiaUNDJcUweV7hQQ3QeC5CEA+jEo1OCHeH9s0bVabn
XISIY5iF0x9KrsMPIw9I7mX9bEcJDE2Itiqlj7mF2pMNSHpvl4vHwSkhL+bBKumf
Uu5sS12ymEGqbgem2PkXZWa4qulJjArpSdvcafexRH0zZ1+Hm7qMVIy9CkHV84qt
gRcvCEPYjegucatgh3dGYMHjiFuplebU5RStShU+aADgRHYFpBLvBEjhpD4nGJeJ
VzAytNpGtu4H5C0OCCSZl9q1zIKrcuo/t6eT2Yd4heooNnf6YekHeLbCaLFVB879
TvGc38mTy0OXzR+5b00c5Myjis7tq432Aa651n2CSa7ojBlDhiQE3J4WmwLd9gNC
FxKHRxHMjj82IVwurJckP5ZIYEOslGEIkq/EGA5IxwT4gWhIhEC16Tb2QekbDBEv
ZDnHersTm+B4q43lHGIuDq2FR2HmbNhZG8V3q7jt8ghjgfTvme0yQw6ne0YDGzJn
uUJ4/eIm2czuFoIhR9fpZGiFgXq0kEmnSIdhMF+vFMg2qKwlXEAhgbEZyq7pJvh/
yEj49R1T0gndrFm+jSGxEN4mBkPD3Mr2+f39XK6KIVO2MMyBp4XuUnj9PXuIx2lm
gbYshgQZbZMpktlTNq8wSjH5jnsi0QGhmR6vO5vbH4Sli7qVZF4qf+974NZJpU0e
ddRRZ8sBBcVUX3JcKO5BRPniUGjyZW6Rr6hadQXlHP49lEoRs3gtIEGhR2hF7Tjw
v+deOH72KIwkF37e8+uncpHLfK2nLKhkMVG9j73yXEhEmfnXmslApsCUDMlhfdoN
Yp0WOx2H/zMmaBxXUtEYRHNof1+6wbF9UX6InIadyeEhWu+zcOA7B5VEHeQjc0/i
vIMn10L64D+dgMeQwrWMvLgIsOHyaqDYZvAg/n8Sm5jUqWASE3v2LZpBCIZxkZ4V
1iDOTmSg1A/KKJryBN5AQqIezriCyxYcUoNfpmVOv8xJsrObo94o5+6Bj/UIN39l
9iwchcRDPmYQy0e0TSB4o3SskeZJG5AQXquiBUvpb36jlVbaTH3KnZ+ntJwMGiKg
UGSitfSMNalntcAthQBo87Iev4JfeFKEuEcxSGoOJia0cHadftpTkxFifNx0NkIh
vaGmBuDKvjwOmZrvxS/X3TGYZBosJiensDX/5FWplNLqwm9D0FQWp1j5iWtfzmW1
SwQwaCk4cXVOBbfBWa0L0xmZBwU/X4UlPLGE0ETvUpIwrn26Y3+eSZXGOBByzqec
DoSwU0da0PdntNSq9gc5iEXKrKI8UvB8V/zyLkFEAQq0+9nElDuZWpVYpXAwCkyo
IkDOCu1/jMg5SXHYNNohBNGGb9d0wh6jpTx5+BlkMDLP/X/RKqlihUh5XFuk6Uyj
vLdqfmU84tlgoAF2Y8lNanxtR0PATdB4jqWCFoKaZJv8FZav2cvZPmE84D0M6L2L
cFRjw62SA9sySDkqiieefOaWhpOdEfbNT+DBe1zflZTIEhp+OKBZ3TJ8H/zynEnn
EbxyC/jZtvLChmp5zWAtjvb8UDSFFJ3MlkCxpjvHO0ea+TMT5y0c0TJgjSnTGLao
cKABujsojtGMw8+jW8Bhfd04akVSuTkZf/Ma49U2InBlbWhNm+UM8zr8IqCtBNuR
STGdaIcfJcehk8K1aVWIleeYivB0fCdPx9cHzVwUIWbhhRA8L8KASiSzo6CXNjVe
CmpsQwkvNJbfIS/X/CO8JKlmdMa/97Dw7FdGWbfAClmfINi/LXgt4omsokFNwWcr
xVTudynRYWrOiFEzmiss5m6oeRWAgWk5NQqXRrUvtGrxIFSAc/MIWhev8m+ggv2i
2NSkGU50rufl1FQGR+f4S0JlVI+jQD6LdbvKY5jNLSQGiTzwDxcGKoQA6LvdIKL8
0WbbB2BsOH9E8JOyLZJvm1Z4/87fcvZ/YtSS7tZgmwQYnWuRa56pE1UuK1rTzI9+
HisYfZB+fWoJHmL3gnelTs9s76CY/SttxYFLXr3rH3MIDc/vPNEyvm7dLCALsTwm
53hHIKKDU/P0dKVrQKWpE1TkQG4UBDIwrkq/trzCo1thd5hGwHyrsOFS39cSqFLw
HeiBWZK3ejIpbomGXLxRaHI9fQQyIzSqvxKglRK6MlQkHgzHAtuRnVwVp8G3H6Bi
f7XuA6Q1A4tqKIGYVDpVYheyDcpFEpNwor0pBCBRiHQNCdEuOz5328SJHHyKUNJ4
1DU+DD0gFwAo8Fx6LxKfZHn3/Jt3XbrH1IEEsxeSTZf+49jOQhjrjQgoywH4v5u6
pUQ4daG+SeEi3eIDJkLotycUZAlbF8dchdKXgTQNM3UikEvxTeSaIyge/SCl36EO
cOSdtyccijR/Mr/a4m1RJ/cWMi+A6gx29yY+NjUvd4KfSg0IAoEcyHpslfSGZ9zq
+Hn+8yDm4LbUfxyf6xvu7Urb8RZB9SVqxcKAWJkrO+4q0NafGWtz9VReBQAZ55fJ
rrl4Vd6rQef5nIpJ1vNoIBY0+eKua+hvjZzQwk8ZZvhG+4BkEtIM6wDE+rhg+Q65
bYtZJ9zr4EkngIVLo2pGs6r62AfGdT+jkd1sK0o+7aUg7IWY0fwGQaVepHa1SR4p
Zvvr69pXpvjsVJ54qAyMFDVRF0eSM7MurfHb/TETcf/Gr8bODpeVzcCOVk4RI2d6
MAGCcOnLAKVgKvpueaEZzi24KkEOszor9aldpxtbZTlG1dfxtQgiElOeM/drbbdl
Jo1XJGup/PF1HxTLnVdqIOhnFMbRehvlaeEsBp+O4923jUlPiCIsJUEB3ng+yHCK
2m9Nt5rhm1iohm4Ia1Gh++daU20YwrXL3/UvmvjILGiWKelW3UUvbyQdPrbTeRR0
YZ2IbBW8F3u0EUESIL6jNUpV0XrifRm04gPPINTM801sHVv9TyV1TmDQjyH3XQdG
03WcHn7PmgTSH3YlXgtdc7OJYdlzDO5x+liHzF+WggbP8vsRvQjCQKRgcf5i2ikF
VMRWc9aT6XuH0LZtHJyowI3ItO+GFyvkX3Ko8cfI+YZxObc6uVM5WpAPS5/l4vz5
jB+9lGCqEHjg3R07YyHPOhV1rvONRievJ5SwXJl5kYyJsSQDbohlsQ7pnwCAbOMv
NCyX07uoco/s7+GtP9pA+OuMmss4v41X/A/tAEbSHvmcmMebzfp+2S0ki/mo4FW9
tYBvJd84BYgjD1cMrGoFCYgl3Y8CjN5QNg+CXGvSKud524Fq44e4UvkzHDw5oQyl
j5Gp+j2md5oBERINoNEbz8QO1yOAZioMg+a9pJjde/2AVULDyUiXQhCctlerj2RC
IqB6Ay5qkhJn4GO96No7Qb4C+Ai/fzsmuhqwnHseSaU5CDsstBpE3Inoj0I91qMM
j+G/pM36+D50uBhKGMF2cFPIdWJxh6xDr4d+5vX5Xjjgp/T9fRYEszTtOk6zVpw4
t0t3VO3UPIMJOgkk+j6sF7gaoQDky6R/MGaC+hQZ25iYtrkmgfDEzkHDEuzmVQIi
6IAMwQ4LwVh5wqvd1jMhpeJt+F6W1SK0VaolI3zZTcBxiPdrqxABD8/H4vDVdWZv
dNUwpi8ttG0lUhtJ5E90FfGTPMNPUzbAQJKN086Uzy1Axuu0m95yZ++BDS52UdQV
ehu3qAkcthhFajRgfNlG4PZrc6hDjqMonJawXKgn4Bn1/RRaEQO3tiZiWUEqs5zx
QdAVVobgPazW9N01zVmSRWQiNKTb8l/aeY4zD3ueRBc5IZXYX+Jw539LfE+NQzl9
0OLRZaGztKvWo7B04Q6s9U1I7gkzog80EmIMmicAgs6wh9OVhN+aeX30tV6LDHEJ
P071omTCvczW8/JZcPoDzFnCqol5T56GQVr2MStU57hn+SaHQRziFyXVwIqGx5sA
wggx7omykHHRHpFXa/yFItvCCHUlMa+aIRXlMg4ki+MucD/RW5jSD3AgjIall4Av
G9RPkC32PEuMhyu7TaFKDAYtE6sjZ0uUYGW+ppVOBF0nix7xjlNfmg4goxlC2B9f
OTzZMQHCreHq7ueXvHYhUrm6/ISE+EOJPPf59O7JDccT0K2oYMUADUIezF2yvlgT
/q6L9sRRihp2Gs2W9Ze/m5VxC4V34QdEFJ6KdNZwBwlTYPqldeCPiut2e3S9OjiI
HjkzfoQfgKF09EE0OZgDCeqsCE0AnariHzz2vl0+9IEZyTr/ehbRBad5yqNSkuoo
PsnaYC1sq9dK/Jh2zNA5tqxno36A67nBNCJtFEwYghmVMjOu7PfTuY4F4GnGY/zQ
KS7FHS2hLYwNBktV54J3Hvw6Wp+4d/nBmAtcucjYvnJWZnWVFvZ64Qkf5fe1l54y
SvAuOFFKe0cPThNA4McB4llXRFWRriTOzj+1eJnKEOyA0DmonzWID0HI0z3Joytm
TXB6Z51zQmZNfOkMkRaaSx7EjffOzh1WWViaS0tCsfIYyPNvuuW359AsoV3oC/l/
Wz8fojxyxqvopToqJkIHF1O8kjV5sl1r9Bjs0VQDEaaRQDhP1KV+uZcn/J3XHnZY
wyTOe5VOtmsOEo5RpuNdHBUZ9egbWSi5YnR6XA07gcZmpUlmHBLsvr1reZXhXBA5
wsnYav1K3Y9HtHReNZmsFrf4raO8V8W/6MtgL9OKsPWVxtG9GcFeHu1S0GUvF30g
znPDkfNiCMF6iPWr6HGwcNHzoqukik9/T89mcSg62zxlp0TmbnJOBY+7WUu1K7Df
IMxvksFHRMzyqkybhYC4HGePh6avFkYXo5V1b9stRNON8PBu+GRhG7ztNWNThbJ4
xgd4uYnCtj57g6X16s31xhY1gO1SmP/R31O8oztGnI0H4jepAIzIS5kzEiw0Yk3A
JF2bdyWmfSUVeOMCbFNox2CoSICgzU4Am5EV7gnXP9n+li8V3KcXB2p2YjETzs6i
Z8iHXq4AolIjTUVZxXjVV8xch4Rv7Bbu7huO5mUDIjFtOxCeseTSPhosOu3i8qVN
+T1zuNxmMWnQJJ8p8cNpVio/Bovy/D35BwpKzdoVeVJy57Ur2+DJ9n44Lw6CwbJ5
N045zNkpSbOgPgBJeHsv2M9fUMWQFZBltYcEsHjKz2UHVqKltrz3pZq5kxGfDb8D
L0Ui+gq4aa8AtU1gBk8nl9pQeNdao5bVecUXrHHY9c5Z7nO6bWcXcsOM4hSigsqA
Z9E5fT2IyMvLTKFU59BygY3WwWuRfSUTJPJzd64LurGa8ijS8LIZEXl/1Hn85CSh
Fb5HsbzIA7tEZmSYuEG7Fg/7n7NiYGpyGwoe62K7a8b0mG+e8RvLdvZqviVUncLY
ODJJS4BnDYwUtda7FY7V9qYAmK6prc8bjvONdexFa2lTTXHj0VN9MsPynolmjzF3
J5NptdI5mVbvcW3BRo4G301idC+hFciEJdkHrRSiscyYQDrRAub+IGROErVBPSY9
0dKyT8Ic5+W1TAxLSMX9jfXToO0yi+tHm4YRuD/rv1qeYLEIcU6XAxZfg9ewwVyy
iKY7mpGMoZtXXe6FAm+XEM1aoDnnhewEo+l08fwX574V+3BpyuEN2LC6pqOj6tt0
aq9TRwgX1a0OO6sSMMbrkRy7ec+vyPVYhFYuMyvASpEHx/e0ghHd0mARjn8+MpJW
n5IQFubQMkazlW4w2Cds7Nlu8712yurdZP7ktikWMecKie4FJj95FZUISCIvjl28
deHWVvaDuoEEyGZu6zncsGGQZ6t564nZBNWwY0cWWySFf5sK/CRBYvqHkrm2Axs6
yURVa0ILSAcziN1uLQQvU43/Yt9ztxbdxzOXmq4UE1gNG9l44WnIpOueJhjkBUMr
Z7Qj/FCGty0HxjqmYc7V6y4DBWIM4tNXlvTcgGjrgpu6Zr+8vJBQ+Tq44spT1/IG
eUPshZfEZRnqDWogi3eUJUhRAqcsFBVJwOD+ZTZyykIP5OpfSeglpojFyWsYI8oi
cI4nArdFzDbOLR8AHHd1RUgovSIthkb+Y0dMFpmDjIwpwcv320SFB6Y76tmtPxhp
lzGxaggAuLnIAidbuAGEhS9fPkgxB7pJWdNMJ/mzptfv5tzI8G7gqHBOdSZM3Rfi
G//MNVP76BDNNBUIhM+fvrGvF3qjeaC2tCIBPGiWtSlx9li71HcxhmO8Z5CcSWZP
d6tsuwUeswCSqoosrcHS1u5npTglZryZ1PbS+wS58MSP4dQY/ygtCWceVwFvz+mR
Es/L4im+QoYn+38xkSOIycrZn89TemLLIrPEzg2kw7r7N2kJrkybQo4h90ULaBRO
bIG+EjFL7qleLgD9EuHAWLwwB4rbmb9A+DcuLekqkMtz2enQr5q2dWRmhirrYWoa
TSVA5bGNWWYYHbi0G5Qj9hl2L47z/cUxN4OkOUuBeigci59b8s+d53ZwWRPreEfI
k3YlnNZVpAay3cNkXlx81HXskNSevXmEt9bQpnYI60DX+iUK8IUMhFubADXIWnWD
gDelJK3U3jOPoYoQYCREXnmyK23Jks9BRmWmGvVUTDOlDKvTs9w01fTqCn7tG7RE
ElFZO/athQo+/pNQtmp6XCiA042nGRfmqee4H87cNZ3D693OH2t/T5Ew6uY29Tft
3A/su5KuxAN+fb+956teh2lAtsfHekP/bX0x1yyRNdPfoazQENSbHq30yT65DOdk
WHYMHeRMgp8vN5PPywzl9SwQthUeuNZwvbX7C+dz8rm4LnF2J2Ko8p5iDe6dZr03
zhGewyPv+QtjjtiHOxFzPIBJgylRkoaC39RrVTfXJGidgMd/j5m+pBqhoHUqILih
uOkge1yAihFoBtO5JJ7J2ZzmN6Z6jd6A0yVCuNPAZCf/k/LK0ZDffqPCnZhF8hCV
3zUZphFcFG7rQ9QXHLCz4n2z4fhn36Lp9AfELAQ/2RZJJteglJvdJ+Vz7jKTjdT/
MOmdQknqWjeUwaGjosXylYUUPZ2nZ8v0LPooO8UDyG/Dv5IJ4WIHhOBG/geDpan2
+L1ee+cafLwvrNcBy3UKjHWz+tbM2H3OKElnIIYUJCdfoXjaCGxvYqMquu8syzdR
RB6idNd3ONTKiMbRrJT987mQumuKu3nQgOxzycLYmaNMYFhnHF3Z1YB6dc6pQTCe
oFx4Ap2fKP7auDt7R3G9ETsLhissFz2b9rMc20qj8lIL1Xv9oLPX+M6wg1+EpzFW
2Yb68OUniV0FEgbM+ps9KDiPpnMw4KoVqKONOKzppC1krExrf2FYzNYi91P0imdF
CtIO+/MAPZV/bnjW/I6hBXulaDw3o7Z/NR/DA/EpakGhgp6NuYxpANhY2piKvyGL
D60AP/DaBuuLOyi35JBqqOUpJhgRrclr1BLg6/E+9Hrg+K6cSKm4UpBRkOdpsZF2
bbb3dTStiPGOrj0VOzgkNk2XFLDSigXzmZCurf1qJQYvIJv1Jexi9b9icxNs1zvW
rubEEM8mJiw1fKO1sY28TW+jQb8OKdPYcHRxGomxBsAwuvK/zV/ryJ9uMaXQLKfS
59Rff46UcMeXgjBCBrnoaNwamTf1bxHOHIwbBtcqwL9aOx6vw+kuA7LfRPtgzB9R
zSEJKY9vmI7fcfjSvQ+7CjEfpBP/MA7rLN3VGx3nbcUxhQ1K8UJS/T5LJtNSjImg
t0paKFU1vCsem9804OS88z/Dx1FOTHiY6gPN9Gh4DcQl4TyX0atbUig21Sg0oTmS
B/GeK0iE0MiSFbVYmzLUn5uij/GAnXytjjjub58QQy01Q0r8wjLwWuXZk0hjxRCl
4r6mw8ZySeg06IM2kcZyztHZzCBPqHnlikkx2Iwq6+VZcymsu3RbMqtRvmG1pEIV
7O5dtAR8wb9i0RV5OemUpK6uq9DuDahl/JARvmiiV3duhtZUgSSSrUv/dYuH/yU+
H2xIdBnFOhWO0VWEy8mIFnnLAI3xv1GTSPNiAKiPHO36gVBwIk2UiU60vZ/kGhMH
ntl4iBCDlKhB/1dKULlc3IKrK8ZJbHjn9Ar9nfzEZH2+rR10KGA3HsBtP61OxUvu
ffm9jCOYD13JnvA/TcafSklxi1UKsvoEMYcHcBEdHnq5F4Gt/RIRRJ0iC1OeYZhA
CmUWa1Mgb/VzUsTnVCIH+bt6ahHA7/4QMnWJpNj1nyVyTGbJAkYiPOvJ7WzGYNOI
8VT5y4HQh4y1IveGqLqf8lk8yh+rlcAlZyzGC7ybOSoY/49aU53kFhrAN7KKbHmo
3qXHtyjUTE9s0LFGg40wRXSLKSameBpMPHpUcfjcPhegsTilbXFfwLBhi+kZujUZ
ONDev3yLlDJ9EJQzzi822yt7u4IKZJndVp088Tg4QnM/qajkow3hSIso8KkVCmtH
6o6pegVgl9R3qC8RM4FzYX9/xoxJUrwX00D5x3hs40HMB84mb2rDemG3vBHYrFHq
h5ncY3nfkNqag8JYa3vhx0Isppn9BnU1RPDMbzv4dMImk7QjREwvdtDLzrAmHjrL
6nbSKzllqcqahvgswwUVJ72H7tFZkVgfH2Qd0W2mYt+ISElnEZ4sRjl6wdjAe5Fa
kQTYEM55FcSZ4W1+q/fqQSMqNzY7BcNehwjTSHqiX2z2cbDJwRofzpXY0qzOuin0
kUiHMnj5pZLkNAZ6dxNw7TN8ZsDWm1m2QyPwkjKDWvZRUhC7yKJVX8a03WGmAxFd
W+0s1NVjNyha7UGYWId9ivgh/G1rlQG7OWzoYfDoz6dMc8Rh7fsXOrElUELhZbQa
2MUZmWgi8Nv3vXyRWyiPleiPOlJ0BOfqZtUsYE8maqDFBD5ZZAU1cjVClV97qYYS
RPPHWHNfyQ3K4fzRnUR9CZxZ/KjZux1UOCBmW0BBvJ6uvMG3cyLD9iK2DACiwK8q
pwwrYbnEk+4SvS+TjzEFBurZPdHOuYlyJ8qVDgjHyeaK4lR13gPwzgI2WGW2FajB
2yBUMiNMvSwB4okySWdIrVygPJX7FATreuIx2RWX8HjPy3x2z6C78wUq/x+mWag+
o1OliI+nzn4CufCPmx6y9Qm6b2YuviLEyPRNijSKBLUdNvJY2LfZfDyY7p+DE3k9
cTkAxzA32xOYUXzE6UguDzYr3ebFarFmnGV0weHUsB7tMo9cQsCgOGoCSqjDTYXq
d3QFP/goJldqGmpUNVn/OCo2Y7qyXxH+xetcB0wdLwMmjGRXO4LY2oTOEEavMEdn
9ImKNWkiWGKa8AoSBNwGB53YoSc5Xsjj4SCP8sS9Slii4XqoSV+JlgjAjjAHTQQO
awu/4/TF4pPF7PqyGl/1fJOuATOxWkSUSEVVwK+Ct/ercHEjU2jpaD8tcZ2BjlqM
3wRgTotjkSJThvqn493KCtfBkBcaDi8il7wYwtP+PB/MHFNHMJV3M1/yvQHOtsEA
urY/pp4wSQpAmHuVFmfFAEKDEk08ZPClgc/Ktz3bT3Ux8fO6Y2EgPd8uu2BqYc6q
v53DqNk3eGUrjABeJjVxxl1lA8HPhxDY4yxJy6iyQOnSz6GCe2hggpHmdzQ5MJ1Q
INMBdh5rCmwYltc7akqDRiYEpsaVhyE///xD9daottcRJXBrLCruTx+oRqS4b+sz
cUUfkw4vwOGGIjXQglpEOHq8cbvfgnBgixOoQpSyqj2LUGU4diALrBTUyvL09GQr
e9UThiU+GTqb7R+UBkPY9T3BotrbuQEDO3d96lQivDEVXwXXY+75PwiFTeeAMpbw
9RH+i8s/hXJz9oFBWBKDaTaHbcaaWIv9MtWdKQYqPK2Zlgj3N1SGAOHGJCqOYiJi
EATbMtTRWZl97vVG9O3jZyfdIAslcFhtqU7gXRDnoDNeWpm891BhqjYzJOA5OSta
YbGGm1fUazwKnocWaS32JjiJr5RbEmwtNbD25kGc8hEUXXw8N+JYDZBjpcUgGyjz
BwDEPyigZmkmKfHl7Dka/PdKHt7aM47qZPDV/LVsoPWKXC+p6SizJ8H84aoEVXbf
TWecIij/kN8WVe8hReLDbL6ODJ3irY1kgwejwGgWokS/aOt9PKlRxxLOpRH822tk
Skp4RWw8KfPTixrDgy3e4vKwJHORVdt0YRxTqXTiHBr1z9WW4dRQP3bNOwUNXNRe
GEKcu2BPMYWqsUUn2Cjy8y7hHwF8qjwisO3Pc7DIdF5r4Xa0BRQrRf5yRd7RzfsR
+HYelXIq9JixvTBK3/n9bV8+y56F5Gnh8j9otb8fvRd6NwTkznyHQgxKv/GMLOhx
RpJIKsyPLnTepcP2kgONuPIsN0BCd8zftlwoKTE6CKAefk4dBKo84LAdnQ9RoTyc
e9NQk93o/w1Uivvir2YlRfbj5zEZ3C6ISmBjF4dk+teMzoP2Ij/MOixw2aaysL8C
UmuUNq5Gl5kAZXeXwRYwi1LpF/D1rWVSwWmmppiId4cPvNtd4jZmZoWIkRbh9vVB
p00Ua10fG2lH1krS25d4DAuDDa8qiMkS8Y97wtGxwdFW1SThvCrsvCkcURZDciWD
n6pCJ7sEB6pqtY9C0Yw/qpZqhiwBRYQzCjBTfM7k4ljbgd03fCbpy69pa44O+ou1
UhWp1pt08QkCdU6C28EDx5vwPHaq806qqMQMaFS6B08x3cqvGw0hq3U3NvLMfRug
zktdfaI59ejH7E2vVcH58UTxykiDw8hW9khlSA1aNf1YPgQ/9Dmj62Jb6qiBInal
GErjECv7obBbrXBoT84ZZvDq5inD7Msjtph6Jdf0Ie724OcZEUQnERU9oErn+uyY
OGlt91a/AndJGNmrAch4GRKla0+oFNxlh0+vKhPCtRwWphumRM89CIh2QQ87pJ6J
t8f0y0mip2huw/tTDrttsrjffSyGBhHcWA5isFDt0eNr5MWatsinEGH/GItD6oOG
B0NOniDa/XNY8d8wULXmOo+ZkN93Pc3TCMia/WDz2tEykqCPRh5wOJSHtdUzrk7U
oRDGL0aQ4plW5ZYR6vOBUfJF9STWkCqvBQZyyYvtFAYJdm9l62POeVZ8QgfMJZc7
Iuni1WLEEC3TMzuWifJoKddwCnQo82Nf3tOMOhVtPV+kVrhunfym3jS52G43dOG7
e0m9OJAbiwi26QHQT3276Gx9GInGlpaDPltVEnA2Sx/lKWSeGFMgWXCS3TUuNKbZ
Wil8Ks+QLvWUqk1z+KUVajrqEHf29DC+ejOpOBp14uNjvuyAvNGvUEbX/FlbUL0w
R//3LSWEjLK/xiZp2yPc4I5Gc8GpaT6gigeql4Ci+kAB+UMlyaNyZZaESulphjMP
Q+p459kXfmRFmYnCQFTFRuWdTSoJNVzOhYUu0AzPcIVpXqY/iZjDbRerSqAPu1US
USQSxOzLIT80EuBbEZiYaRak3uMkTnXAg87q6eauC4V7cnQwCtsrtg4/6B+qiV3J
Hi/HZ8BeB70ScSq39GPUDZweW2IHGLoINZZRwP5p8R2EqpF4ejOjgRk9M6hdGEFm
uozMUbsggQLLdXUCNa/YYDplCGZsuJTCh0mY3KM9OSOqKHwxyC9x+W9MQZHawGdv
FssaNEoR9hODMyaMXpnbLmWEGIA/I0jR45vtgFtLXVmBOQdSmTyq/u9KEeyI5nmx
USJFcD6C32bgJoF/WeDVupWJWFS36czqJHtoFnFFtaNvr4bKv4wAh+VQfrMz/D/1
64dWA7JA8M+aeygSlMIqeQsRVs+VKNaNWkzwYJC4/ipXZpRyBscYdBxHg5AI+SsT
iqVWJEEZLc3EE6FshClpiUuYuSHaP6g5FF+MMk8fzTkkIbiIN+6/e+zRvukdAq7c
vP6D2EN0Ta6lTSW28BNJhyDrVB3mPAPpte86nBmBZkddGgLJnh5lfWeiRMWLvxqU
7oDo804SbI0k9n1I13wDAzHSmIBuPsJ3aPUIFV4MNe0DfBfM7GsT78MomLEOQlVe
epQcOUE/d/0xA2krYhjBXEzuYsOX0PCRc4FiKUbJ4eaKoyflotFOmMltCFFmwGiw
Hs4vhpjs0N5o1pFD95ja4f63SwMOZei3biN0M5V41UMfmt7HxRYWBSc5ImJNq2Ob
bUEoBhpU5LDGh4XG45ENkVmvNzrFsrN0B6CzkMtDIZKebQUSKprTK9rvbhNx8e5N
5FgGdWPxgIJJt4G/xlEGdEHzyZ9qSASYGT/zggQguf75Sn5OmjAl0qwhxh2VBSe8
rudZV2Z81+gsDhc9NJHpTjCFxEj3DpeQ74431YHGz7Jou2nNb/CpiYhF3toTkhgU
w0y7XKqnWsPZNsxSMagFzOT8r/K2oYHKD1iOmWP0XUNSUQlNwcadyWTdIasno3oP
7+iHTg09oBiEwpTc+EUo0vKjDkaUcMp7fDgKNXpYw1o1iPR+UuK1nLP8nVPmBiPT
ybmyrUQUCiWpCttAFNwuca5mlD4WbYk7tzE0uMIoBFgfbLpA40RDfQ6E5DdrqgsP
fao9rEeHdoApc/r+JWUWDlqc4C+/205S5u05ipGTPTarUasQEa5xbNVwcS/s4xbc
yXWOIYFV2O6rRaRA/U/NudtWoAYnqL2aL7BcoGqVrthhFmyCyl5C80RuGrcKgTaz
KXisBsxEIsPVNxZFTrlCyI4ePsBiY99hdAlAvq2Cu5d22596tUUgYGshGoSTWWxG
DLizM5xvEBGPGMBXVwQ5z5YJtRPoeTgXyEqXHtIQpsI/WCMMmnZDOdllUie33a8e
y7t6x2ck6uFzEVHaf3f+QKefMzvLUdfObtQjj1Ntsel0bRmhxmrEpRuHZdxsqqBe
FT1XQ93le6M9oXLJhErBQNOwSOai9zoooKNWE0N02mio0u+1IDYCTjMAoduOCviO
dt0WmoSNu7ZwACZItYNqUpdpnTWz3NKjLZeKc1yvvauZOxHxfwL/bp9bKd0a6jty
kKYzNdJ1Y2YXLOKB10MnaEpIW3urlcClhviBwA1PcFQMbTFcqMT2kZTMK8o56k+F
2wtgtBiMHyVkl/B7/RdTKtRgl8IaeIPix7Pebzol/6GFdCyZzb0vB4A7RCeHOsGl
yheguioewoWgvH7KG9pbOq+LMs8smyno7H1poJ18spnuvcvfI6YKzdz8c7zLjKbj
Lsbr1JlQfamqytVf/TVuCuXX4rfTD5WP9ZJEGCIFDa4mTdPUDi0kMKDFwcRewcbq
H0P5zx0S7Gtuuw7sYpgbRgcnOAPO+aysfDU/nFP7wsIedltIRj4Wlk2GhZTEiLRT
m/ARYzBiqrdQ3td2/b2G975CvBURpbn0+VOo9wIQoRE8D+kWbd0ESMDfasQZXXjw
b3szHYUQwmgYcVOkUUGtZ9VLETV7szaNGzdZfT8HjHXpJViYB1/B76gWGe2OzrHN
aBl0mIXgUcQcM0r+gpUKCm65Ia5WVQtC2LQU9qkvPR6SZDXn8pVdl80ZpvX0d1lz
sLoq05ZoIT2MxWwENIc10x27RZVht/U92YMEKz1Uh5BaHdjdR/LCadfs1RcJKcdf
TqPcokZEzlbidhj52bpvFBH+9P9NUqftZqjvVJewtXyI6FBCoTzc3w2j1QGAhCyu
X72Bf0TzzDPVG+y9fNnxgaTIYMWWuC88R1uMzQ/72GfZPrUnhqhYvV2cORyLNOTS
Q14l+NqXDhMS5RAUqXzhudvEO90Pxqts4mh4pNn5cZyimxleMYk03ema61YJnAwu
36yUXl7V09+3YwttrDdI4xv8AIiAPllgfrcBdsi2jffgxY2Mt8N8PMsfIlanQepX
Xy30AnFRC4g8K27O0wMeVIt00JDC2A1TBZLoWjd5VCXgXHU8KDg3q+SnmAPQm94F
kI5uBctxhd+ar7/ZbbbyentmgedWqBnBn6sMI9SrYG5zCHZDXvqu6TsiwVO5r3gf
g4ByLnwLN4ftOKpRvEo200eqoP2ZTdse8fj8gIip7VQaDWnI7Gde4tSxszMsx5j3
oZcKZDLm3SF0sJ9EIJOyA5hsOBu6k6oaO89aK+V9LBHIzsgtKkoUHBr+pG2baKXi
UlKDXoYwGvCjaFd/sbZMEEeysZDDebHZQEBOqpAxtVGl355lMs1jZjnlRb9QbLZv
h5HHwX3a6qXSSLlFqDeKH5YVD6OkrCeeDvuzvwUoQDBKH+4/lRTSEeUJl4j5gHXd
nGOHGFX5XGJEcvhWy2gVeV7gvwwBwnRY0TVi03R5VuhBUVQY/5EBwwiwKGwqbbUe
NXh7ExSMTg0o/StsNeAUd4VdBC8WACYn/GNOm1Ou8UN62uMwFPCU/ij8II18w7PL
YlMg3fcr6zlSMAB2R84Xog5CQS6Pw8cDg5ZEkWIqKo/Lp68FntsYack2Uf3tARRU
R3oalfsE3FBD37yFAEEocYnQNyu50IVbkL2+BaBEOhVw7fDt8czPSMV5yrzt/bC4
85oR43wHEnXkTk0QLMlDuiqOLtSKinBEMCaprLlq55kEBt7Z5dEOwgUcLuL0nT4U
h6JUDj4NT1yxxDuXUmobjq+pX0q13S7nhVjQWUdoXlJC/n4yEzYcYwlSiBTSV11M
hiH1sQuW0eOrcso6d7OFTrfLahgsHFbYwVaRzCtZtvBPKbSEbivYnPSJAetvFuVg
hsuMVH0SYpMbZhaJUsJueowY7jXibWT4FJV+qeOCwKiN2aPdiEOLcByGLbaIRmob
ZbdIkqzDDCtC6+OGORYuMtaJEsIQAH9SpL06qVTt5v9fQiMCEWgdupe6J+Nar5I7
teqkMj6k28sPOqJ4/QehozaGL4GQ6chopHF5dgv0hJnth3Kem1en+rlu/pkeGmgY
JH7pbIcdF2flfHEQYOL653yNe+ZfUKaOYTBRvpGZxknzJBcUs8EGz7PIGhVCaDmG
H6bNGPW/EUDF2zhFsvEuw24LVF0ux4naiS4r/31MocGtjn10ZvfgrJcLLA8irD9T
EMkojc7BLIC1gxtNSJK2FxU31dFty3P3ROqohqsVBq1RWNffG5hU5X7tRlXsoueo
aBTtFsuY84I1YWJw4wTVHWJpWef8cpCQlPucx/i+Gz2NAL7uET1DY6cnymtaq97f
3ZjtBG8if4CePFMbgzFW0+xHj3Vt4bZXopsARuHFShgxyg3mzhCih7uYXSO3Rr4x
cwSQjo1aKS4/cZd74bFI+rd4RH1U8O/60DYi8BoDe5HzteyNWR93pLHTNpmcUyKo
ylyssh17bELStc7d4KKnujWyYazkKTzAljIPuZrDoPzWIa49XPOhoow+IbvQNBew
74MMwi/Mt5uIbupO/BcBWegRWORmY3/7ZbQUX62Kwu6gqHYKekBcSrX8a1ILLvJ6
IbwvGX0h5K9ZPYUpaby6HbzaRHHvfwig1OdRQJiQtlDuaRmJp5SHxNyTQE4A0TX0
tN3BquOxS9rA1N26fMASAHJfJZcQXyHfP7liuLlBvWOIogso7DKQSwmA0eL4JoFt
v0OPuAx02ctNU+jWZz8oB/hSeOouaEM23waRVwslnFOxKNO1qg8A/4mnpkxms4ML
oVNXWPDSt8haYlRagxqkBZj/DImBqojIdOJvEHplCWNUSpOCWMtuglA8IFP0f/kW
kyH6UQ5IkRrVlGQLiNSst+mHDmJ3vx/OtPLMasLagnfO2dS4p0ydqx9/i2GjHbg3
io+oevLtzfksHl5+PEm3RJZKm4eSOyTQuR4m+0vfrxZ8qi/Z1UQ32sa99sx3tGFt
xuxvmqFqf3NyeB6sDNS0XK/NF1L4xrXDYtE3yLQbsKRj/TrNw83nmOgivezFnlkc
xT59Dmr+k1vRFf+ZIFWJLvfA/Ytc/R9vPo0atm1JnJZ9J+lX0Vo3vfhgc1ejnLuB
r/fB00vF6/knegt7chD/npFCZpZfodpVMyiJwLxMXZ9Tuen9GhczjqRywuZSPkGE
/rfqJK8lrDaWkaH22ygXFjsgZM0kWG2Qw0too5+Ybu9YQCTw9H9QGc3tEgdaDBCM
8+c8jaV2ESPZtmb2P+wnrROuekAMLYIT9dPK1LUTSeC+0bGMqRzipxa6vDkmZQdN
5iRJv/a0jhp3i/rULJMKm/YQOuTjAjHHcGItXg5aQPXvgx/Ivxf2YR4hot55UMdb
tI9+wdKJaFQsNLlSKPqYexKVnBwqVc2hgLM4375SEho8hQUWGZPXB0avBq45l2lq
qSUJkmDnbHFIQJrZo5V0/YJIQRi4Czt34hPZdlWAiPTQ7l98r7l5O6NCOxBl0LpA
VM16zjjKb06PQ5IESzaFtsOU77HQm2lQJLolUulcAIs1JA+awc2PtdBkCrlqlTyc
4vZevpsl0Ux66GL8SIks/dnv37r4x/0vkKO+2HYtJO4FlV5JOziwX35EQEdNC2uh
QwOIX67F3uvOPijIghxMGgv6Bfb3/b3ICX+VNuKR7HGWjX4H0TmCmyOLQma/Fy3M
K5blhUAXR9pFQ4IKt3GGV5cIGlPNDViAhvOQ6wqOH4IE+WuAXosnLdDPdTK+QGyk
/mM6VeApgB9XlGrh6P3HK8emy8/OjicR7dSH+uKNCBO85H/cZn6X+kHa8/fzGeGZ
cn4VvnMaE3qtWC9TEgtHzIGWgq2Br5a5dca7cb6kpOfbaxOY/jyMW0LMAbB/faBe
XYxfiyAzVVsXOJiHcSZjgHV4utls0d6PxHBE33RgejZ213B+1F51QmPwmp93KoFO
g+YLxkbbpum1Ir3yzW4wGzwF3gDd8oONIlWLkND9T0CxjwS0KRLIcOETVYbZiKnG
LaxCN4tE76svgVfdVEhq4x3q65oylg6MTrxU9Ijd2sWjqvXam86qmzWpfXSWBg55
htGpgAHtTXA+IGwO6EvL2AJ+jWXaKm32oQXyDEVMGQ9ZM5G6XskAFjrbicHi6928
M3kYx0GZUNhtX+rLLjhFZljl34y29sftBP1mj19Cs4IqheF5cYIBtZ52qHIuvlPF
6NpQXuNlQa3Ce2wgRXGkaD6iR5smF4/DlOkzMSk6kuvg/DOEqMyfaNtIc3sna0iJ
0VBABNovYlacjcgu8O8d0XwhmhNfgAJc3t8y/LsxCLRP6wc8cHffeEwBRGnDuB5L
rZbET8I+DVW+nq8zP9BtKsoD7dPVdVw9vmkHcEw40dAgivWhb42gk/9Z0kuQFtKf
ABQkZ9gG9oaOmODPshQqUmkd5L2YkVgHsL4EidBfyltjPlplHkyZXswBrI5siXUZ
SPwnOauBf8sBX8lYw2/Fxe0UwHJdezndItQxZZAwq00TciyzWmRstuQlo1aEc4Jn
33b5NsLZQZASpXuSc7YDYMvy7N/gooymFCSKGyA9ZAvVyWq54a1u9GD/7hQw0h1F
FHCczcimm4HA27iZOkXpRppLYwxvJ2lQPZZSUSd6QrwB/Ug93LPmXoScQFRFMsBy
BjBA96eNODU9Xy56/YuNXDdE+MDWgutVRLpUt3W+wnm0AIdR4k2cF7JDl7sWYcNc
gZnuqKI0xDsywDfQS4ne4LriH2vJiLX6+AsTsYOkxKM5Fy5hUhpPyoR/Oa8A6oso
Lx85KnNWJRo84nzNtgvj9u6uRET/gQ2vzzHAI9mwMK5+T+OiGiMnYWboeg5JWQC8
IHL0jHvCXrqsRXtqLUd44AzImcF7RT3HD7fkRi1Y2ImIHZHKkoVqFs2SVk5PcKVl
yfTixU0HlSwCt6YcJZoBb9wmDFoduNGfW7NEH4M7Q8m07OFluFelLIoZNLQorJXj
Qs6ntVeYEn7P6irHquN2l8WQfXOP2esHrRMk7FVsIcF0VvxDGzVQa/vylfvoTikb
qo0qSEfoBgR2/7Qy95jmLxfqwfxBaWzutepLYNDMkQYP0rnxTU6y+BefNaUx/xEN
/QVsIf6MGFmD8QGDu5WGkXfSyZTEnl7/JmE2oRlZ4afTToO67usIU6CFJfbAyJXT
MUbgUquSVWkRSXfBwrA7LeLfCgBkgFgZFU1mRTJAaZ6P/Gqobvl+WU0t2NkDDfSZ
UZLYANvU7Gn2D9pk5vlElFtd+58YdEyzRSkMKaEzomGxosNCpHFynX0z6qYEELWB
QWwaIDXB/A0NMI9Ka40mfSCW7Zh6D2VqkfV/olYwlCDXKzaOMYMBqr5CUw8Mm+no
47dF/YUF8qoKNj5/JL/9qrcSUrqIMMQnwXY+32/93EUHbecJcbUC/d/YJBvkwkTO
UtibU5lqrnyaOkebIVCCcVtaOvT13OIVqVEE/bB1v/1WIrT3IK/BMMHyVxG068/V
gvtKru/jYMkb6TqWmfARRHkqAl5X14B/9JK6Exnhx+ohtduBNdP07pK31gfBG4GK
qaC6BBraZ+0uvzpFcPPWXKMBWIcqmldDAlMXFWTU7jMBEbuKcb0cu5h7lZ7aLW7L
uqYlD7UTG3KPTFZpLS8hhud6Q/YUJwmEpwAf7ZRTfTDHnfsIXXk7F/+qPptbfT5E
eUagWEhUvb508HXK54MJ41PE6tQI07jA6wbQ44ZtSg94NPQW1Q92j7oO+uZ2G2cD
L6qGyLgZa00xAwZKkjwt+6fdPhDxr9AGJ4zrPd7hVaeI23NuzL7IgsIKDA+gVvjw
SbEztMPwskKJnrcZRf9O9kPdw8wXMUwZY3ToGYp7Ju3EOWYCqoVF3Xq9HOC0YR22
Gur98vqBLGn0xIsYos5Yj8Cd464j8GI86ELDQcaBYzNdmfDoDxEPkJJacJK19loi
TtNM5KeZkAzm0Ea7PbDRGNeH5ZLk7Vu/UsKEaTjeGtdCdw5DaA4CqNuw9tnh14ER
F5m4EtuQ9Q/4RLMDfRKm6ZXtzZoDSlpMqs95FE63LI+lLmGRv6Dnq/bt42W43yZ9
n/2IIclKp7XRhgVETi6EuvYFuDmvdqHT8fkYa2A67M1wnX4qZguRZaczX0rEj1sY
nwNOs3MCURqC06AUH56UszB5XKLs0GoowU8bm8icRnS44yF8HNjvR73mrmEtGPfB
yjNHMuXfYdVnwCSHOKu1oOqLuMcJ3LACpWSLH2KRhtKnY4oe2wry/mYjz4+BaXX5
lG7P0vBJPr81jF4KhaBA0qiI6IK69gmivCsHHcDtwGl7ROTkib/WF26jQP0txASJ
tBFu3TSMQTWXPl/TPsjM5tTwhxkl/b7tiyFpthBhA6G3vU2pb/QeKmw+5bErjFDY
49nh0H/1YtWj3+8WPODYNx0mWN5afkveU82dYwdp+aiC2Xs7hUyczIGh6p8b00LK
g/cbud33c+X1mSgaewBXedM2wjdrvWUaqbTgKebP4zZuFyCNdTBqTuhv28Qs5HTe
MPbwWLjQbQKYgYB6yuaR7q4ZgcrDugNRofgN8Goni0PYjHctWi7ZdsGhcXIyeOJi
cm642hQdf7+raRolB9ouBkeN/K0DCFOJBjm5IKPz5QMUta66CwvGQzMSbmmd5NsX
bW39ig9ktbyyRP2/zN/wYKV+FQS3E/zc8dMESzNuV547lLM7cEJufzKFTnPu9oas
RVFaqWP1A5ZJ3TIGAsR5EmUY9BsVFLg296FCoRBik4qK1/ltvBPYP9tVdXtZqK19
TCpy6mV5wrACyfXg1/3tKdMg9DNaEi4sPbHVPKM/1gaQO38pCzoouYCkmveQHg+R
AkqX5dIFOo9C7XA5lVpQizp+I0bMBo4Nn62/9TeXoonlozrOdZpe5kO9RoxJXLL7
+VAZQ4Qf/IsPpKOOG3hiaVtyLDZuBnSkzb3BaSfrdtwOE2dkcBl0eoHS1UhmDTIH
htKnsYE9tsrC84wGLu3BPkr9pFeZIip2FipJ2EezvyeWTl84lSZFut6Nutey9Zh/
4MlZfrdBvSRVss+z4T5wfKLvYKoEuAO6JZ0EoUFED/YT1n4T5Vl3Vhliw48xxx27
G3UUmXLrPmH7xjr1jhyms5otL9e1PA8rVbes4b4D2KlyO58CQU05PTB1v6RoQvQu
RmxEqYEy4uzItWKIiDSbF6rau+7vDTWgQ2AZjltO3bTLt8da3Z9zCeR7JHI/dmb6
QzAxf5r8GmVjvB8Q7PRPso330meMLj3txwsOINqeX+r4OGpCiKKgrUFvt+vJDTSO
hVUh/OS1xR7FQI0P22iIsYyK0B1pg43tI8RYbRsT9oYAV8gWjFONICWlGeoBuERz
4ObhF9i5ZWPlx4JIx8vNBK0YMMWSMYnBGMktB7R8lFWv3HK5/jnqzruAFd+cA8zr
evhBlj8OnFvsUXh7eVi/TOigNBbhELGoDec4wPGBX9JQts9UBWtJcDcNT16+8ZDQ
0/ORjJ7FO7NGWptVeBjBGNsgEkJaiooR8k8/+wY9lfJB0hbJb0JqV9PZxjAFTy2o
e13+nZyNivV8CXtN4iaWVJ08QOr0psQq2bAVFMc38jN5J1esY2OQ3gACT7OTp6sa
x5nXbw4CFJ8yFXpSsyPo+BENlr/r5kHjmn7/RIGwv1qAHdr2fBPSZaC8x+5liEoW
wTxtWt8AuDS63+7+88B20GyKD7IwmHgkp0vL6JiPf1TiajqDQDvcedFOn9x26MFW
rPEU2LRZ43wf4kADkVxv0dQHcYagkDYHyUwgiZuJZwxx60+yYM6fBJwbXFDqsPwZ
mzqlPExWf/ptSqUnLrw5Kc2D5AMY5o6YM5c+aW4k2Ww/8+8kmzgDOawJ5HIMkOTw
OANb2DN5/J2I7lkEr+udbkwqF5G0FhBYzCOhIIVZ/CLaME0AVv1SmtCXfosiIUVM
k/X637DttkGB/Mm+qoONGkitsqqSYLPL7hk9ZOWbK5QeOX06SFgppVlnf0xbORZE
Xfm5KekcctdvQMWnn197T7QWnZhucyYFEuNkckrwx9YfRkchMdmdMN+4JdLd4ReF
9vESdcVaK8Sr9SFenHZyCCFPd+biQDtSjJxYQk8Y+jgB9JxG1Sm/uyiYNY++ueEd
8JowVjr0SFQ0PnENObIypTUzaY0Z+0WGBt+5JZQq9Hvxir2RtdU2kmJ0PY7UnNhm
2WZh6Vqhsjyztr0fSyqaR3COtF9GPaXF9oC62xaYMqN6UCpVSRZUqwjIO01lC6Y5
FVPp/rfZ7u1QcBwHuAc3/vbwVYUXKfmLgbiBkjXVTt3mR/cntx3CEgbyLAs2D2mL
zkPVnRf0u56Q6akbpBUTB8gHomCTJ+7WJZQgpXwgplM1uuqaD4EdblZ0v6wBtn0q
YaO/EN3igT6xgCV4vZoQt7UjKJvMEE8he1+3AYjUcu7/YTKtI5iK9qk8iH8BXJUD
Hu9nItrUz06Q4mtdhOtwOCemYJwqrK8mbxs/5ZmtZZfGWP2BX+xlALV0UGEw9xuf
8iUi+tup6FYTLnAEqt1TkSW21T+Qn/GoDlUMeBqXRi0QpMxG+/Kqe+ORr6Y6aGuu
5XMTVDC5MXr20Fp1yNMVJitB0PuAXcU+eq+oDaJgcLjNXXKbvMwBktuz7opkIduG
XX1r4PclPRA4nWE6+kuvX0baFz6qJLN0i7aQD88L2Weryrle8sq4o7p8lO8/9HQ6
10Fcqm/m7Z5ul5cooe7+fEzX7PcXJJ0owDY1XMW0c3t/+6LAjgCKX6vtb6vCY2qY
Ox03yi5SN8ynrnJ0D1ZbrL4y9l61fGtmF4PAZQCdfKnLssBdTv+RoRRerc7aO6pT
dcvzrtMKWdeOQCNuuAg3yyZDQpjx19arkg4KORfvcYZq6CUHzIVcuQONs0euz/id
cczUZ5G3WrRMmGi5vNWrBYhheCpsc343FB80Dyh+flSne12sWM1PlWh3U4/gX8ah
eKB+3UQbuRx64kWHOZgPq9wd8ZgKTfsDQE5/53svRogxL06Nxid3N2RVl16vARzV
E1o+XKH7GhPDrmE3zv3Lw3e3bVPRPKhXslI3paR1ezAa5bvXuol3qijtr5PWV4Lq
8AxP5OFsKucEMkvxYuKbiE3QDh3vwzOCFbyR6AZdBUZxuyonhIKIMsHzckiVOhtZ
CJvljnUouRwCWM7IOxk1AACQEI6DpGkPaIu4/qqgQzzPF7A0b0VOLCCik/RX++VF
Wimnc0vG+eZbXVpsRQummZzhFS7Szg18fw3jBRYq5YC97ShWDPTnT5rSGEMJn9Uh
kOITnAb40HGkjBsdUWtpJPjf4ITufTwEtMmYIprzs81ABQqqJaGEutW8hbdCLgWa
vwnNqD/f5V/nDdHn+IOj7bXqgIsLJApp12qtJ505cHV97q3W5a0y7QTkSqDaaQMv
5W18lpBFh8GDRUoz5IMU+80mr6YPELLT48v1klHLRfSo09Bx6GerVZr1/tSjkAR1
py8FuAXC8VjCiiJA4jIJaePpBfoJZGcbNPH/srOoL4m17b+DPcGxZZ6CUMAqcJ17
7lUHwwSuhcYbkklnC9ZByPbVKJAn7ktf58rVxdjx/k++GwNtViYx/r9Kf6VRnbHr
hYJnlaI2cMZh/qcIFF+bw0NRlCLbBs3biJjuW3IvOZHmnO1lZtyS42eAGIJOYFe3
xgmAGzJDma99p/KhWaJD591HNPSDwIma6coRsBgt88zgmOnNcvxPNQvN5USu2wWT
Vzh1oe8ucAXrSmdBQ/iXIegr4BtegRsmNsMa7UXxdcnnTR624K8Qa7QsAPHz13yh
KyKAu5wHJhPUM9XLern1EuN0rYmdaid8g+a/+pshCbzGp/9q1IKVyQDclReDPG38
7VgpF5Y3lrWX86whykeKaJJAFqwo/mPwfKyHuXx9dm98H5z8M9gFXj5LOTKZ61mm
Zgv3LJl08EmGvc4SU2qi9z+6Y56Mt2ayRyb2+tGcNQRR9KWvCS9Fl+gT+6mntaUZ
rJnFWtCE+nIANQDGGdM3mcVQql3dgCxzBqdyDM7m+TPaLiCs80KPzi8Citf4T/6U
Rg5qHuJH7ZQFxDX9DrHucYokYArKOr2NZCxDmDq75wDqjD2OPPUUfo7CyAqBOCZs
BHCVE9k1DH/8QK02JtWu4ZDAiNkmeJwr8eAOB/3LhhdkbYEQnvhJT0mqwu5etbjC
gZPC7Le2kuNh2LE4wWkZpt8ZDWveQcRvO76EQY/uyqUIfTP6nZ8pXZ+2Fhmtss9c
6e2Tk2wiEuaxuqLXhqVY5XZv3WPrId77MbhOBiPKtm/PKmYRqOJxDc0jhKCr5leu
MPuFzBHXNbZqm57xc+V/vFBa0Fq5U+A6pjkzqwUhnRN1jV+5HJHfZ9PZuLxHmIzu
mhtWEU70wOvOXvvUH5yy1TjzV/RSAZ8lZxyXTdHihLXBsm/kc+Ujbk1uDlF3uKhO
xpdaZRT8IGpls0CySETtKiOkZDUIrU1PBtLMsxKSJvYfM6sHj40k78BJ3Ks4q9M2
8fANJBqnA2kHmJKc3ycfi1VPqGnqtW5ccppZNmhb3kY26UbW9Lfb3kJP3tUjFWFH
XK0zm0ddCavCKmzcEGHTIQstkjr1sCBmFuPqp7whbCxgwixSDo3T/DvoMLJylsyr
/E/r5Pt8o0EuZTWGkkmIN53vMBcoAtmuhvm7tILQXBmSz/bGShiaNppLGuS0fybp
xfgBA93GidcHNxQDF2MgOsZUxjJ/BrKrnemScbnLve8abrTut2L1G9Yf1Q9ZP/gU
ZpKVFwPuYpXJFJb4j38L9amEdRLmeG6ZyzVY+ey/MNwBiSlykIJMTI5E9QKmbMRg
e25DtFHFKl6BU6Da7GSnTXuRRD1QLI9x/CKZA/OAFOuH3A62eKnxmENFFjS+JRzy
5pFMxtX9IzS3h9Fu3xhEzLUibDWh8NjCXnkXg5y9CUQKDrcUjR9/mILxuLolQ61v
dIo+8LL+XR5/qyuwxhVnoEGGjGwZSFQRxophCnQErQmRvYKTFc891/JG6Xh6H7N4
6nM5ydXJ0xna6J5Nb3bM0xUplwwFzPkQWO8dGfR6zJsEz5iZvwwjx7GjJkBUeTrJ
oHyitqyNMmYedy9OCFJoLZ3AF28udqAi+apUEQsbOb/uI23S2Ksngv9TrmgWsMdj
4AFXniuuEC9GP80Ten5V9aHSEAXXjsZfy55hNjgkYvTXUQpTbbEueP5ZYH9Baola
wINRqfofRR+QRxNwPn7RQJpRXPTisFUUBDcTWMoiX2GYwnfSBXEMzdGGbuMDhNXM
mlyY5DA8hv8t9LDMR3QdCUcTY4JpQnh7I/R4ur3bRcd2+SwZU99yrPRee+yKOjmA
RqNDYvQCzMnE0uUKHYabH+SeaSikURLMo+OU73Ssb0UiGd8fYxRovTzeMcHCWjPb
x+o1NUAkIOiN7u9CBsCf6Z7y/MEfAeLMA3fX1zTeQlHIkRKQOFE6vrmWg6mcFEX/
12pskEhW9Y+sKFNkSdqbv2syQI3LZO6Zn4AFjk7xnoJSim5pXfp10+0tQ1EmtxK9
y6KCtbJOvben6eWBdbu0t3fhbmpgfUHO9wPV/t+WdcJsDisCWIcn8udamgbUuHKR
6PW/17SWOGBXv7EmTRS3v8ZiIUZUN4f/AIlm/PPYljPfoBhxSz6Ml9WNGOvgEIPB
4Ot/sRezIaFjiIg4tgEBrbz7Zk55/HUwm0iDYmFPKC8Jayjs8mFCH5gxVSPJXncb
0Pfsbw5YGNHpMGfZ5X9xaUXZQ/K7WEhUKBbuUcofmCd+KeCLFn3FpX5eX2KE1Epj
bn3HKefBgOJOtxtwuEhweVE9Q7hqMgo8B2QVJ/jtQu1xmERZJwmFHK+Q0tzIKgNu
K9QkDZVKEvwX2050RMOXNVECowWnXt+S4sU17QGNk8VQgmEcJ3ZjybgnUPvZQEoi
a3af0hJNjk640aSYTJ2bsfOw+TSk1obYnho6y9sJHkLN+91sY8hWvQ4sygx4ck0R
jxfRoZHcwBSiHjsQbx1oCs7dG/Osqg48Jpq6rLPBnxtRRSm2bfTDCuE5i+Y3Yil+
r7YD3LVnoaW+QL/OgbJP/wf1jDUMxC3eYFZUxtYNASqxcAgl5dwTde9sFcJiuscc
PTW4sbv+D2S7pKA6GVRQ5vQrz7WaSHAV7gWG3CG9PNxo7mAp7koNfL3qRMFpyAKz
9xjhAjnzz6EtF2SUUShdNvcIhh46mQcvemZbxHPZGyX92vPcXm9aCz5NNKWu5KAX
h9sjRFkF1sL7Q9MawsA+9ommuAD2u24vclCrSdCetCUxjUYfvE79mQk1rHG7x7eW
VlkLp65deHrBCN5Ct1CkYqHBZm0hy0ROCMv86PhRYtf3fTMUDtcHYB9oSBXsov94
vdXKZGEWjkiS0ldb4pqsiba65ovD3lI0QiATl1gYRBdsAkWI+FK3iwYWA//SwSso
W7BLTtZdJtN9g6zfKR5OXf2QU1IKf+yJFZlQlE/72f2LEsNB9AgDar4Coey50TPP
/Fft1qq1kWJ8miL9wgSklKUN3qJzkP8LC7QLNUXstiNFTNijRguQJYSp95JRF162
ivs97F5TPxVNEMfKKgRiTmfXP08FrfMh7TcB726IvM47a/bAkAKQtXdv3o5OMv5j
+wLfC+/qxmQuOC8REi+h6/IMezKY7+fEC1EZ9ezvSPO8cbQpWvenaeuEG4WfiUrO
s0K9nJRM8WEwiepJYcWGdMNOw/hFD6N/AtVzudVLFTjBiU1Nlz55pjUJHePZkUSM
qyjIsWBbocHo7jz1fLemnFxWiNyD+5P9z52wB1YPWL9kMVFJ9YVktz7ASqZioc1n
+XLquB/wSKZtHCxq2yVwabjnZSBNZoYHUGUDkLF0sQhkk3lGEZS6qYg1V5f08fvQ
I0jgte71QjeIWCuxQJb/e0ZRHVcek6ZtaH4Wd4NPLLkkzDIJKT/hZu/ovf9YmABP
Udj2vg3o5LJy4LM4/xpupfwpk2dKmFkuYbb8wZUJ6swfwpZm48CIqRydEXxhvl5g
9+DmR6nVOKgYlX5smvdCseMCNFUbl8LeVz/Q3753g1qjlQHY8KRvuNcyvHsZTie/
Jy55Gv5jKlIr19prZIfvlKX/qRZ9VU3Ag71GbFpOjK5UHn60pj+n1MN3khSkd+Ip
TMJoNoWsQwqEUqunT2Qv+gW847nhNMXgvuewMNn7HTVikDT5T8KdhWAhjeZWpWGs
kO1UFmPwpElQ+PuJjQe6mnW/OLsIoE3HUZuSfIkx9OG9jry4Zx/sSOJPKTsKfApC
e318wh3wKPKbW1hsXGNfOcd5eBiRR5rqPhgihuFpz4jKAgAR3P3BirUHNoTpUZJx
uIu9TbvJtQ+oQRdQ6WlIRE8emlAHN1Ikv97TlH3TfzL+IN8HBc9GF2hnVbFEOAbi
MMP4TqvFoi5mlQooxwQy81nKUv6F9rWh8y6kak1bZjzmFpH6Gg/hxenwZxp17fI3
cKeK0v9vv1hsbv4QfGRgoMd/Er0R0J7gOrFSdnpJZPPwGgtOfoNMihb0XIVtSHYP
Zyh2HYTga9Pvz7yCtYIx1xBrSGlZDCJ8KEPviQRC4LR9NxyZ1RvrYX0SOQfd6BVB
EH149FF/YNsNhmLUrcZ8cSNXnOCv+R8UF1LkhPuhCOUgqH6zCeWXWYctLHS7oOfZ
3ngs6MGPDpLUmZWGd+WZSNVkp3qkRzaPAlN4z3AffeVUi9d+ssJrSJiX7GRwB9SW
qtcGSY8P8wqq9JHJqjrDlubv5AD2s7LOOXNbGNmwVZuIiyTC5yE0RJM55UgyvmZB
nGzcoRcNFzHMBYOiGXEuqeSj22h/yJpEE3uPanVp5kmvukMPfbrBTYfuxUZHikaF
jX7lbo7qkkTkMrBeD15YH1DslAMCFJs6rcd7kL2xDTH0EJhPhfDlUazp0ODplCbz
ZEkArI5O60iTWGa31Ko5ZDZj5/VOQQZev+YRZOH9/M9PQNMQfq8QbjRINbAwha5P
LXwhK5cfCbhu3DHwfxr7VSF4JIsehkDYciXygWcAOr3OMk3gOBbpVt+uVZO9Crd/
RPTyg7TST6k5IeW6Y4NORVwoBSFd4gsi8gtFnc1q62trozxWNJ8FPMRdNQLoQaKv
DdcnJl1joRXxLrrhr+VLSORYPQk6WIsDr8LA35edPaVPZ5OVxmzljX67uHYkEXEz
W6fwEbkA11QRFoX/A2S0kYuzmzsTw1dAPC6La8hrkXyPx0Tx7UwwHI8MchYK3doP
JPOJ+IGqHqk1Q04kztPzKhUhoxcwbShF/M5wRyfQWXABw+Q8aXqWBa7qsxNj971D
Romwxp1B6kk1k3tUUqukFE+9ELPQB5rNF8OgVigAsACGCb2q8qEQBUao8EN3/wsc
w1m5veM3V+wtfzblG+fhYz2E6muKzfb8qCAB4FwPCbok8gn4/7kX3AweIFXxWeF0
JK7YekVp9nmbZI6eicEBxWZEviJ/RcesitQamiOFqau3pvokF12LdU1rOORyPtRz
GuHBVoBCx2uPtllTnpZYc7LEoAjj3KzD+tOf1n5fbjvY7Zkr3ncc6DS3D8p61Bwq
L0JW11TvlNgb0VwYSx/JX3H8fYbZ606HWZDOTX5/Hq75ELZE4RsV3c407C/rtJUJ
3Ykl0YXczKn65XQbiJkIZRJnYRWhKpDj5j+LgmX+idSEQKNZGXwbbSUJY6glPACL
PkbsQOQXNonzgg+5j+cvLGVgpMWU6F33Rr1mgirDE339VYUehO8XCwcWc/hELfZH
0VHJDjTS7jr8nHk7WqEmbVBb9l8W4A3ou/iQpDkZ97/RTTUVnhG4VktFtGAAFVzl
uP1QTrPL9mDl1HfZYJvYszO42boLuT6ghx3ZVEypf7lrc2DzYf1PzR9uH9A9CBSZ
CIkP0PiO2L69ufmYNxeUp8QNTtiC5aFFMLKsfqpWYFiALleAorzbjbZkWOL3ye+W
UHTLtFT21hBosYOa2ePC5/JXe0GedSP1aEthL48sXJ8v9RXwioGYmmKTQas7unkN
Bzu+zeWPP3M2L8jEgLZkHpoCKfBfEAttUPDmSiZhZSQ9x8ipctXV2mfvl7J7/+BW
sF1CSEgsDikbylZtwnv2llsFYVm8lKiPX3dFC9EimQPi+A39BfqWyw4HlSgnZrZy
1ca1htMFiXetdNhKKBsaDt7qAB4egtjrpJoo3PUTPhO2TXLqpJ9dBRZ2vynqBc0E
cqsBU9dJ9IFz2NVE7uOw4L+gdwFqCTCadn1dX938UQLgF7iA22LoMXKIZRc8dWfD
5mP0bS0IPEsXlEmVL0lB3JHnFxvTK7YeJA7ob1mnJRIufn1Dng8Aja1Vr2Xkk/gg
/moWazOj7W8ddA8hUfkx+1DfYBTS3qIomxO/rlZa5ZsoDpODK+W1K/3tAtVJoxpn
VEzW9j6uYRKPAYm8gGWGnUFB7Ni9FmVDxYY4Ax47xPYzt4UCIBo9ulr8nskgf0BO
/1RUKyrZqtS/ssHp6j2snKo2MdiqG6XpeYO7p8cT+GjQdbDGDE3++MRCeHa40ot5
ryq496pJ4tJS8EnJFIvQfXCrhC7z38nB0UlRRTTqi8TDJs6PqiIKw+t6emcT30vz
QZKaZm7bITeAWEhHdT7JTsmYEVlAlXK4W7KlBcq5tSW6FT/+VWnKTYGE1qfOEuIk
yqZtyXtO0cHeAsOOyr6rQO4TsBFIACLOpL6e9CPGc6M7Zeyr+h1nUSFlRrnUkz/8
hdxmcGXejKARJs9H/C8INBYAHNY90iPnB+7ukhMmnL0/MGVC4yj57f+uitVSexbA
LW8NwqRDmjswCZEoy1DCriH6mHt7Unhk96faFdD7ma2QEwhd0CBg9bNyAKT4mmkl
dCl7X37CjXORQw8qXRmlEWDj1h/iyyLNt1ybC6fGd3qoM9lhtBmY/3q120tMayHU
5X6988FJRPm++v6zKMFXpqQvTIQFj/ebrGpF06WlpeSRBeF2q0BdyA8Akg0vJdiF
IT7lAq0kByQxXWv8skDnhxUH2mV4QqgiBL75v0KhRzmH2o0ZSfNdS3cGMxAlOZeN
US+058Pgl7/MrOpx5zBadBYdEa3SuYE8jM2XqcC+UvggKO5eXDZA3Yk033NjaXTJ
RIXULM9qLF0QEeuJen5JSNZbuRKCJ7AESg9SKADiBp0Q0JclMVE+TTJNcNXb4Y3W
y9HM9F1/wdyiCA6zgR+jSRR1kHKhWJjwb4iFRrXvxX+J38jLdo/JgLEZ4Rn8704v
N++PSla+DUhcG4Rnu3NNoUAjWkpqvYmrRWk4XK4CHoUf562i57vJXtLUALklTC8O
oqeuGGD5ol7QUeBphdqaXtIFvSmVDRDkOyJu2jGt9HNq68fWg5NSe5j1fuNpwKjK
oUWGk+P5efEzpjWd388Ct6qOM+4S62G7I/5DzacbXJwE9nVmcmVur4ysoOKBrxp5
2H9GY0uAlKUQ+Hbu4RwZuyRSCWL3ibvfWMYaS8JnotlgXH4CHbwbkMnY7FJbfiyd
xQvRNgWlTwtqwRaVmvK+52Ds2VJoJU5x+0CZR64wP1HPNjvGp0vi5/wYA9nVYTcP
MKyfeM6GhuP2DXDbM7dAnQnGGsioMx8mfFWy9WHpOHHQyJfKLw1vsl92/8Xfs5a5
H2Z+jMNrwiQU5NqOBf4OEckpctUmafmFEqeBl2SodlL8Rwx51Q7iGPb41WHZOdqy
fEkBa3vE+TszugyhegKIVZRojEETxdrmjJ2QEF4v3IDDnuUhmdKrS2DOCxvlGJA0
WQXufKrPU785pnM8g4M3ZrhmDDzYQxodmSWiTVNTMgymGD2/CIVIL7XwvzmD4UZm
cS7+2VEAT0zexyjYBxPZaGz4MjWSSHgIx5Ee6v8Ao+Xk1qhGYwVAA5Mg3Nmo9a/x
oSlF7J8e4SmQu8oRBzBk5JE2+GQv6Le3cn0O1nMmm8SP4KnCgy6GUk5wymIh+NyW
4UDT7y4rKpJn1pA3IG5m3UN2jPHKyp6xYFpGM51Kekc8+LWXbbhLRW0YmbslQ0Vh
KO2T5gGxNky/E5zEtacGss9DyUwtZEajwSIPmPQF3nVn8QLhYNuom/NRyo5P5gkh
3CHpqyYKUQPre4/Y2v0K8OrVN083ca/SdCctgvpGOYV4GKgNp4nZfmiWzUJ0YnDr
+UVb1cWeFImNH8m0boSfEu8ep8+kz2TPeYa0OOkLv4AdMMYWMBmy9EQRJivG7g0G
yYNDfH5xmCMYAEzsucYwa7K8fPIVOo2YspImRVTbSPfR2FPPh6wQuDaRTTRCNRJp
7CTm7uAFEAFR+WQ7cBPrMrTciIdVnI42grdTA3b2ohI+5PIhUc0XDDhGko4lF6Fa
CW0Sn4etJEGagXuRyNzNgh4rehPrOzTR3dsEkKYV0BzhIRpDpyXrKrVHYv0ZGR8p
OgHnFk1ImYAa50mby0UBAtTyciSfQZF0rfIsxbEZCQ3LPkG36vwDb1saytglZJy3
lQCwXA94p0odhIWafGB+IkQr5++SDXD4/prxzqlUv6yuj7Ad2g1rxelv/F9j1YS5
aLbuC0EsTGlWc8Ik6QoXzTUDh9tK+LXRiigRVuTSIsaGuWUoUwrQMNhnIdD2Ghmh
yoswkvtdnu+TbKMoL1BglvdXYofsNztWPiM5NWdrgcLxJpREYRJVECGZ7fzgZveA
lDZcl8wN/mlz9YH9SY6UZqgAHJx4k0Frpg00USY/yu4KmwVtX+o0XMowF+YgEk0m
ZGAydz+PJoSU9FXrRrR5wf9NWR9G3J4YNU9j86WLDaEXjBVacj1EEiApll3ErLUM
VIChxfHNpAjWKZ0hK+h2C2NyXwsttRiQpHnbVUZ7nO8WaRWJlpUkOXUVtpMEekLP
GgM6euz1iQyqX2I9UUN3N3cKm95GFr0lIqbnDHXkEHEgjhbRw3ucAfsBMliId9EI
fZ+9I1/V6z/yzCcdQgNXClFRm9utXCFbMW8jdDSyV03cnkO1ypb/SHbm4147hkAQ
dwp7QDZqVPfcRQLoF2vLwqkKUQmPRFXXD3de8VCvrC6W5D4/U+fiGyZMKfOziTGX
E0DpBTUKA+x78D7hqoLNJF9JfBVbXXugxikiJpR/6HDznzTFAMKPXnlbi74NefqZ
K/I33/2RC4BWpws2g0yb/TR/OIp1jXufUumFwfz+55lVs6iTL4KuQAFq6BpUjLCS
qMkpZTPuQicYZF+xFJK1yuSeQ8ll0DGWDdkJoCuy4C3OaHIGKWNZ8dCC0IqNdc4v
XkJtOzB7dSW0SnQWNFHGy/2wulIrKwOftcW4Gl2lVI++ufMj55i0HPf096HpLBTh
SXYOK7+Ge6a9CFpgQzOFDngFSVEi6FWaJGJkw+xrmaSnLKBmxxnFhGLBGVS1pWbG
/ZV49mmK0pRwIOykBLvWNUJYpThWm5tTooQP13WWVIzK1uYmYgZ3dnu4HeporPFi
Ac1QEZSIlAQImPsug9yv8j2IGk4q8H5SH4zx/HghUV+NUyP5hZOtuhFZfRfjaTuw
qGHR1dotuHismTNGteRyLI9e2cr2lRfaIwSyifcFp2oa5IzzKUKtKQMLN45lS9Fu
k6Nn/mPhg7RNtHPwH/k+VEeJX3TQyPCKozaiWEW3VqdHLVhThPlx2DrI1ThMPhOj
juA6PSpSeDsM3XN/Z+unk1mmVNvQ/DNkcBdSaOKszKqx9SYY2Qg/DXXtaziZgqBJ
bwfxnlMtsjjHrBAzal5OxbjoXQsWFzkDRR5lI2f2nvNcW1W+Gft5H+KzI0zq9mbf
x9JZe7PJT0b7GQGO/nAvWO/KPJcDoNKUsDy0TgxSJqgE2qTA4W8K+T1DDXjlKaS+
LKusdxxBqU//rlh9I/UWbnWbyb488Y9CU9CjuAH5rmVsBRAubpDYXnduWEMrlpwD
E8mdRRWoGiDTOd+69EU/SnURNe197+EbqRxtonTv7vVqmKtFzuFjR6ATltN/J7Wm
tEEugAmbooHc7Dc9Vf5EnDyONZs0uiS2pKQmaLVf3GOQSXwXq+2yuKBObFawas0m
f47vYIRTauRUBIUk0lL10oEzRkzXQx9QBIPrp5rPerLHBaIq5RnsxEPRqquCuwwl
YTZ+ysiArXRg1IGVS5aRalBWmuQdAyiuMtHIeAJypDgDTmLfziFI/KlZY17IrypJ
Ql7mZOMODqmGpZXEpPY5C9/kGJWcQk/9z+YBQCheOoUomdCM5dz8DYyZw7xyqwb9
Axi186WDieLrCwfXxT0mIoft9R3GebzDO5mr57s+D4O95yU3GDWYJI7tdIdvS2hN
snOkvEN/9bR8SpIShw32Bn95fdE516zNc6RjdOrsIiKNdtXzpmowS9DA6YejIrLQ
cYzjNtr/kgZLtzAAqrn9dEvXW4HvITC4QmFCo8aygUeIpUpTeDN2nw4Q6ZS1eIX2
sdt8jeLS6qlNajb//YLgo2/KX/RlzBYHvn/ah8lfTmv3+G3WA3KvOHY1H9Nq7NEN
/e4oSIzGnTepgZP8LIbhLf/3Ak9aUQEWA+1SHPbkcDIulKy93djvkc5WQjJ8wBzV
cIH/j7XIPmUaxCJGX9qVsoSTl4ih8mCuomYg/yulA4Q7IfgAo38rGqF5syYvgUOW
FyQ84ZJX/UlnCy5ykpBNLzcnlERRQM59xPpE3vZv+aXOLh/RrvUMCe3/3I83n4PG
gEt1XcR7ux9pxXBdCTPTGrwS0vMojN1MHNVvlQZA5G3JnPixHH0f8d3tY7t/bYrb
00Yeqvbxe+LffU6XbjIEyqS5TRUvFyzulzADMEiXARngxd4pDCwAVDrdd454uUvF
aZaAA/WazREZehy81YNDeiyVgssen+B4LckDY6BncJsP853wJh47taGMVhnpTm/L
zmYog5nb7UsehD4CawGEbuxvpuIGwOHL+BMRx4zPXHfyM7rMYbh2OeGIw1C7KZB+
ty3kftPQxZ2t6Pc4GfG3QnXNX50TBWQKtIjMddiVdesYVGIwehKEhOdNGVV6lzzC
NY34DdZLoYS2qsYrVMBHJ3bmWzfjdq+UX3haPsTvXk9wMnqHSXGWE90r5KhXHUQG
f2063e9eEEmUNA6e/BDEUcfQIJRFk13tcgF6iaftngs8cdT0pHgBJ6NelKq+jyiI
Q5/IsYVGYQiI712ks6xDcVXPOQDS/Hfv3EbNaQf69GVPvIL7eBTSrUxCtjMdp3XT
R8riSVRq7UpWPSoPtOX5G1yDxZ3SpwZglDViRbl3Zf4RN0OQKrc3cdOY0rodWqax
PdRAe9g0/pq94j7IvW6WDWn7hMXTIsI5LsQmwqL7omnqr/BQuDUEf7sGVtfpaYFW
ME6UpobrraYck7ulF+/6Gpx4+lD1VaieHu80yDYW2zQaJI1kHABesL8bPljydj88
bH+p0C7lndunAOl4KH/4ePCVA0MZw2/4dmAMIidbmj4d0h1WZXvXLFoluRI+lSdJ
zD4b5pZtl7Y67NSVgsn1ib92TF+MKpY3bGX20VLwQ9NWaCn+Phk8Agqpxf+Gn+dN
vx3D2UGBsico1QeqB2v5EjDEh9rq0VGgo7gurR+HfjR+/wTEVNvyBM7Mxh5xmlTv
ardKkwMHO2MiU6Ur1xlioiaJm2lbEayDFvhSCQnvNMiOOML//PscfDgDx5P1ha14
y+Q0iqkoijnHvf78Z/bu0bb2sf95JxwsbdyayuRTGLOLgO01d2ekLS5O8Jbi0KvM
G1vu+0E0vJJX6i+epgIY3Bn7oCm/vPw+V+nM5f/dZdUtwHF8ZzloChknruaC++s0
Ew0xSM2q2KRBdwPXf+FsDekQcUs/4BrtetFw3CLtntKVDBVoisyldMZe4/ZaTIiP
eA0CJWG04/Py9xZKrbrm0VkdZ6e8PhmVxNt5tfK2CoZ3h60fA8uN0cpXqVAraHzG
o8jiaOi07tn1W/zx9LYRu62HQYAp/AUXCzCZyY/9FKV+x8vFZmgZnCsvdYcZDUvQ
Ie6CBQ7zpAPddQlwS+rgkoqXDXl7qTZHrChSIIeRe6lu0+V12OFWUrQVnbDpo2vk
9ZNYtFFPrMEyYO53pQuX8vi/kyCdlmWU/ZiA/RvT7WUkCvgvo30cJE4qzmSVnhmY
jlBgm+WEqi0+KNnhWKz3/WbYhvxxHGttzfBe/ZsswfccIlGr+tbtgBqKi1v1GVxA
+3aBOtyVTaziAn+j2A5gmwJBeEJwWo5MbBdvRRBbuGHTrZR6+gd2eYCYlwub+sfu
+rqjiICaZCeLUrhds9hkBvBzM0EgmAQJdrDleSF65mM9kO42eWZmUQxhG8OPEfOa
vJMlFWq/3PAqQSE24lryzWfR7YYlSD3Q+5ufJCtYZ5pUHg3o0+kxBF9E5Pzwkrda
+TO18rn7ZZav/leuQimpUhthGlmRyk/ZNL7Gv7/1aW4P6ROp0/Xp8innYg1ywLbU
+6ne6LSgCsoq51mT9QZkZgQv5P2rEOWsmzyp6+6TaYUzGY2M5wYy1Pu5yK+GApAK
JYLtcgoj6lcsAOzoIqp4PTii1Wng8961P+pp3oW3C9MiWJJPAsVIui0HVe385/Sh
eC/aREA+UQKAgE18GrrVWQmeWhFLEugXxlZPNzSfXMKl6PDyQsRAOgyqe0gf+GoB
T5H3hBcHbVknfyLoU3Axbnx7061bXitEdO9QomJytUn2PlYqc7Otb1T1awucQEyU
l718OL9jtoOBhMN73XeDw57kdAeFIFFM2CnMwoZm2Y3iTZbNq+bBSyEaqabKRB6K
kmd1jG/kjkJqPkpa7OiQKFeSbw+rNRB6kPU5sQGzsz0opStL0k4Q+3JzOjOJyPAf
TtrioLr6YCgaWJG/XcTW7sJo7sizo4M+uujwd8IsmtJpdqXRNGl99USIq674io3n
LYLpLHhpTPUKBWH7aen+cm/VeOLQHMCVbLcI4IBjG7F/Umir0Nqu3ePyBL+cxUqY
MCyPH+pCwpQNzSHCR1HCaOEZejFjDabdytLKbiNpQs5kOjnj4DAyZQrJU+3Nov+X
AwmLM5ronXIcI/tMOBw2lVKq4Jmnjmpoi65gYBc4y8yqjLJJyWcRqt7BG3q1lqnL
hqeMsqLpcg7icYfSCt49+fiKyh6Ob1pegu2r4YVWZxKwkDaYMWs/ekORKWpj8gZ1
B2a6CHF7bahNvpk2fwMYa1Ac+OTVzxe7iAhq8P7Pv+H0qlJigW2jid7IWerXs+hC
nH+s5itXQsGDJppJDxp4nR6Yz44SYaZNYEK/YqexkNaYzW8zOgcgXyLAT/lfajl8
AQXtzGvB/jvoXIOI/kWoi6oWMA4U97OG3K2gL0dQc5E6sUp3/UBID4s5H8N8SVoB
IL73b5Y+7iglnuOi1xKM+TYj+vugx2pkg3BcDjHi+b/SZyX1nxp6JrxCOOYLFHZT
g3UYN+Q8Tv3wIkbnmCNuYAs2d26KIS9N/EZhfQHhPxb8+3WpyQtX/LhGLWRvqYGJ
KToVY8bDYTdgPwfpGZCw/7OZMePNBuKsM/DZJY508Cm19GlipB99oKG/QKus5kQV
kvsct1aeCDmBggENUY/rOR7exxvVA2ejMGwGyEgP/BQrjkDwtmQaLAzr6fyK2hap
iqn10YJcAfEA7lHswdQ00PSKlz9yedO1UvrGSrHE/KEJ0U+kn2fljn96vzuBhxMF
trAMWPFpan9X9UgO2QIdEZzXeE+BAL3UEzmocJkaBG5/wzo0GNUZ3OLYkymieg2J
U7L+sSEoGACXVR+oSJ63GwD3WxdAfFj2poPhf9gHPQQXpdXTZmEGgwj5i+V0rs5C
7Aq+9RHK4SgTKUuB4zQY/FDwkzRPWRHY7nR7KT2Yf/22B5HxJCWAgBDcV6CGxlup
HefHHtKFX6XWTX8/+vfSU2HHp1BLdat9EyYlvQCh9XhPsrAOV4cqLArUo4wZ7ffj
gqeXwNso8Mz6gKtMrMPwFZL2XzqZrkVfg02rhS11YyCLMNCcYplAZVquXOKkwojW
X3y0JjNKHmtatweNOYUJcL64C3ewQiPmKblDqHp4zy2RvOiC1K7cSW2JJYwaMPmP
wMi05vkfwR3DFSPHwN2vFeB47tblhkeIVlMPBVagP0f2HTabFH99bp0V0SBcMCCF
GXhVA3h+Qq2yEPQ5Ohxn9d73W964HpueO9G0LeOioEHjtqjkqt8y0dR1ojVbsgAb
9Jfzl075q9B6MNAR7b3Tnz3siKtv2bu/WrL9N9JZq96eDsgJ8ML0c1vti61uzA2o
SY/ptlJgnLeg3CZmE4XNOQJRtrrDdKVT7oBBTOhTW4MoX8turxkyck140IB24wGk
3WWm2vPtYse4bMBop2ykc4qZXbYylYfbjvd0l3BfzWycMXP28Woun5RW9L6F6l/W
TjTBvXXonGrl+RY9GkJSfgcTwVow5otT9qtxV+K6UI0USlP/kbkokdyKgWa/iHRV
TAQugj2TujiG2S3tyPIVsVyHaRdxQWphZHERMI5HrGFa+uMtdfirdlNOmKkzdkqD
fC7HIDKphf8m7V4q9DCunjTwNhVDvO8yHBF+NePcGe4tkUcgjYPHV17nPB2Gy26b
D+fcZROhMDhBiD+tVfN4qjw5v62x5Lqol9Hyk/w6RRHU3ZWBB4W/NslruuZYEfX8
RbKoixKzi4NaajPb1D1fJNieWkm2CAl41RD7aqZIPh1C0xUedhOLpBAluFSEBXxw
O+pCUCItReuSTWKyBNgwP5QJn2qSQp+hw/UStc0GNuLfsBuPsK2bed27bNEYDLRo
aBwq4km9o/pIhcdyVbORrG2Fn0U4qPXUvsk9qGUMPRK2IHnM0AYYecxeugL7p4Gg
1nbokntx5QE/LbOOTHqeTLRh4TKraHH4L0yaHmiOqe4k+8f495XOYAFgZvLo2ohr
PB70jlJNm0gbMaNRHEG6TT+uf2yRaxLJh/M6kCo95pJ29JWZgDnFyHBQTQ/jXhSN
H2sNGPPxZ5zbaOLLOvfFU7pDO2grWpkWMC9ahGgEaaLozd6/U1vXx03cguetRUJW
++uKNqNaoP2W0TPzztVoOsBpNtIyT7GJQwPrDUMjxufkdJZPeOH1Em7l7m8CDRIs
X5QHQTVtZuIFBNtCsiuMtAaPTVokHMGIYFYKxB5mz7HYqyAqUQBreegTc87Hv+0q
ktLaRYQdv1SJ8SEoRiJmINoHjdPGJTSqmTqJUMYUBK8O80D05krMKf6HXWosicda
C7ZxiCNZ+6hLYPFQXnxYXr+bDc2HzrgxgwnqXYzxKrnGo+sDqz689DpLRXZF2S/N
vGPn3kr1+Qd7FqbKkMVIe8brHCBiAVIT/M9lHO8itaQbVrd+WAYWJRhMIERb2uMI
DWUQDCnu0zF2EpHTBeY26XVfi3abiVJYanpRw9C8qMbnqO9UJuBdZrhshvk8goEZ
OkbRHPA3tJjRplcTlsDnbsy8GmuzUm4f7lcaEL8wINMvRauI/Aq0MqvRnQukkmVp
aUrDBMpr8uPiZ6e5UXyeGPLZOhpXZ1JM3Qoalm58KKBzRkuS4RBiOUZsTN2LUrDs
+gTs+NhqJ0NoD8E6uiNpc7NNKb6/DKJ1DFFPVWMaGdzywq3teq4//nGD+HZb/VG9
ylJrS5EHDX7MAtfL0hw5o9viHAB8wYjMQwHPOyp/GUzGmHxLp4m6zPmIdIVgJIZz
y6c/oqHjo/Ikw0c63DJTjXBP3RsJZYwMtjgymsyVfbI+R1Rv63407szW+eolgNYy
ZIP7acy3Tjmgu1Jk/XSM/t/2ctj8CllGH4iTTsK3XZ0ScVwtE8RtiN85AEsNzajk
A6wuZISeZCXKmugmVeZKw1Bz3P01Y2hUbnuOUFgnACLO7OaLMfeREynAf4/mbbok
shuL1iOArPDYwLNQCXFissePmn3szdYlpQU0FrF3kyU8sJVq4etaRhgI5sLsZGtn
vrLDpagS82L3rk92LHTfsEpU5DW9mvzJx8PVNiovirdJPOHIOgovSQwJsBigqR1L
y4PhhG1maEpEWHQL8Am+i2hQHBQ9kzaMxmaboTKSYOsLIBULYn0FcV6mOhMCRPJM
pNiqVdqSkjJpG3rLklXMNV/kuewwTdUQEz7fGzRKVBGEaqqz4C9TYdRUzKbUCSLy
zM/SK4UzsCKyzosVLam6irfX3WXwrOEuLyfBZBMjVfOPP20oNeG5HlJf5+E0K/c6
rSNz5Jq1ncv3ZPBgcLBwShe1hiijfVF0UHpmbJe4ZTdNgf22sg/jehauFY6pLhp6
wExPT4JgZhW0Sdt8KRcnAyoh3LdIxUMWge+qZC99wqHADhZhl9WR7CavT5B4bFD9
K4xfwUmUbD8keSU91WtHfivr7ZguPKhBpw+KoM73uwyQoejaTsfzJ2yd3CqdEioz
Xq0HGAZziBGadu9m29sNCx0Ps+MFyoGZFMDYEplbVHIN2cXqi+q/TzTF+rvnshYW
npDv2oX1hNMPW85rkFdw69ztd/vi8XQKLIIa6p3DtssTebzX8+T+2raTn4PMsf/c
6POj+EtLl5CEsW20zo48fgaWhihb56NRJ/fCwkCK0bWjtFynCbM/tbEf0vVU4H4x
X7KQpGeNBFw+Nw+e+VvuNac6SZfI0yiiz3QJlWE8cCLO5wY1MbGc36Sbhpcq/1hG
HLNwn9AN+PbFD2vLrvHvWYraiTP75RdbZhhsNxvZuYeojyUAEZj5magi+tFJfYLw
XB0ka4Hbqg18wwPkuFDaJauYkF7cKfZKYYk87xYoJO9xpcTzrc4Q9dfynC5yeea1
221Xq1XrKvy1hpEbxJpqGGETBsHdNB+3H8xcT7cOiFC6TF2GoFLDPFb7msEzwuax
hKFgkRG7UX8jhSCaOU6C10wJ8uW4QmmJfkOhOMNRStCmHGRCePS5peMlG7kzMdrJ
rIfB/KRuqKI3wInjtAedXg9pWGdmbTSh6l3yJG0K0oxZwZD5ueNyPMIYNgzQb7Pe
ZC6CM0tCidCdMOEeXoqx57QwPUFqfmtjjYaimSQX7jfMFoNlutL6S5ReT2vMmbTH
9drZWe9ZF6RuRWH5dLtML9YocF1Gj5r8FA/qVOIV4MeFtHdybYQMpZVzEyelsV7S
y7b0quH/zP5C+qB0gTAwaYv6z42EXK9rHlb1fNlfHqK4FNDECRyGlk/vQ40ta6eX
yx7nFh2u9HrfPQ3TQEvKbYOGtPgYLgg+tMOv2f8gPDkm7IQDkxJXvbnUcZUYmMOW
mTxb1iv1Hx2zkhVV2AfHU4hcj830kJY93KgNNdcxaQ0TlafJ8SXXTvMiRa3D6UZn
xibl+u+yIMWsFq8kIIcumzD9rZi87GmvDzIEYnm9sHboOWeOpUIg0Av9WqoRE+5O
hl/5IJ0HzsMOZlc7e43g7Qus3MvjmNTeJnCH8ZCmj9HDY/dVj/yIV7Ode2bJ2M+7
z9b9OKxeiTp5OODL3wdCq1q+IC9lEULyYY66XIrjatjwZWoKkIaLT470vIavTU8c
aF4gGkM+3lMAT7Cmw7Z1CqEUC6I/ruTbxurqe8BRaWhTHotvaosocBe+ZX0Zl+d7
d7TUXDXEgoo0HoaloGT69aw/MnS3wz1cE8zUTaXyMagowziMs+6cljtYmzpg2zZ6
LoNppj2x/vt51uWi/Iig/0jYwu5l8CD3M+NXHsXc3D/n95Zk3aQ9k/uRJAG24sI/
0J1VseCUzwo5uaxGSKz0fEF4OebST/Sd481CiEUuU+eakh+nPXZuyG52skXyTwsF
4TryZ+e8sqlGhbJv78rQNxWeTjheRkHk7HzPhsfr3sw65f619QaedkpDGtyn5Ama
fLlJmYmfk6cq9INQH+lBXFdpK81tBWJ39WYid5oHnEDUMEogSx2sgz7nmGbM3FVg
PVPmgAvx9rBx1R2+WwnCqgpjim4Hsc9zbuV481YnShjls34ptojui8nTi09joUKx
6vmfrbadwPgof3jts9TVZ2+OR4XNPDCK06aYTryFUX/hb9tgFmvGa1a24f3T+yQz
vBqxa9Y9xc7JxxdHlWTE54g4MH/ad3x/eEhzBPkIB19FJlQD3noIzUoCITIHLMvF
bFjEHi0HjFvB2R3gV8xO5nFwl4wBy8/HO+GKZFHSrTsL2/OOnVRdv3LcxG+bmccO
V6VKGsTYx+Q67lge6KYiQbtgSG18QzTcRbjQbEnnpIqH7SCyqnJo4ngpm4NI5HSI
QSlcF7uxa1YbL4Iam/9Ya6k6VV/xZIlFobz9CjoIZMtrZwU2wPAx4U0vZxhakkzm
+OQt/B3zTeb8skndJhcUP+WaxBKd7OdEjAnairSNGdDeCqQ8RmJ8PImL8SR4yGEB
fh3ZYJX3CFGctw0BYaMPtEa+JxFUbS9FEx2Wrkm4Rra+qv9e/Ce1bBYxZWqiwyVb
O4WraUqbqUKok0sDUEc2KeXWY4Oa7ezuJGIvUAfH5AxK0cEA8wlWOwBhANPNBXrt
ZImhrd2v5tqMSDzIkWzJpwhUg8fQjd86cJuom7gd7QJSe2TYAM9HwyF4ZweoJIfR
rcc3i6Hf/q68F0Fzj1XOyCI3cowprDyvoHxnhhbN/T0BCaq3tCKBWKni91pQSGjS
2V+lzVXvjf5Dlyt0sB82CtP2DjCQGr46tUx5f7pM7d20C4UxFnhPhaSVc8KDcyxP
x/igjoLdbPA3sJDNFuIKF5xbr4kAJEiusxZy1UocacgFhHzXZcEqVxFxlfpKfUY8
bHN1oSjJRhbkRhm99vuV1wDbBNyTkkvsicw2SwJCZHU=
`pragma protect end_protected
