-- alt_cv_gt_latopt_x2.vhd

-- Generated using ACDS version 13.1 162 at 2014.04.06.21:10:36

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alt_cv_gt_latopt_x2 is
	port (
		pll_powerdown           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           pll_powerdown.pll_powerdown
		tx_analogreset          : in  std_logic_vector(1 downto 0)   := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_digitalreset         : in  std_logic_vector(1 downto 0)   := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_serial_data          : out std_logic_vector(1 downto 0);                      --          tx_serial_data.tx_serial_data
		ext_pll_clk             : in  std_logic_vector(1 downto 0)   := (others => '0'); --             ext_pll_clk.ext_pll_clk
		rx_analogreset          : in  std_logic_vector(1 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(1 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(1 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_clkslip              : in  std_logic_vector(1 downto 0)   := (others => '0'); --              rx_clkslip.rx_clkslip
		rx_is_lockedtoref       : out std_logic_vector(1 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(1 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_seriallpbken         : in  std_logic_vector(1 downto 0)   := (others => '0'); --         rx_seriallpbken.rx_seriallpbken
		tx_std_coreclkin        : in  std_logic_vector(1 downto 0)   := (others => '0'); --        tx_std_coreclkin.tx_std_coreclkin
		rx_std_coreclkin        : in  std_logic_vector(1 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		tx_std_clkout           : out std_logic_vector(1 downto 0);                      --           tx_std_clkout.tx_std_clkout
		rx_std_clkout           : out std_logic_vector(1 downto 0);                      --           rx_std_clkout.rx_std_clkout
		tx_std_polinv           : in  std_logic_vector(1 downto 0)   := (others => '0'); --           tx_std_polinv.tx_std_polinv
		rx_std_polinv           : in  std_logic_vector(1 downto 0)   := (others => '0'); --           rx_std_polinv.rx_std_polinv
		tx_cal_busy             : out std_logic_vector(1 downto 0);                      --             tx_cal_busy.tx_cal_busy
		rx_cal_busy             : out std_logic_vector(1 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(139 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(91 downto 0);                     --      reconfig_from_xcvr.reconfig_from_xcvr
		tx_parallel_data        : in  std_logic_vector(79 downto 0)  := (others => '0'); --        tx_parallel_data.tx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(7 downto 0)   := (others => '0'); -- unused_tx_parallel_data.unused_tx_parallel_data
		rx_parallel_data        : out std_logic_vector(79 downto 0);                     --        rx_parallel_data.rx_parallel_data
		unused_rx_parallel_data : out std_logic_vector(47 downto 0)                      -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity alt_cv_gt_latopt_x2;

architecture rtl of alt_cv_gt_latopt_x2 is
	component altera_xcvr_native_av is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 1;
			data_path_select                : string  := "standard";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 10;
			tx_pma_clk_div                  : integer := 1;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pma_bonding_mode                : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0
		);
		port (
			pll_powerdown             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_serial_data            : out std_logic_vector(1 downto 0);                      -- tx_serial_data
			ext_pll_clk               : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_analogreset            : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_clkslip                : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_is_lockedtoref         : out std_logic_vector(1 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(1 downto 0);                      -- rx_is_lockedtodata
			rx_seriallpbken           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_seriallpbken
			tx_std_coreclkin          : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			rx_std_coreclkin          : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(1 downto 0);                      -- tx_std_clkout
			rx_std_clkout             : out std_logic_vector(1 downto 0);                      -- rx_std_clkout
			tx_std_polinv             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_cal_busy               : out std_logic_vector(1 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(1 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(139 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(91 downto 0);                     -- reconfig_from_xcvr
			tx_parallel_data          : in  std_logic_vector(87 downto 0)  := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(127 downto 0);                    -- unused_rx_parallel_data
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(1 downto 0);                      -- tx_pma_clkout
			tx_pma_parallel_data      : in  std_logic_vector(159 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(0 downto 0);                      -- pll_locked
			rx_pma_clkout             : out std_logic_vector(1 downto 0);                      -- rx_pma_clkout
			rx_pma_parallel_data      : out std_logic_vector(159 downto 0);                    -- rx_pma_parallel_data
			rx_clklow                 : out std_logic_vector(1 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(1 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_signaldetect           : out std_logic_vector(1 downto 0);                      -- rx_signaldetect
			rx_std_prbs_done          : out std_logic_vector(1 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(1 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(1 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(1 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(1 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(1 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(1 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(1 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(1 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(9 downto 0)   := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(9 downto 0);                      -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(1 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_elecidle           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(1 downto 0)                       -- rx_std_signaldetect
		);
	end component altera_xcvr_native_av;

	signal alt_cv_gt_latopt_x2_inst_rx_parallel_data : std_logic_vector(127 downto 0); -- port fragment

begin

	alt_cv_gt_latopt_x2_inst : component altera_xcvr_native_av
		generic map (
			tx_enable                       => 1,
			rx_enable                       => 1,
			enable_std                      => 1,
			data_path_select                => "standard",
			channels                        => 2,
			bonded_mode                     => "xN",
			data_rate                       => "4800 Mbps",
			pma_width                       => 20,
			tx_pma_clk_div                  => 1,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 1,
			pll_data_rate                   => "4800 Mbps",
			pll_type                        => "CMU",
			pma_bonding_mode                => "xN",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "125.0 MHz",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "120.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 1,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 20,
			std_low_latency_bypass_enable   => 1,
			std_tx_pcfifo_mode              => "register_fifo",
			std_rx_pcfifo_mode              => "register_fifo",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 10,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 1,
			std_rx_byte_deser_enable        => 1,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 0,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "bit_slip",
			std_rx_word_aligner_pattern_len => 7,
			std_rx_word_aligner_pattern     => "0000000000",
			std_rx_word_aligner_rknumber    => 3,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 31,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 1,
			std_rx_polinv_enable            => 1
		)
		port map (
			pll_powerdown                  => pll_powerdown,                                                                                                                                                      --      pll_powerdown.pll_powerdown
			tx_analogreset                 => tx_analogreset,                                                                                                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset                => tx_digitalreset,                                                                                                                                                    --    tx_digitalreset.tx_digitalreset
			tx_serial_data                 => tx_serial_data,                                                                                                                                                     --     tx_serial_data.tx_serial_data
			ext_pll_clk                    => ext_pll_clk,                                                                                                                                                        --        ext_pll_clk.ext_pll_clk
			rx_analogreset                 => rx_analogreset,                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset                => rx_digitalreset,                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk                  => rx_cdr_refclk,                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data                 => rx_serial_data,                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_clkslip                     => rx_clkslip,                                                                                                                                                         --         rx_clkslip.rx_clkslip
			rx_is_lockedtoref              => rx_is_lockedtoref,                                                                                                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata             => rx_is_lockedtodata,                                                                                                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			rx_seriallpbken                => rx_seriallpbken,                                                                                                                                                    --    rx_seriallpbken.rx_seriallpbken
			tx_std_coreclkin               => tx_std_coreclkin,                                                                                                                                                   --   tx_std_coreclkin.tx_std_coreclkin
			rx_std_coreclkin               => rx_std_coreclkin,                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			tx_std_clkout                  => tx_std_clkout,                                                                                                                                                      --      tx_std_clkout.tx_std_clkout
			rx_std_clkout                  => rx_std_clkout,                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			tx_std_polinv                  => tx_std_polinv,                                                                                                                                                      --      tx_std_polinv.tx_std_polinv
			rx_std_polinv                  => rx_std_polinv,                                                                                                                                                      --      rx_std_polinv.rx_std_polinv
			tx_cal_busy                    => tx_cal_busy,                                                                                                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy                    => rx_cal_busy,                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr               => reconfig_to_xcvr,                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr             => reconfig_from_xcvr,                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_parallel_data(0 downto 0)   => tx_parallel_data(0 downto 0),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1 downto 1)   => tx_parallel_data(1 downto 1),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(2 downto 2)   => tx_parallel_data(2 downto 2),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(3 downto 3)   => tx_parallel_data(3 downto 3),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(4 downto 4)   => tx_parallel_data(4 downto 4),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(5 downto 5)   => tx_parallel_data(5 downto 5),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(6 downto 6)   => tx_parallel_data(6 downto 6),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(7 downto 7)   => tx_parallel_data(7 downto 7),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(8 downto 8)   => tx_parallel_data(8 downto 8),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(9 downto 9)   => tx_parallel_data(9 downto 9),                                                                                                                                       --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(10 downto 10) => unused_tx_parallel_data(0 downto 0),                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(11 downto 11) => tx_parallel_data(10 downto 10),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(12 downto 12) => tx_parallel_data(11 downto 11),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(13 downto 13) => tx_parallel_data(12 downto 12),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(14 downto 14) => tx_parallel_data(13 downto 13),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(15 downto 15) => tx_parallel_data(14 downto 14),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(16 downto 16) => tx_parallel_data(15 downto 15),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(17 downto 17) => tx_parallel_data(16 downto 16),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(18 downto 18) => tx_parallel_data(17 downto 17),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(19 downto 19) => tx_parallel_data(18 downto 18),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(20 downto 20) => tx_parallel_data(19 downto 19),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(21 downto 21) => unused_tx_parallel_data(1 downto 1),                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(22 downto 22) => tx_parallel_data(20 downto 20),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(23 downto 23) => tx_parallel_data(21 downto 21),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(24 downto 24) => tx_parallel_data(22 downto 22),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(25 downto 25) => tx_parallel_data(23 downto 23),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(26 downto 26) => tx_parallel_data(24 downto 24),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(27 downto 27) => tx_parallel_data(25 downto 25),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(28 downto 28) => tx_parallel_data(26 downto 26),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(29 downto 29) => tx_parallel_data(27 downto 27),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(30 downto 30) => tx_parallel_data(28 downto 28),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(31 downto 31) => tx_parallel_data(29 downto 29),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(32 downto 32) => unused_tx_parallel_data(2 downto 2),                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(33 downto 33) => tx_parallel_data(30 downto 30),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(34 downto 34) => tx_parallel_data(31 downto 31),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(35 downto 35) => tx_parallel_data(32 downto 32),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(36 downto 36) => tx_parallel_data(33 downto 33),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(37 downto 37) => tx_parallel_data(34 downto 34),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(38 downto 38) => tx_parallel_data(35 downto 35),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(39 downto 39) => tx_parallel_data(36 downto 36),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(40 downto 40) => tx_parallel_data(37 downto 37),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(41 downto 41) => tx_parallel_data(38 downto 38),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(42 downto 42) => tx_parallel_data(39 downto 39),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(43 downto 43) => unused_tx_parallel_data(3 downto 3),                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(44 downto 44) => tx_parallel_data(40 downto 40),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(45 downto 45) => tx_parallel_data(41 downto 41),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(46 downto 46) => tx_parallel_data(42 downto 42),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(47 downto 47) => tx_parallel_data(43 downto 43),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(48 downto 48) => tx_parallel_data(44 downto 44),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(49 downto 49) => tx_parallel_data(45 downto 45),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(50 downto 50) => tx_parallel_data(46 downto 46),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(51 downto 51) => tx_parallel_data(47 downto 47),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(52 downto 52) => tx_parallel_data(48 downto 48),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(53 downto 53) => tx_parallel_data(49 downto 49),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(54 downto 54) => unused_tx_parallel_data(4 downto 4),                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(55 downto 55) => tx_parallel_data(50 downto 50),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(56 downto 56) => tx_parallel_data(51 downto 51),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(57 downto 57) => tx_parallel_data(52 downto 52),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(58 downto 58) => tx_parallel_data(53 downto 53),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(59 downto 59) => tx_parallel_data(54 downto 54),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(60 downto 60) => tx_parallel_data(55 downto 55),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(61 downto 61) => tx_parallel_data(56 downto 56),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(62 downto 62) => tx_parallel_data(57 downto 57),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(63 downto 63) => tx_parallel_data(58 downto 58),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(64 downto 64) => tx_parallel_data(59 downto 59),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(65 downto 65) => unused_tx_parallel_data(5 downto 5),                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(66 downto 66) => tx_parallel_data(60 downto 60),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(67 downto 67) => tx_parallel_data(61 downto 61),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(68 downto 68) => tx_parallel_data(62 downto 62),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(69 downto 69) => tx_parallel_data(63 downto 63),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(70 downto 70) => tx_parallel_data(64 downto 64),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(71 downto 71) => tx_parallel_data(65 downto 65),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(72 downto 72) => tx_parallel_data(66 downto 66),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(73 downto 73) => tx_parallel_data(67 downto 67),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(74 downto 74) => tx_parallel_data(68 downto 68),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(75 downto 75) => tx_parallel_data(69 downto 69),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(76 downto 76) => unused_tx_parallel_data(6 downto 6),                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(77 downto 77) => tx_parallel_data(70 downto 70),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(78 downto 78) => tx_parallel_data(71 downto 71),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(79 downto 79) => tx_parallel_data(72 downto 72),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(80 downto 80) => tx_parallel_data(73 downto 73),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(81 downto 81) => tx_parallel_data(74 downto 74),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(82 downto 82) => tx_parallel_data(75 downto 75),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(83 downto 83) => tx_parallel_data(76 downto 76),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(84 downto 84) => tx_parallel_data(77 downto 77),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(85 downto 85) => tx_parallel_data(78 downto 78),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(86 downto 86) => tx_parallel_data(79 downto 79),                                                                                                                                     --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(87 downto 87) => unused_tx_parallel_data(7 downto 7),                                                                                                                                --   tx_parallel_data.tx_parallel_data
			rx_parallel_data               => alt_cv_gt_latopt_x2_inst_rx_parallel_data,                                                                                                                          --   rx_parallel_data.rx_parallel_data
			tx_pll_refclk                  => "0",                                                                                                                                                                --        (terminated)
			tx_pma_clkout                  => open,                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data           => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                     => open,                                                                                                                                                               --        (terminated)
			rx_pma_clkout                  => open,                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data           => open,                                                                                                                                                               --        (terminated)
			rx_clklow                      => open,                                                                                                                                                               --        (terminated)
			rx_fref                        => open,                                                                                                                                                               --        (terminated)
			rx_set_locktodata              => "00",                                                                                                                                                               --        (terminated)
			rx_set_locktoref               => "00",                                                                                                                                                               --        (terminated)
			rx_signaldetect                => open,                                                                                                                                                               --        (terminated)
			rx_std_prbs_done               => open,                                                                                                                                                               --        (terminated)
			rx_std_prbs_err                => open,                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full             => open,                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty            => open,                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full             => open,                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty            => open,                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena           => "00",                                                                                                                                                               --        (terminated)
			rx_std_byteorder_flag          => open,                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full             => open,                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty            => open,                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign         => "00",                                                                                                                                                               --        (terminated)
			rx_std_wa_a1a2size             => "00",                                                                                                                                                               --        (terminated)
			tx_std_bitslipboundarysel      => "0000000000",                                                                                                                                                       --        (terminated)
			rx_std_bitslipboundarysel      => open,                                                                                                                                                               --        (terminated)
			rx_std_bitslip                 => "00",                                                                                                                                                               --        (terminated)
			rx_std_runlength_err           => open,                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena              => "00",                                                                                                                                                               --        (terminated)
			rx_std_byterev_ena             => "00",                                                                                                                                                               --        (terminated)
			tx_std_elecidle                => "00",                                                                                                                                                               --        (terminated)
			rx_std_signaldetect            => open                                                                                                                                                                --        (terminated)
		);

	rx_parallel_data <= alt_cv_gt_latopt_x2_inst_rx_parallel_data(121 downto 121) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(120 downto 120) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(119 downto 119) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(118 downto 118) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(117 downto 117) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(116 downto 116) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(115 downto 115) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(114 downto 114) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(113 downto 113) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(112 downto 112) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(105 downto 105) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(104 downto 104) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(103 downto 103) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(102 downto 102) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(101 downto 101) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(100 downto 100) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(99 downto 99) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(98 downto 98) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(97 downto 97) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(96 downto 96) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(89 downto 89) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(88 downto 88) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(87 downto 87) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(86 downto 86) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(85 downto 85) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(84 downto 84) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(83 downto 83) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(82 downto 82) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(81 downto 81) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(80 downto 80) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(73 downto 73) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(72 downto 72) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(71 downto 71) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(70 downto 70) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(69 downto 69) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(68 downto 68) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(67 downto 67) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(66 downto 66) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(65 downto 65) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(64 downto 64) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(57 downto 57) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(56 downto 56) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(55 downto 55) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(54 downto 54) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(53 downto 53) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(52 downto 52) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(51 downto 51) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(50 downto 50) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(49 downto 49) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(48 downto 48) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(41 downto 41) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(40 downto 40) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(39 downto 39) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(38 downto 38) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(37 downto 37) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(36 downto 36) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(35 downto 35) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(34 downto 34) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(33 downto 33) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(32 downto 32) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(25 downto 25) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(24 downto 24) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(23 downto 23) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(22 downto 22) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(21 downto 21) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(20 downto 20) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(19 downto 19) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(18 downto 18) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(17 downto 17) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(16 downto 16) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(9 downto 9) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(8 downto 8) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(7 downto 7) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(6 downto 6) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(5 downto 5) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(4 downto 4) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(3 downto 3) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(2 downto 2) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(1 downto 1) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(0 downto 0);

	unused_rx_parallel_data <= alt_cv_gt_latopt_x2_inst_rx_parallel_data(127 downto 127) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(126 downto 126) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(125 downto 125) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(124 downto 124) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(123 downto 123) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(122 downto 122) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(111 downto 111) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(110 downto 110) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(109 downto 109) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(108 downto 108) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(107 downto 107) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(106 downto 106) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(95 downto 95) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(94 downto 94) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(93 downto 93) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(92 downto 92) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(91 downto 91) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(90 downto 90) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(79 downto 79) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(78 downto 78) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(77 downto 77) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(76 downto 76) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(75 downto 75) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(74 downto 74) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(63 downto 63) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(62 downto 62) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(61 downto 61) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(60 downto 60) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(59 downto 59) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(58 downto 58) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(47 downto 47) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(46 downto 46) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(45 downto 45) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(44 downto 44) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(43 downto 43) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(42 downto 42) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(31 downto 31) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(30 downto 30) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(29 downto 29) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(28 downto 28) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(27 downto 27) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(26 downto 26) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(15 downto 15) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(14 downto 14) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(13 downto 13) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(12 downto 12) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(11 downto 11) & alt_cv_gt_latopt_x2_inst_rx_parallel_data(10 downto 10);

end architecture rtl; -- of alt_cv_gt_latopt_x2
