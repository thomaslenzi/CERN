// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sfdR7RJ2HPvTnJp6qJVZ4aeTHPZ0EfVZTW6HR39xoy3qisCApJsP59RdvU6bGVcj
kl/iV9muZ94Y0F9SLfSfOLXCk8G4sKpOwKQ5DOumGpHxoy15xSHyyOmUgOvuRfRO
I599tBQO1YkEj8mj+i5fUAAziFu2jSEtXv6Lv9ba8/I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6016)
UfuF2BHLqoijPFho8eQ1O6UfzlYtlViSwgpmOfoihBVwfuRVL6bfCUmT2P6SlWVt
AgvktFyTi4rAOP+lVyfxdXe2pGaTLUv5W9LOr4tt4hJllB1wUnjID7WX/666oYWS
oV/uACL8H9V40zX5gVvWcQq+zfTYtlRvXJooz0X9v/GfjbGx+2e1gP3RyQ5uU9FV
mqpz7QNI0c+AUH+4ZwP7Zll6gZKkEQHGLe1UDa+NxpC/XSAkDF+UqXL11G+XPSTW
yHacNQ5uzwCV+f6565AqIS9PWr3M8GuqzWUjcOIb3XfeIfWaQzQlMlXzNNPF0Qd5
KUNnWaxMTJ23/assL8rPIpJO8WfW1+iZzrLP5tWKBUybGGv6NnMp2wF1e7H71OY3
c0nAAe2SfKKY9wWUdCEQjQeI3jvJmiN9uJa/Ts8NlN+iLGS9gSVH9US96VN+7BjI
qddcGaHFDEaKTm4+lS0YsGu/CdpHVQFq23Ye+K1SHQ3wJZVAPtrf/K3hPFdWDrl5
Q4IXWFaT/ECBxSJmm2Km6hUuiUdDdjfmi6AfbBq/d6x3INg0MePnam4aw4iLETvJ
rqrWukQCgcqi9PZOpFe1YqMujNcKzkFv04itGISFI/k0QmkfNOjQldiVA1+R9v5T
1SZZ0rM+gKZ31Zv1NvDzjSumzO1TibYfTUXOUakqD/Yio4n1xq599K7BGhE0gtY8
KV6ej+Ya704ImNB1KVEz8LK6Dmsg57Ot6W2NmQ4pIM5ZxLgH014jy+Vtbj8EvteR
53t5wyzNemCs9Kddc986sMydkAzod06vsBIlQ7vzoiXtu3GNVafdbepeB17sP/x7
27wfv+T6hxDaQbUFXp63QbjFcCHNmEJYpbq/QKToHxFSDMj0Qhcbq23OKHyT0IjK
Zbs4J44VQNmgld7p4YZvkPZ1bZKx1gSCmTZvCB6hvbgSEoc8UXl2LJ4oX+eezZS/
gNHzOb+NpiEgGmEIGYU1E9phjUNXWPLtkppFz7o1rcKv/HSi71EE63jHVLyNf9F2
e6Px0OYauqKCNDf3HMoQ+yK5t0TZeiVWT6AEXkX+GfyYJpH8FmaVexCg/hz/udss
krCIrFTEujeg0Vr9LCCwhHTrb7PwZynteVPp+p1XePMu7uNeZ7iEC7FTLNNpGi6U
b4cpNizIwQlWEK6jlccRqkFNwbncXGD/BkVqVoxsD8JSskXf756EChcC4r0acZwA
lhUoGJXdNy/d9P7cXVevS9ULp1/VVNXTK5V9/pOE5vKrFcyG+WmTvMnJ5Vhn9Kem
wY5AOPYZYxvgTRnsuZbwHxh/vQ5pPQ/F3m0YVqGJjY8N8fK8SFyUaa5ZZjCIQ9W7
xtkbq8l6PFv1Dv8uIcb+qQyAfqGE4iFTRmXwTuG7etdGtYekuM/MC2NpVrR5N0Dj
VVJEQE6iLOJAzJfG0r2evXD/xzGXmZ+skyjqXdij5k8Cde9KhHNjgAmEwNSXhEFL
kQAx9Zhzk+GqWocJLloxHU9MmmZDoaHDe5iemVbsHLuhIyD7oCbdWmLatTcDikf/
lUJ+VhJbSpEycB2tuK+Ni1lDn9Vgz4peX5DUFi85bSRwqiOuVdhI/uUhmQBgZWa/
OPrZeuVQvUrJAeHN2RaLl1am89Qxc2J8aXH2962sc3E7Y6Mzx9LOFTQNiB80DO0K
4x8lKFRQpza+Jl+ftkkTGWeQZffe3soHC7bTjrlBUgv6Y6YzfAFHUjhljp+WdMmm
a7kLSStviYB5uSUDtsONuqp/IvOhlJEfLVJmDj/BjiFs+Dwo0eMc6hmzotwSNenH
BbbGxxYM8nozotTgGZRRfMqgD8gAZx0YmLaaaJe4ag3o+TBiB4jCDPSSLGF5IFly
7eikkaob12s8AKulj6kjmVzGtRAc6RfJ7DIYe/YEx7fdCTXyjDWSHSzGG6RFlRNl
QQlWPVHY0ovlI1YMSHib79Q+YCeGFwuucKhQztn7wmJcsyyeE8IOgFGJI8A7U2Ih
+8FFqqerZKbJSJV9Ba3+zXqplrP52UNkza7iJ82Qdpx+5B07f89VY4XaqZbule6+
tBFq+KmCZPJ733hlkJwTo/Gde6Xp/G7JvC9n/J/N8p7RbzZurA53zIvxU3L483/h
h+tRiDdI1OkJVUcq3Y1aTNgVRogJSB+VXNfdTEAGL3/S207uz23OKPUBeNjd5Okv
tXLpHIOFIgihCzsfPfHswB0BN6yTTSkprrAlhcwXYKkz56jqSul70MO59OX9INVy
UFf56KWCYpOM77obUxxLHgvJDTZOX06+z40SGSrt7lS9IKDvwBa8vMI61qUKhc/4
/CglpqmoYsP67NIIGVyAhZan7lbBcIKZ94U9HMMERS99BEu97iFiE0rf0E7Qf/cF
Uzc+xzif/3pMah8oCHOiS9bq30HGMP3tVzEGRCLxOdts5rrDz4tjjWM4kFeKmZQG
HdggPtwbLdlDxA4TIP+KEIiHt1S4J3XEIh8m34Qw3wcI8TWYo+agkHjosX0v1AM9
RUSdfzSc8SFrdp+qmQU5rxXfft6TXDnaEaQS1zSDprnlb539atp2z7vny33ePIfs
CitNprWX70cOPRq7qwvhJIuzl2BoVq5vM2wd56A8PnOwhfI1G8Rj75xX3Gw8PqKQ
i33vJH1vRiitEffpsNA8IoPgYfQIjiypgnvjc72vvHS0PgwdtI+raeykUt8s4vG3
pkQ6whgNyPqF4wKLDLSRJ01BvBbblj5gJtmVTuprfC3eu7si7cIaI6M2LgKZ4j7j
VIUr8+aXX4FEkzwmzeunZFkwJT6CN6uVwWjkkLAuEsOd2EmUJ2ie9pjTG8iOYHCd
39cB1sgUOmOZ+Ly4+orCZEAW+fRcumwni7Y7uaRtfJsECIhUVjimBOwTYtHTTFJl
hskq3JEbUgz72juupUCu5S+hq25Z0HEwiHa8HRo1jsA7KeJUreLtaa5zEh0YY7/r
mjVQGkZz4WsvkOzPtuQX1sUa4HK7266Me+cAOrU4dFczgTSBATXUUd9HAwDse3rA
wcHZgmIYsUvhZRhc1X3AzLN9Mzlo2h3bsCFg46S/dpK5WpbosY2xzOxyH83n2ZAE
G93ApHGfOYtZpRBCeJS5ApgWXdoqYj216jDlVqGi3GQICBonBTi1saDO7/KH7X6G
R2wyp3xkZNJvvfU/kHChakPLemuXih9CQWrL6ofIgqQvCVUN1E1EQc5vJ9f5JAJH
TVVyPfRgL0nADZLTIwS5EvYOhA2Z4K+7uORoycVSF6kSwEmZlEjPq+zMr3h6kdEB
gs+H4OYf3XXuE82vBjrNojZBmj5T49JRUSA/wOBR8oo5WZWeSvkdoSDDpjx6+gRN
abVBiU8dioFTittxQ4IkNAVql40Qqx3JDnfmae1Acrpn1TdBxo2aGYh4v9auq8vl
fC6sBTrX9gwlWVGd16tVngS6HKMXVsGg76h1GwNw33MAFv4pjMXRokq8ArClYpNH
sTHAJp0acvnYFM4sitTkApbEgSbbrAVXgygLc0FeVf/6s3qmRdmAgMgTpWqi+Ora
mlHgzx93X/IHtNk52Fg5f3uQqi0ehGdxwnwwoRWV/AbKSFpTqWlSZPdI0gYb6O5a
AayEIyvPpvMueYahbPgzO6mpprgu0ouOeSXpsIzmpePpvtuo4cTzLxQ+n6Ctr2th
tJs2ZHiLer3fMnzrxusVTSF2AJc3SJIPh3RH4x3n0DAunuOyoOuY/rVZU5AlyWwK
JZxwkvbhxFD1IUT0cb9YyxrdR9XE7xdkBDWkXXzcvWRTh0uuDd4pI382DsKju9d2
p/00HHe2iCqTWaSPii7DTb1K0wo0dCzflwoerjFLsabcwwZTnIftN3Lflvzd3l7V
ee2lDWhFMTzZVh1yIts/wA1p/AJ8J3+15Jgxa6lhrZx9GdZ63OcPrIbErutr2F8c
33Bv7Tz3TYxR61uu4BOPAXfVFaJY6un/NB7rYKOJ2tltE7QV4hyqAVwx1JBm259V
kQxLxEl2jG1jruFeK179ENDJwV/R/Tv2Dgr8WV0BSAD+kh2uw6GA3ivUiU9aZFVA
pEUNSDlRQzV/BZ3lMFQGDLPKvBpxq0PscCM4YUxAJSOMe4duW5eCYbgNLz3Dmdug
nD+2Jc5KMmEXjSiUyR/Q2PaNj6ra88OOx93hWLLy5BtHaJq2b8SOKkvm6/ZpbaPE
/vnYquvE4XSNUuaUClnkrHsY+BiC39nL+U1zuc9uh2MOSc0b6aWo5EllpNm+Fx1q
kGBQ74iCoqW2ksEf39mA27EwW0IZ6DvGscNjrEUJ9qFpL3WxOkDqEc3bVYt64mDZ
ecJkOkbBq9v3H24ykAodgqEsHhRZCKemSHrMp00rhgp2+OP08Vr9ujzicRM7vDuS
hsb4iC/oVd2Axx7oN0Y6xbcSX2C1THBzmFqStRJP+Z8bSrHnoP3yptYXyhqWf8BY
Ky0XXwuCl6siUJY+wAh46p0/eVAFdJOtptRPh9GtaA7JX73AfeL/NNLo4SJOqWdj
TqRRV+ExHsHcIQj7plupNVdAWMIkIznPH8rB1i1zV+UUTqXJj1HcLpcEHBfY5m/s
8CLldKEsFg12vfvjOjcmGynqByFUVjWZ3csyyh5HAyTNVWKl2oLBXthbdNfCmrGE
8Xnj22Mo+2DmaNKYwFIiuKNHVzfvCc0xvvi3vfZrJX0T8dvqDSSH+pwpDfzTEZ2N
d49KmkqyaUaoH7CeAi65LW0LDrktS/CFSwK/98YiNN9Y8ty9WJ7XH/Brr4Mo0bxJ
UjZQhMNGOMGc6WLWJpgS5Ov01G7dhk4FGfziWlvF6qvty2J9UcumCcQfuYMtq010
cKgmcNo1Xf5iqbwaSKFmJg+0iEGf4/rs0jzdk1iFJFLAtAiOF2H4U4aLHqq5Cjv8
tJSf/C+D90R0JjG5qGxLwj1lUxLYVgWUnlTsr9E5mFkXRTRPa28rxRbuXz/1hCww
SDynvvBRsgyLXFrSmpXC3g/alqolzNjhLuDx1aEmuf53WdUwlz23DgHcm8jz1b8d
QF8aXci83U029gcg0G0hdSWNYqt2A4mljVK/tt/HEn8duMR4tTNX1eZtkQJT5MgH
AiEwUmvTceTOifPx+hWIuxdC6WVuudZDSkwXTZFqCX+NZydmJHFx4d4qhLdEbZkP
L40jtwkQMVwDwirq38e77N0fXURAGgPaFl8Qgiwv0VG7T5OheRucsz/BaUN8WwC6
1sKN5r0U4amr+XZp4BhYSnrpKIpvEj9cVx7YSeb/abUzLOu89TdKUggu0pybMfsi
rie61cmxHTHQjvriBhN+vto1OOqmeuqGPbml54oIjpzsOEV5DeAaWngtBSz5Lfm2
dYyVeu60H16UJy5cykX1vNIR23uQxVo65AtRSWHfLWmJAo5oyxZbAlxZdmWwTE13
Sfwizo0asNXqIbF+7uvLl45od/ZFI0KZRXnRXOmx26yVcMmTTB1VQ0G8C1JnDLAp
G3NIUA6M1AfzIL4tG5/6Tvrk+zDcg/mI488Ci666ZJ7HPo8Hl5g7cx0x4fqUTaIQ
wzcC8mrQCF4jDCD4JQTYHYkzkqjMmINLgWsGRhTrKHaQgXB6hWSWfwPqL+Yzv8W0
qRtFUaMoF7//EIew+08d4WcUl/0bXHaiOxpHdphcVd5dG77kQTtDN11BDxN4q0I4
vi4BHe0znyHjvEWOz1fDxemKhQIN7cApwlaO0jgdQFZ7O8mlSIY/WOj5CHQoUTPx
Z3bC58nkDDD/JRUvuxEOUt0Zqhn3qiIVjRCTPJbsvVorjsdNMfuEvE2NsY0tBmD3
4UoOu6mGFmndJVFlDqiVUDWiTv+AYtLo9RFMNeJNebVL3KJvkSTTC4QDnswYYNMs
ZLFpiolU/YxM9JERZ+QnDEzpxlshQN1/bIwj9Lo3slh4jfNQGtE9OakPWvoLRvNh
gy1JWMEbRrrvrBnHlvpq2ERY5addihsMIBJNOm3xK1gXdsqS+SJ/h5jK1lSbGGo9
BJQ9eLKTHWt4uP9QX9IE4y4wwNTU9MffJJNoY/V4FO1mPq9uP0U/IQL1OGrCQBpa
fg69MBO7r8P/OT5Xyq1th4GceFEwTknnIaRMU6x83A6JPx0vX7zEP46BWomSWhgL
33gbo4sgz4kiJNR67VNYv0Y6wa75pK++KsN5dQyluGmPiRDOVA9+Cf9qqmSyAR2m
ay0bfMcnEeY4Vhr7FLfW+19tmStSZmkVprOovL5QbT4WE9LqHrt+XTNoJaHHeJBe
UQza0BxfGuhvyhLNGZbhqr01iIyeclKJDNbscgNDQSkUErK8taNeXK+GbjVuVwTy
6tBntI74nvuEEwW8FPINwIVqG6Ouc8xXK4HLOCympwjHCzEa69QyhVrVZdOaq1du
pruqyQVMCFlfN4WQkJQDq1eErutpCTsafJTk09c+1Z7117MHYQKFvCeBXFD5nzlB
ANy+L2Mjaf+Nbp9co2lkSTA1pxzu8sk/9qdOPL5RrPiQHycNa3PlUqW49LdCR/H7
jVcjqWfirLzvmz99yDhG0KHO8ENjwkcilztSGKoj4Xc+a2RQCw04p4o1kJusXpQC
OYQajCyUDdIYIkGzgtOvmAsqygBCweqRb+2In3SJB/Wh8cRZCi+b3x/iO9K1jMnl
0ylCFVCLaDphiAu+v387coyKQaZE7fggnZlYn8MncEsMYdEK0Ck4Nk2ZxDbyffLo
198J5L5rcGCXbOX8mZxHSQjjafRbW45NLKyBqMVE5RRIr2at4JDZczl3H8zIpU+G
OvEBZMuKb6N8u/vabDWTa0hQCVnKvmUsz3UKCdVG4ote9mQXJUXsoAFStHQDAa1c
3EqtZM+Isa0nCVFQGlv6AJtGCxivlz6RyiUQHtYMHFecjaK3QTAYPT7IJWL7uUE6
1lj3ogDC3P78/yTRlJ+iy+4jXdWkF8ZGNwCnJ+5FEz6u7WnWhk/g2IePRvHHryD8
hgIYKb1R1STYuqoQZD5wz6AS00FWPldTaZpQeNKQkiM+hd6QdK4OnvAxx2yBRFaW
JHwcc5VtgiiMRk1c8IWJmSTgasQQTpcVK+Y5WMFqALj71HXjDNV2VTp1rCYhD6z4
wOOOkrJ4zSMoAjKv1VlCAl0/w876mkNPjeF/XJtP2H06/Bkxo9EAuYrvLzo8W0NW
lEbVj4NB0ZBd4+v1b/Gagwr17eMDFl32NF7W6YCtRULDTttu/kRKAmy8D6WZZhfs
qW/TDbxfxgowanJFkYVuopCgasEv3vOAu5i3TILqdfhQVaqI3uheDo6Qwv2xcPFa
tuvU3jDJnYSJ8qoawLzTW1VcOSEjMERmzkeIhuo3k6wYYrNlVdGfrUrQvS1dviUB
yfW3vwEpWreIfi72+IyPCQsLyRL+Ux7Zp/EniTSzfsm0NtxruKPTXlwIP67RZjme
hsSl12oVAWfkbm4Na4TFJDengt3B6h63RmHk0VfDm/pAEvh+KZexUGltnPQxGu/z
0ViFjSvRAfdPMCr7Y2erW1M+02CxY8IuXyI3Ks2rFXMZg6qBJvQM3ewUl5iLQOuc
eW5hyCsjDIsGA6WKNubAWrn6T4HrIN1gxXd8LAByGqK4dlG8RJBe1vc205jlWuGg
HnDTgZoxA868sK1wCXyq1SAaxxTVkdS/LlztqsG9+m6mS4IEmpQBxw3QJmW/usys
s6ZF6wOwknl8UfChLv6hYHMSBVS4iUSXsD5+EAkpJvvvv5y9WICQvJdGbR0jdAMj
MtYQk/BCzNzaxNYS4q149G535OOQdTgEXWJP12ouDhsrkfiny+B03DR6A17BLCT3
u0ZK0DVfYRauvN8yYkyWRFoC4aluWqvoY+8tWXzrPdLHDN+KznH9ytfVT81f08En
0sgmyXpyvykKlshn1IKtpyaH9KbHfGuBS1/egGmNVB/HsbkA5fqPATShY9eLh80o
Cv1fQMCz4wLQVO16aje8XCrd/+Pad5XqO07dYEC2E1sAlAWw5LNWi/IBgQQ925f0
c670lqdAUZ6J2vnUenCHPitBD++ZihldxMclvLZ/7KsIiwQCL57mXSNPwhtMLzUm
wK9i5D5z3MB7rJf2b7PYIA==
`pragma protect end_protected
