// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dGz2ey1QN7BWIK1XCr8EdYqMAyZb2eDIY/Ua7S/mq48FFoNrVHwFX6yFRxwVEM5z
N9J60IAzQBODM++Uy/WM2gCCJT6ieF2w8msYVAqBXAe3hXlltYFzR2c1eh4BNaTl
vcsWF2xNM5x+3m4/IPK2V/V8aOtDVPXqjwG8h70Wclw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5216)
apXBYx8DNa3V04e04R1ecncJq3mjlhSAchP9202ZZBqPyMKFK87waBoogsx+uKK2
GU9LoPyNbnEvjuSn+zJizcGAQTbOAOKM3+TpZrIflaUehymB9YbqPVtZ7V+4bhJu
ifZDLbtRr7kpd2auEpdpHQCIUfmqKwVGs4txT9/mJ8gVq+RUz/X1mTkLxb/J1S1j
QjC1nLeQ4r/fvG4zzuv0ZFAeqQlPrrdaGBhWz9q4GSxKNKmUiJ3DcI7fpUihz2+c
tkmeNl7O5bJTf/izR17WFG1Xj3Oxghc4NAORWh4UeD85RFSRYhiZoYmZDO+/PbGG
drX4xGjNv9Ze4+E5N7Iu2dkcha7LkgC/XnoCuQYlGkOPUKnS/MrQXBwZI4d2xG2/
V7kNbVyVjWB8YfFmoLYa4h2z9729i0gHgou7pUNTKOoloGef82+NYPR4X5SFkiZm
m1X7q9rY1eGaWhNlFlQhWN/DomqrN9CbsHbHrtMbcpGhKDV6fRBg+zqJknS/CMiN
oIb5cRcrG0+fXJrDVGRcxR72UO5VLTtfC9Ku9+zdjIEbpFzC7BkC4IdZV64jYoli
zjYtjGmZjyyYrfiydsH4h47flFEGh+TzHueFVxmDN2ZcwU1WnuxuijcOgUgvuwFY
A/Get1HqBuGMT06rQoS5XftDbuPyjaFrUwQ2RPfR2REppols3K81OyWSu9k1iKH2
per5/gIqDtQ6XBP8P8VXtAkqjLrD3B/t6XmqTV21cwh5932zmMu++Or/U8a6Uwnv
Pyc6/Ap9XOZiMiGkOnJLDOhfB3zEKDvupk68sCoGT7cSEPomH4lzA9wG1VNIkgn0
x2tiqe5aWMbIuXjfdUC/palk3tC3qLKWBjWz7pFXEXOHJexprRS8dmnLK+6GTHwG
3HVI9xcz31La/ktqx4TdrSonQA7m14xWzrFKChAVxRMaNFj3bY9jxlaiOfbWdPqn
KsRIWBGaBnqoZ8irvrpxdXuY+r2Djcrm3smsQ0PGGB/l/pmCz34jNMBswH93psV7
DomXDSuqn5kdfRyHmOYlskvTSpmhaSjFjRkEIhHcIEfzLqg5FS5IQRR4whGXvMKh
J5W8c1vcLQVJCMaZFe8zaARwjW7OZ3+0A3NnALXc6/svzTJ0LgrBq/RSL7lSv95V
fIeAzaUdxR8MQ8ce5eGF1cfgp27ZAqM/MmjwKRtr/wvw98peB4imFIUl0XSdTS+6
sHZPKOZ/Y/XoMyFVF8FHg0958b67NkXJX7JZ2bH2x5g0paQD1iU/zA+FWWa2Snvi
V79cRrLlD5vTvDQdJG9rUijnbh3+tGnRahW//cxo3nBDRurd+uCiOZjqx9Zfvfgf
73FhRckrQrE8wIfXC++MNpFtFOCQgPojTWbdYNeyhHlkCLsGjra0phQ4+OlTwRZG
lLYX2AKNMxwzqq6W2akAhOzP/hPHwnRCFidml/Nbo+cRLfmE004lf7lcBYafGU3V
hokHNGZRs1bqA7v4Twu9Poft6jl51RE6zR48IbqUBl9k5g59XwiQUKmfMRXIsIdI
//QpgESPCyz96EDfWwTVN1Rb5ciIFvymoLpkI+5zdpq8g122hiWnCcwsWWs/5yC0
F1GffNwXnccXanI3pB6lMMEqduhh48IMs/UcBteVSYz2FIDxourhXRxdFL7TU+Ti
dPyKK/Iecw2FndEtdRB6vzG3vwxeR2rcGEpDnGwHN5G22XiMaD7x1HACXU+KSDAw
LcKiLaUhIXBygYsfjGJxnQfib6Bg5M4F1DPKwfTn+t/VLH/sO0/ElcqKRKTaS35o
rx4AkTzlTeRSWc/9DwNgIuEWsx9iNXyg1/cjrAK76ea7KaAYO8CyA8C0zEVUzpT/
gg/uoozx+wCN68bPb+rfrWLSVMTQz12FXjgt/KNH9MLXtCvVjKUYR5DEQpVf9b/A
MsZSXBjuVOM72Gyer1p0VFc8cEs5zSrZvX93lXLkBuULhzHadt6kzKhaEL+aiBEX
Vaa9hF9nLgLj3dSe97oVJ8UnUZJpOr3jwEFdLcoV6TWNnoPPHuPsB+uMqcST0mCQ
SCLNiYyheJPStP7nqncNHj8spViUYBlvaigTwEsLTIcq5Fj+sER53fzAj59RjU7h
5Fwn3Gpk8LAVALLeapGA09Y48Gy+VCVNs+n0UwtWKknsOeFxePMCcc1fa2e6rxv0
JLZcZ3boOTIyqjJsn8kMKMe1urc604B+12ubcLOEpt0AZrL6A/Zy0IRkmQfTB2sU
UbBqQ/j92xm5HyOAKYbo/SmoMmU4HZukJZJTQRMTBlYjm/8mrTbNcHv0Z+XqXvS5
snUc1rPBLkroX6PAtJpJb+kLH8qq76ZWN0MZvEaEGEmJJ17B++m3gIFNSDK/B9pE
W5cZwQWwgUngHW6c4tKnvspAvvV+DT2FfDQI4wZRJkbmYsqQWBCUN+fgURUMdrPx
Pda66h7B98aWX2d0706XxJuwuVcs2lLhLwEVk/Q4/3DqPn6seMrV3bO4vXa+Ugan
XhKT7NcAt+YbzSBU11eHAyBaP0qNpMKgXzSqiPu70K8W+JAOKdIivLs4Nzto5rMn
5S3LgJL9Fv++yg5xXJ8ksIqSumDAmycrDk+YNfRRHoFgY3mCYj1AbbG/dCjmtLot
F/MdyKgE6Q2B45jtRSV94FDvWGBPQEEHnSfa94J3OdV/Z4EGpLkPd8alwHjdUar6
G9Yz3+mVqHDmS2djsT6SpQvGXPtLKhx1/CnJXqyuO62pcLk/O3iyXN1+E6xMT97z
lITIv2ltKC/YaheIjJMGjYpmU8kYMw+dU7zJqJQUXYdo2w9e1O8R8I1mcU6eFVcy
jzSzzldPyKbcC4maAD/heghWjpSfO69DUHO9NqZt8ZODpS/UHnv195DAaNIAfrOf
psDIi4BE/6hXfGT+Jl98FzHYDbqulmwLJuCo/jwXF+B0MIuOXI8ZDKZfqkM47fRa
7rbB5zJi0dQFvrIh/zLAqVWIzqNTIkWTkxcGnJ1WN/scUxdpWUjAVFd5zCZGxI0+
MZFJGChBQrgZ5iUMmzJfRXk2+/pkXMVMpiqb2ueq4lCAtqjlqf5qmIHqoEh3aUZq
oA30Tn/pSV652ndd7wNO2BXIFdPdp9WavNp4NlSsNLfiLudKeR5zp2QnxX8C5wdv
/7J6s70HtXYXg8sNqymeTXvjcSMh6A0dQkGRlalApd9Spd9kHaLt680/O9xhxNp1
8kByFvGqR36BlwK6++DjTgo9yMasgWLD2LiqrV7w7Lz29V1we12f0FhedQuOpBMC
GHtTYYcT0LWhYyf6vBI1UKTgH7xozo4rkl9Oxq1sUmMR6/C0D5hzFQ3uT/mQZrhz
AgBdv8MD3fO7M+cszrRr+QTq6F5O3U4zo1MCFzT/k8gZ/t9mqOoitnfRmN6bVHm6
D0a0lfOGgrpMqb6PkOAfy6Oi87JuRylCqhBP8kkiHy8WFXX3jtyTtLDFD6uuYuPE
9RZHgHcaApNtCE1lkJ2yjpfEcNB8Cxarmh3v6fQksBqNW2Oq9FBwRVuhU2pe+e05
LuC7eURnWP/lJZfTkIEQa7SXQW6aR9DeSpdyUwxs9jXwEbTT3+MrxAN3GMRL9igv
SD2xHau08trxQeSHUyznLa7Sa1UusOvT1w9wEAlFlOGdMkN+BapUptFMiGDLFxyx
lUjUDVFzAvafSj6ErR0T7uNHbtLjQcI9N95K4nYhlgLgIVV1eVQZL+KM5Eobd1id
wNK0mFmtIzqI+hfLWTePCQP4VSuPKrga7uuL1KYmkBaESfCR6p9asqUUC9LLMGKf
8LxGLrkO9q+ABHsJax+K9XtQX3teWTduL7Nl1lX5vVYpBWYK1ZbDghYANBEAfKll
ZHeRGFr0u/+EZb7t9LZx2ew3UU3tLvqBpvKNhfDdS2r4dYcWCxH/4mhVOMgzu5Lz
xzVN/QZSCvR38vcrV6QruOoyLm4F2qzwB9fXqwA83AsB+AqfhrLZa5uj7ZwCFEGY
X83GwsrvzsUEaCGIWcHDe3hBPEROuSUFEgEnhiCwmjAuOLM47uC2yUxArJu4Yk7X
YxhNvD12NV8uvXla2M2Kt7sKovKwxxgOkw8YKGJ0Y639z5iZItg2Ng6uWGEjzRAL
Vxtv0EUavhRgFnrYk87tCtbifqx8WiwVYN1no616lBcnETDttCGfLDEl0CFF4W1C
q/dnsY619Wui3ZfT7oaWrFe8jTnPEZFo4GYwq/mBpdIeiUMiKU6bBDAeDTo6TzpL
7VBteGrBP1EcI5ihqTSlGFg8pBZkrsBrD1kPY2IfIA6+hV05OXLF9X4oHpAtjfEF
QxPgavnFEj5KhiSTM+veIQf8y86x/kXTHutcifV3Li+sCQk4pBvCmedcbnoGVI2C
bqKDU/K7FXpNZhlzbtD2Mp5EO+CjhmvBAVrtn0DxAwHcZRb1bTX0kx67vpumLYAc
2kQz91cW0epMLjQuKU27zsaQawcx09tY+don49r1DwD2jvIfwMDAFkYtcZEi3Uc4
0CzZx9qfycywLUp58Sg3HD3d6K2tEQ9B15TQCHq3LW7e75X3KWsbFIUMZ/EGt0Xj
o703MDvVjEE3F0fZXNYSAGD+W2cSf0PlSOEXufHtDeW6SSlX8CWzAzTibKoC0Uhh
bkhWoiG3PC9tguiN4FMJHMjTIGffivafCQ1rV4XcKcdj6BBV/D0ZG/FHnOte3d3X
EAdVMv1VqoeU9jaX1aKepvjx3PRy52AMLJHOAbJW56hMBw21pL1Zvnjns57o21NN
d780+GP3vc5t4R/zB1JRD4kxqpasshTiyA70EagxCbK798ed6MWAfawO89d9ccAZ
6XlC/GkI4tSjrdUiSw0dp+5KSUg4POJqjFPSaF0lBy3wTAsdApKbzLZQd4f8vBJi
lkskfDelnujsjeYLkAyiYVAPNNDLWB7Ey3DOTEyAnA/109HLRHTpR8bnDLmkgLxD
2pp/CjDSGwrlREli35H/jaWQvPKTAZqK7TDmkXcTvkwLKyHcPiZulSTdqwsZUdYu
+zyctME38B5jSkte45F6TTfnIBdRMDXk5IwP3kV0rqUFa970a3oi00PmPKZVMyuR
QibddclmrVC7QwFjvlNHvZNqiXHIqRmDcl6WELtmDkUXxOt/a1b7IddPr79wwGnE
fcdSE7N01QHMspLFswMU9S2haUCfwuVuHkbshqDLKNclMqVYOB3GNzwCZskJfs5Z
hWspNo3B2/+nlm7BZBqGHqh+KuseUVwjLZ+bYtHJ0Afjsro/ZMIJlEfKK/nYeohm
g09f/kTKigAREzs1Wf3hcb+WoWFXaArm747vlPv0yC7AJ3o750nHhIlpf8f0iJHE
+8dw4EAWuaC2WHX/cuE7gJ8jysVvJzmTiKavDJ1L5E+h9aP+aV6PxplYIA9Qke4a
JelfceZFM4Zcx0jcGXNgwJPUoirFSV/yJm3HNou6TrOt85jHr259/3xXVUgCBOyf
It+OWFYZ5CrcoCRDAh9Irj8u0/uoyJdQr7s5LgvHde8J3GDLMXHnVTPt0l/fzbCf
iyxQTEbu+0HU6XGAXNXevC+CyfSM1VUVoMkiRDJnaeMSk7y+ylQd5E318T7jz4uw
YML7eQLLCz0aXvhsTZPvUYgmVhCxJtbCin8khT/obzOZbRIF/nV1nJnVBwFJqzgH
2wcvQq4PbxnAPJ5jomPP9k1GJx21xfd6Q/rXTA4C1HLbjoENiWR7l1T4qGTK6Cy9
ttsLztBmzjnMs3zpiFYdP3itZs/4nEBGkCy2MZRm7vPWFMLGVRk5ae3CFnJIpB6T
JzNnT4S6JsZmr6+JX1Ew//XcCfWwzCXvsPS35kjlEt6ReQT1A84pcadaV2XZ3Gjq
y3zQuo+weZMPOi9EqbGLU90MGrJnucLjGyyW3fXtT8CWhXRpeivpaKG+y1Od/06e
Jxf6qGBTIvXLhonE5Tfbf75sjFbZ5tVeJx1ytEEZKBx0FskytrHBX10VKDql7+eF
ejiFzbSuqnD0l0rCDcFJeHu9p3s3QZjgxQmIlPFAlElG/NlXagLRsFT06qu8f8O5
QlxDXmstPY8AVAkYkDVbK6SUQVlWGvj3OPGNyHb9A1MCnfP0poDwepPe/SsDw6iD
FFJVnmtyu8WTedgWShm10SZygdW9k5s1B6FNYLtlwFLUQflZx9kO+m89DRWbOCkE
Fues6ogF2mtPBjs7yDEvUlDIrBmPRvEFaJXLQNQr9ad2g5P8bzmXGiFxmadQo7nh
eoSQLvUWlASB7gz6A2HWwqcJZcthuZtryeQ0NiDg+s7XkrnLQ6HRPxhiO/7QlS5O
c6md7oyERiHlQAXF3LOUCIJPVEX1HiA3uoZNKBmRgg9iq7x1HpUQN+jQV65KDh9D
B0hALESRkqVdqrrG2Odc+MkC7BJz5fM/4XGZbPy6VSUazUf7pQWA6tKimBpXnfff
3CbTDkv6zI+sp7bbUfKAjIO4OGtVMSBdqhVPxiBD12kDQxCCfNxNWlU3DKpZ4ksF
DhozSX9zOYxmsHk/avvSAhBEanuH5ZNxOIZ8gy7ZJJzzqd2I1lA5W+5vy82iA2iT
iOpS3bBFATAgBp4H7LNP6Uh2/uJheXyloNNUKsVw6Uh+4E0X0P+ijJaDhOdz6LwG
bpWcGQV1vZ4V8qHJlX9PDPfwiZN+/EKZLuuBVqsjjhwlyAGmU+k8cwzogJpykcVI
Apckttc7rFnlo/+Tza0fcWw5n24+7E+PxnD1zgVU5jwA7j+ziO4292aUzV8PHZPk
lnYJau37/p3TE/UtFnPh9doPeXKRcGIwkB0TZSwOToBEMvcxxWUrD3QqXkbO83OV
EMfOg6CvqLzLcv33sTz9G1yzAI4ZXE9uumI4WdkyqOU29t1yD+2OUSmsS8swMdOw
m0Zfl2XJRTi03YVWgfNAMYMh02rUUdMWs0qmOgCMdLsbbqVvLbYaqQm7GJ74lHDK
RUzwePCPUabiCdPjGJLV73ed4lVKh5T+sXHxJOJmV1o=
`pragma protect end_protected
