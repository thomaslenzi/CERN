// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gAFDygF99vMRrdDWbApFHspW6R0jPhDEuM7kZeyH/s7m4V1Sng4HvyLP3jiMCIQY
udeqA5p/Zaft6WXFhGYT6wQoUQmRJmRdW/LTErsIw8vqs2jO/ZhMBHMSaPrabmfq
+d/wKEgZ97sVVdp3RHh3d+08JHvAew5rVAnGe7WJbeA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7504)
wXyaqZusZyMPpOt5yoDzfvM5KmWMBBkIssipgpDWu2lXgjWe+idD2tUGn+X9BM0X
Td5U+DipaPfp/sBYnles4djKaLFMaaaoUNSSr/4sNrFz00zKTDuZddAAKObF2zM1
FIE8WpZF4Gk6i0EKLZRuN1NEzhO0TfMoMxvAbx5YgbwckDI+M88ZqNX6k4wUVByc
5p/HwAinZDiISJBeoyjlIScwNIkXQknlSPyQ8vEuEfbv+jOCnXyfMSilAnQkMf1v
+Cmpt0NLZClyxDvJaocfcHyhPCeippgrFNZt8RjGxjYsf2Bmn0MSopNiePTse9NF
13cNG3v3XFyykDdgFg1a473pzN+/modHgfmhkSjORUYy5MjhhnhllwIgwHSckTpR
yCpsmsWChGQ05HlQpNxFk+R4paPXZ7+jlLFu3t+eny9K1FA29PLfJHVDsPAK/i+y
db9AEVsBd6rxox1cdsVE7jiE509rfJKl03HFpKSmUCr5P94wro+P0+J9oJQsM4uN
QhPz4JNL/FbZbO8uX5PnOOjD1OvGt82GAb8rvAnmZ5EtNJZHThpWWtRYvtxyMCi4
cgy1q99VRj0iutqJ/k+3/JYRk2tOjkJ2rBznSuphkD2Ntr0XodMyv1xw3XHnOp5+
S69HojuJz/9O+kgRi/aIxekjJdQ3ICjLZXRvLGXYwr72dQhG28HQsCxlC7u4x4cx
u1QN+RoYGRcFBoAT99LztlOZUD+672beHV/8VHg6wPFJjVyY3F4NpatK0lvn/nhT
+y2jt77ccUcES5DWuN5QwXId+sIM6VcTfBLcEKmL3F3KnuBm8Ahcv5d8mdtPLnJN
T1p9fDUTIdAj4Ikby5fLAcrfHEWC8HTBdfOkey2lm/0I6EKD7vgHqBb8g8MJMGUo
yTqISQJJfOcDBEtCnQMUJL5lbZWixhDEegShasO72ZQTnuArO87MR2kZYvzv3BSw
Qmp+NK713dZfF2WRtBLaINOmeNpSSzxfcOVzydSfwFLevCSpgDkXvozv1oXP9jx7
dhV5MXeN7dp5kA9m6LzUDeNBTk9rYqngD9guu/smPDWCN4LXVk9eoaPgS+V4h1bg
ZIKfkGyETX2DUgOdZh6fMYaade91xD0IyxXjGzOmGs6J+liQypNluPS/LpcKvC8W
x/ZW97mx0jw1imVFuPg9bvDkW4nPWMJS8uwLGV+P8I+jJrnGcjy7PbdqhWG0bF+Q
f5bPSQp88qHCNtbwiMNQEodBdBXREqjcAheDGfnYtaQjWkMWkZx9WnajnJEYf8HW
IF0n1F+XXgPoUHTPI1+Zpm4vbcETTrJSuNHjJC7hpnKmLTAk5d9C4LrxLPb5RBZE
t+SxLe9MbSosGE/STPXPVccmdrrFonXXdhRB4yfY+NHXmweGS0T79OPSEqilgDDo
5kRNSd1ZhjYguCCZR0e6omr/uLFRcjZEP7QE4DsabOs3bo2FW7uS+/utu/Gtek7U
y1/GvPsDJjzV3xUPdWgT1JaMQkOU8PGqpXYJz67Z6wIFUcLNvZxpg3np9upPOp3E
aAXmbnkQMgo8HMKutXMUbFeOmn5QqhVtW0juiUudwI0jD+i4m09PhdbvFOIEw3UT
sUHbH3N0jVfq37UM7ugLPS7RJsvNQdCsSiVuYxqXsL4T/uxi8MCAUU/CNRiLLI2b
wCYacV2kbV5YSRWoVk3XwVGOpKD0OcKpe4xowxZuknNPnevrv3CKqlpxlYlVTytr
+vSdEa7Sykv37OmjRNJdbqxfwM0W3LCINKvJR+oKJmXpwZx4I6g0j9k2Q+KXk8jM
7BbyzZPPvYiyuT+gM7TnL/3O2uP8sFryGIf0xz80SlHgztOLUCQXNGmhdBF1l2KG
an3uCuv56YGR7fWI7WxH8L+dmix0fmkb78aPyzdezbReangofuzeUKNgec3xm9xl
z0RQ6E9kd3jf3HbsAdQwA+mUQNf0vUOsV4117PF5yEHt8ABNsTTW5U1K9A+cJm4u
c17cfI0MPaisTjgJ2YkIvzEmvSh32okxtXkYegRKMWjUd+ZRQJAy0SqeOfNGT5Wb
t+wOpLq9L6U9YVAUpifIrTdMROU1Ok6RE0YKKr7CMFoPJJICZ3h4rMbZa9t5EfQ0
W8BiTtRoF0xe2K13+A0VSJI7rXqkDRJu7c+WppAyyzuukzd48x7eVupwZEkQPDUn
1EiEk+uNhQ5bF1JRPtMkjeYRJQK0KWnIFdo87PsJ62EQ9T4Y5+AQpaJ4YkMSoNwr
pFX8UrrpAonOvK5xXv+boXA6Ue7hMQRT84HFotxCjNSDSoNbVTqmgMzpCenXgciA
nrwSTsrB6NphYY+aRn0kulWp7z83VtHHZrk6WxRHJGZVm7HId/A7OhjsJDe2QgIv
vnpCzcWvh9tt3Fb/OSFsBzwdz8mCRwrVMsYLFMjvuApxHFko/uLEDqKuIvETf6Wh
cplZ2dYnRm5M0q3ql9x9snfMUHywuvYCnY8ewm+y01Bz2g29rwtrmrsg75FzWxCf
Am6mc7mpBk6+WYn3EiCuM3V878lQgGEoIPVLTiiQb4maLVcYTQ5hoY/okw41M8O/
F3scIG1sx4KqiNB503Tu4BRDAK6/ubZ+Kucofzn5+Dl/gukQPBx2e9Yxj45DQON2
XjnO1GdECS4CuVP2ZFWUy4G2xN5WQk042lazkqmvg8X/toW+eSOm+3uKAVbMZE05
JoxzYUEheSRstJ0yLV7WI8JlrolVqR6Gl0K7dRcUkAsUdpOoQGE7MCfcW451k5/2
xKf8f4MzYtMMQaUaPkoBICsd4/geStG3Z1ESX5QX+o32TryKdC4V31HJB7y4fD6/
YpYhq/35SdIU67dudKP/xJWD8saAUTnH0hYwKVbudDe6gArfkVFVCn8VbhKmqDtW
uO0NkOxm2eILsnsYG4NLx3tmNBKzXqTQgbAWXOpBVdbc98RQK+YU3QGRQKsIMYN2
kcQlAUuI0TevqpMSJjQ+AU2Xgu0cbAvOpnN8+FtiCJ6eSBb+yiYDcMup5DqUo2Xq
d4CPaCKDJs/2VjIAkrEQc1x2/Rb7TigMltM6uqekwhn6lGrCGXEN4+ftT/bv2y+U
G8p8ZYx2ajWLP6b9QUsW+jYWm4JxiMMsdpxgdetUd+1jkajMqxfHJqrerCZsab8j
taFMP8VB1mAoYLm0+srVUz+v1pTJO7jUs9R2rBue0dR9XJSmvSc6KqxEACWbE7cF
/RA3VbDz1HijgpY6Vb74w+Va5S3pvc0VL+q1wa0rF0UGtoSjNb+LLnqwhXPWt0Qf
ZCoJDx2RUrZjlY8Iq9vavX+RokeSqUnAJYGM/oMqtim8bJ+FaMivZJJzKQ5xVjRH
bRJ60C45C1mGzBT+jsJ9yGNZRQzkjsSNLQ859+d4JJs2sBTDsbaJfcT/km7btCac
E4VH6KMqK1w07MNkUsxRNTTxNI9OeoWnrUkBfg0c55OeL0F6eXK2GMeP9ca90rz0
w9U+R9wrxsecAI1yleV9tbUZFDSXo2r8cPSehiCcOJbbU/nYvSRRGB6h3Vn0GyuY
RnDuiFp2SNc1EP8R+H1Po2jydf7moHmiX7c1UG5ikBmemG3uW4TvFXHA1e4w8vBz
jj0bd2x0Sy1dZjYW2Ex6uXruCMfusESYG3YbDN6roKkHET26vLCkWnp9A39GUjVi
ZsRydpZjo6SXkiSVtf/1dQ+wEQSwUiTOh7nZs7xa5+mX7mb6XCD0v5f1FLom2gBh
gPzR3r3x9WhAAbOYJSSXh+UghsInUzsmqSf9G+XNvc5U2J8FQxLftnhiaEbSOUU9
laIMPrcDRk9HQNylqMOlymX19Kp2P2YtuN128+O7lv3Ob0nCn7WmHUyzstYyzk6Y
sqRK8Oxm9o2Y0kW+X+CfIekrJtbWW4ZTsVqJlEGYiRU8gvThK6heMKa75toPjvKB
fKiXdXm8Uvsb249uUqv0fQUzD0Xnt0TeFXfrJmNw6KnthB4N4WWNN/2x6xek4IW0
uT51GASoJljRf88j3BODfZDp+iEkaxT4GUTE7XLGTUqxFEosRBDqhVIatR/kr2NA
KIBrdEQQWrY/oT9U592or4kB7TcRm4on8rdq0ut3cY+h5QBki4MfMK5SiX1WLqPu
Tztl2NKzA/oA1DCOzpQlS0qGpJRqGLjvSKMRlDr/3vPi4SRLYvrpLyd/cL2pboYM
I9b8VK3Qvdvn7/eJRlQ8UwHXV8gtHEq8vFnyi7oN47nkf+mc/rsBldXyeRlQ7e/O
ekeOLTErseiBg3BnuPpd0W3vn86y4SVZqqkcw6fK/Clr90FsUaRQAizO65imp0Cd
M8vyYYCizQ0KwaOFXUyc7Y6reQhtAqNfTEEhOiqQXaar5yCN5ad2wi1vf5dbJQb+
QfANxbttXb9o9xBVyQ3cBvLuHCCEA1FJVu4ocBjafX5M4F9K7WVXplRJ/z9HZ1/P
atezvAPtJgE7zQrNZCv0XbkGFRABx+oXJ4sZSQqZQHPbzg+8F24vXr9+nXDPgfFx
AlD0ZwUcQVx5alZv3ycTSnxW96B7Axc+R4L/m/2jEZoPD7ah9X82+TiIEeSI8iX0
R65yI+nCvXFH/OER58CqeGeQh5aXjyKStAw/phX+3G0uh9s4lybtqiJTI39Iclip
vXVvkV3Unixf/JKnMCbbYSgxB4nRTwH0SNF8k9/K4XOszvT0qnc26u/fFzkHJHBt
RyM0MOk6WyE7Ay9sEvN7BpVRe7SrpM4rpwhA/hU6qPsCnUZZ+fVMX90NsHDhm7Hr
y4WjyvlzTkf9A3MhNLVRO3I4aIkn/L/Goi+fo5u6dibh0USktJNuv5n8Tv0dxe03
AdbDFjUwbIjkRasqQNzoZsUArPIr4YsJbdk9N5ISWrnJzXs8sWgf/f3fiXO/lVf8
OIw2hqIoWfbOqlT47nr391cg/tt74HXeMWQzM/u68VBmV3bveAAY3aJgKPFrbMdO
AuuIBnPiOzLySdIgJRCe7szeQXaVZb6e7KXTYFdbdLf4Kfu2HqPYFMU59Nz9BV7X
oUDxmV33vlfyEJaSdSF+dYgN0HAVKe1ge9v6vXVn9VVpS370UFxqJNhEpSSUjlUN
2NIz2d/sQF0iyHTbyT18yki71aeDaCbPriF7pHD8ypuwBmNLtLeWDzjAZMAILkFp
GZ/53sWWNqn3amdx4kwC58q8Jhi7yE5OpioOlRY6KilHwunFwX6cZgS8DUtv/Olv
Q/uhxGRAG5TNwSRdcyoU5pef2NUC+oJB3WA7+j37pyAghnjF6yIrTa3nCcoV56g1
AqLifNr2Ppi9J6A0i1xY6ge4ebaK3p7NpLcgF4ZrZe5+W+NuyyT1WQSo9Tl1WbsX
DDXo7tt0Qp/qwuedwDUhSppT0oUA9aQLXBeeieelFyCqZOsPq9b2MJu8LxGj6P9I
aSsxLEvgZZpZ42CaLUc7gmi4gSrRTMh5H1zDtb+XyQXlPDWrtRMf/z51g4QfqPYr
sz2GlMCg17JCNnvhoI+l5P2Al4aooiBJHsMkKoFSm6oSRw3/s7Qm52Uj6xrorOpd
5nbAb6S6GB1HY7OCgIhv5RHOl3FzXMzOQ3lJMG5oZBa0Svsi9YPLf34xPA7XueaV
720wxVyd5PINarsY9KKitStuiru1wlRy0j6KADRBYpt2B6VkNWba6pC6cVSxRP7/
5/RkIZ9cy/j1KYr3JbmEUWyHsbXhs80s1gbITzb12LWDjTj/Z9kKBOfx8koLbDEu
lEU99tuTm6FQojVB2kR1BgS4d3L33dY5W4rhs+NjXGZLKxhN7LWjd/e/+Tq0QxoX
Q6gKGMTP9MqlllwV1ZW5+WPI6in7sECcHBAdm9Pmy8LSnC9W/pCGWwlK3PqPi2eu
afDjSi/CRJkRSnsR1yEb4QVAU1N5Y6mUTG99FzEp8zSXzcq9DlFtxp5yLKcM5ux1
UGmhOUhcLqcPJhADUbELaYQIHx+fZ5Cy0upwr6+kGlnRR1qvlzVBaLHxhLaBF3pa
adzcv2lFNds0x7LH4LxvJKxu6EyjGymJxIjwE/s2SzJEmzMcs6fkVW20LgDew1g1
3QAtrOl0Byg6CsA3/VkfetxTdmYRoayKSCoIT/o89ULu9IR9ABN6qeqIkUziFJ2/
wqfkXPH4Iw1Assx1Exgu0CqGrI3MxQ2lITLnyUMI/4btDX0+vnY0//sbsHPUpdv5
QrrmzK953zHQ1Nbg1TT9IIZjOSW9eAolYDpQUeV7DQ5/snuoh8Tl5nwilUV5EPlk
jh+VtWUtNMdR4Y7A5+JbEmJktyg66QqqGUlIvv4NmCTr33xjwYP7NQQ8G+0dxB0K
1oWSp3oxQWCode5cSxxCwdiZ2JWbXu+5EuE8tsIS0AhwThvV9I/VnxtwpvGRH9x4
5364EDB1/r9y5G0AbXGZe5bs1Eupc3Md1KhdeANOoxlTF/kg1XtU7Gfdr/8+faIr
QUtyeV3RXefJzN2WhYc0uLWF68t1sai9Tp7qOvGJ4dqkUGVaTUb5dvwlsi3maxxO
EBffXR71oI+mFQjMZnYEuPRifWJOVugPadn74gWJhCJUUapcV7qW70laWCT92jj9
L0t+bqyLN6snD78mhq8FXmMBo7zEDjUu5pJFOJbcOAo/bfjnGm+ggbIl9+MElECe
xUVMhDJ0FSWyWL5PAiasoQUJIxj09t4XEA4B81I8ZDQndElWacrSmKAQZilqyNCs
2hIOFndSiVaVnJpLlO5R34psTAxhDMPh+HoVPMfXq3cAD42DRsRX0hc2FsrSDs/1
RGhH87H8P0+4GWdyobLQw5DeuSdrUsFOfQCS6cPbaSGjl/fnm5dJoIO7ty131xUe
31dXuUBkfRQtpzvPqBr8PL/orq7+uxY8vgYFkD5YOPD2G1mxvRXLeuE9/c//H4M+
nuaThdrFNtpfm8qSWehedJEWkWrQKjiaij2uNSh4ryjfN9EuhgDf2i3rCwN9FE4G
ZfcNql6W3XNW96XHTFEsN7Ue8DFe2BfYQr+flH3E8MFELQ0mpJdfrlv6yHBZF3zs
v0nbh9XUl6LNAhyxwHCB0qaKDGTBFdHn02P+g1In/3X+ssvctYRi0KtLVSMLtdqR
tG4zKh3Qxkh6v5zzM+3ytjmDqhhDxehKn2LOFJHSIfzu+xfAqyfZfcLQcTMvbWts
KJ+melgIiv9XSVkl7yGSEt9apNxT+tYBFvoRmXQuVY0a0fYDjRWUccjlPPNq6zmP
yW8PmffNupCxEZycouiMK6KkaIQreNOReaRofUryT8btdJ6/VRSiFt14Ao6E/pMY
Nbu6t99xX1ODzFXDHzFsdTUyXxXbsQloYfhaqVdY6IVaHUIlghy0eV/+nib0dWJw
8OsifVy3S5M+RwUvNaxZ33jGzcL33sctjj1KfVZY+0seMwLFBQWuNnMUc/QCQ2wR
8WqWQMgzpvNddLW5VJ3MLhea6OX7J5KkkYndIqxUkn1cRFbOQ4FbRp6KUkJ8ABpo
x6E/IaOVP1aF1S8n2q3pssGmyLkH6fqYHzO1+MYkcmu/dAbMRZFrdLnJhhAfYsq1
u/oNEvRFpNJ2BRNi12WvRRVscBkrSg7mKsHpinhLPPQD2IZrEUYbSIT5FS8KIPcs
aO9OeU3Ft/uemYbYLRm2bYwDgTq0atm7nIS9KPuiv+WdwIEeQd6J+SL1VZzhkQNU
wpKfJzLAVqpUDcCtTSXXQlCU6+dtQG222q3jzeKVLtTYtaUgCO48AQmCtvtJHSsW
pROu4V4H4eOD7ToNKv+hHwq23kbNxGpll/MVUORuMotWOwTI5NHPCa5l2TnppVQG
oE6scnkUzO4MchfbF9G4jd2inf4FITxdzDPEz1prN/h+Fu3xa1aox7jOffK+pNHV
YynSv6kIUW9pF7UzBGL4dGJRiOCLUvsdd37aG7BjrZveyabs+dsmuex3N1WtxVqu
ulYKJrBSeZoQsjL9+rFe/8CyM0abQpZdsHggBX/Z0jp1RItOiGzdqLu/TsB70G9/
ZHx/uAR6g8wXHyUT+FXAPIkeakZYJ1UPJrWCbppd6hzswneOaXUbOxPqWt6JvRXl
YAQbSwH+LbAHv7F/GrYxDR2Frzx3adPH5CXAof5W9uEVGEwiIjufWod6jXwCEfc1
MXh9bkDn6j7kuWEqqbGCt8vlodDqNB0oXAhb9Xlt6UENxY7SE/t/B3lzxyNpVorT
/XPvInOTMdsPaeP7GyFIZWsN4nmiP5h1hfpmmIynoOTiCXbag43R6Je59yU7k4hF
tf3XcgfsdQxy54C6LG1OvlfWVf+9bsWXRKJGkVI1FYd8EAeVf8NQk1IQfe//crW/
7aPhG2SG/8l/gCLAD7mpMWOGmvLR5bcIiSM8BjgwECkN8unnfnq49u1AfGPFg0DO
he2G/l+q8xWENhIMYVdKT3hbaeDfyTJ1UhnyNYPISG7kQxex8gjqOICGNQ2U2E+A
8aeXbJC4QrDO7weKl5mLCy3Jjq33CRtsufeNWrjVehdsyVLOzU6N3xdLV8dLlQTl
NCf/SQudOy8W/hH3JjYad3dpzGllFkwgi/XExxhebkBnuSyvJlcFU8HZJklrgECq
+7XdxM4uAs4g5yVJ1egRBcLj4MUnHe+aSBxWTjks4mXoy9mlXZqbMIm/9jdsnc8d
Lp44rRHiv+o4ou+4vOTFTbLzTdPiC5qYMlBgbpkBmJpZZGd36VbPBJDBxNre0Ko9
1e0tlVLPL/rLGN1vLmhXZUWfFLy3JP3Mdz77qt/vrU4v71RqN8YYipzjspLej1Nk
d+RH/ruGYzgIdZk92vUhg2X3eeOcnw6UeMP9fXS8TzudGN5hMwW7m7Eqji4z6fZp
y6l0SerlqQ2OX3icTqgtIf354LG5wrKqHxXdUS4zD758wPahNe+/GVcBIM5TQtpy
Gl0+K+WSRIyTYO1P5knAWdUshdvcXboRzR4xhV0RkbYB3dNvIROXHhnb91jCLA4L
PioOZzcqWfOFCK3QE6p4qGWHLjZj/88BE+/PLh2mPu/QM5YVcxmb2Z6tG2EM18om
fjLqcz3za0/GZl3G8w/4/JuwxM5RCat31B/L8abyNtpCV9+nJ3M/cDmBn37G5ayA
ZHH/AwQd6EFMJe66Synke/Tfhy1+ja0umq2WSDaPfvj7jllz/H7XCTHGnJVPCHGn
1YY4yqrV5ChObsrsWHOG+PPOT7EcaNqZ1wB9Ch/SSUqwBSJwChxW3k8aXhCdlN8V
rQZ32zM2BV8nb1Uq3NtZ9Wboh/45PI8PX+K3ZuTTe2/5tV5LSHzZSEdTMp+BPc1B
7UrvVp/9AYlzUgfB9g3NVKbOnzo6sQdm65Mh5EZDICSRWIhtpVJPsA5/+rzZdOAE
m7zRCeDzd/WQmAEb5TmQPyMUAEJFSej80oOILudz2vZhQMoYeU0hTZC/saXT6ZQf
sfnvSPROHYcrtYX0LVAfYctYfS4FGKhYMUMdB/8TbCruQvjsne2tAY5RyPqZjdpC
vSgmRCpZfNdP94pWwxb2A8mzYTsvCF6GKPI1/qVd/8Q7owxFP19LUgtta/gx3o0o
FOejVj/OLs4yahPhXO5RZyyNn7nH/siYJE7UHKtO8DKicpyuWXFl3B+cuhPqOjEa
7KvZ3TyVbO/wvzEliL6sX3Ecjnzk7yDaNUUH6F9oNT1zGBFPjxBK56JhCyjPomS7
QQZIgbisn82lKAju5CoWfaqUZkr+FR+8LGx/wEouR1mhAAN68mzSuvSlOAVDE7x8
UAF8KjJikTeLy0Ox9tb+hk8qVpTq0wvDbxQH/uc7OeOFTwI/ocvOeCsU4lD1RwTD
yYpNAI94KGMQFQWxM+qS8MgEFQzKRP9Jpt5NcqThvj1PVjiH+FWSgjWnQOoAJ2Ly
a0+V6pV5zsKFvv2Z9WQkCf6LLQ5duM2Sm+yf9Xp/XczSOgFM0RojiG5yV3RDNZCG
SXItgg0yIdEnnexS3EoQm0iU1sNbrZ12DC8zCPiNgt45DZ4CvioMd9JW2Qpujdkb
6f465CEfzBlKBXPNEKsMDaxbledo6fb5CQRhuOYUw4FXz8LZCyZ6IM6+n+vqvbbV
AlesiZCBb+Idef+DwHBLtg==
`pragma protect end_protected
