// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GWNhR7gKbLb8OMXxanF3nDJ3nX4tpz+99+5bW/DuQFH2u9A8b5kXyB2PlK7D0ajh
6gjo4U5G3LjUuEIxk8fYHS4V5vWfC2LmuNqbKiP/9mXcpQtEMGmRMmVr4krOwx2Z
NaOM9GB3sUnbRllV+XaE0TOJffRDkbh/f97tQaLrBJQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30576)
7tmUMRt6a3bMWxnvKbNHBdAe1VT5dh+xCKBEB+8z1+yDv3dMFl3oVXrzga56dWxF
lMpd+lxA7iFXa1j/SrQKnXB9U1ty3/1w08hyE2uUv7T7ruqshC5QGky864I38rZ3
KhpteUTXmm7+OOlNf2bu0kkXfhVjUREshANJltqB1wKDqsmd/ENJhrldYFHwBoSX
tEMGga1wRy1CKOiUQl9hYOJ7WZymKf+UZK1r1dKC9660s7PDimVXMdg0SfEK3XVF
S6WaeXqS4QX7YRDJ0Ji4bY3qRMvibXW5xdQONiCP/P8LFv/dsjn8TuyzjAfPPdUS
MgtxCn0JBHH9oufmYI+9SceJR7xDBnbmLHXLRSI1Qdv/Ksc4Kgp0G735vOHFk8tH
TZa1edxl/6LA+g93TpjGqBuFeTjyxVBVO/t8zw2VmDAesiMWomYnJq5vO0O7RPJb
Cro+2N3vtmsvmc7A8b78l3EEV8dNo/lhloROLPL31hFVwGCVHRSsju2f/w0j2InL
KeizxOmwc/92Y71MoxLOYzXAtyimppLV4pkAkZiNE/Rr50l5oYOCY64cnuE3MfiO
ZXQNs+eMzJV/teoerLPRyKBxq6bzGBa9GFPXAxKVDa5SItHJjqZEbLjieuHU/TwD
0gOn+kL86xMwwFMi8pXr7I5j4mdwlaPEcec/o13bZDsuAcetXhyv7yOfmBvd9MdI
D9GJQnFznQGPb3/Z2IAViwM5L+rR+Fan/MeKJ2wlZpIxJhfhjLBU6VZ17zv8dGQ0
1kn/XjevrKIfQ70tIG83gQnuL74/g2qk8OO1rlW2EfYmFO5QGkDGcdAyJKkS8VA4
6BQWHdeKHQPI59PejujsVo/VAvsYRXQvKhNz1UCdHmd3mn0+aDOYKfHFGKINjdJ+
ghn54wt+JZGJtxLHxdtT+fPvVRe31Sq7LPN+6sHI4Hh+sOLP/9R/05H+z5l6X0B0
k8H9IrIYKjos+GCoSEYnc+mk9+i6e6YqRYWpIXUStSNpaDnUykwf6AaUyxNu672u
lGwB/zcNtQI4PukuXX6Ht9TjjKNUI/3as7dW8+NkCPKqxFlBWwlRA/2r54QA8Wg1
Ve8WMNCmxXtiEADZX/O1i0f2ju/UHJT1m3EPSxbyQxUcHQ40/Fhy1/oAvdrhKcF4
KUPGsBGxyAp7Z6q0ZOXsc10tZT0Ux4Vp9W0GML59V67vWyiNBVIeE/rGQqJXKutD
sgLZvJe3A0KoO9yxo/OwExOEHBL+wwL+2X6lNipaGOkFiD9lTiTUNHQYbrEeB5+k
HiVEKvX+onwsYjvfdGdf3BeCnXz37TKbYNtbrEyd9jQqNP608YADQL5N6qw/2EyY
q+rZo7PGl6N6k9SXdhnBFY+ROVLnpVF6gTRKf1RZ/XmzB2+FB7wTUzA0BR8d92aI
8wq/+HVIdyevai2E73eUoWOc0AOxl8bUzZ3Qz6Jl26jdS1ooAY9tVqc4u9BemODG
nQ1ME0QJ4UGEFOzwVhkAHI81QD/vVjpp2X5PzmR1BOLi3EI6uegrI7p/e1gECpPf
LGGevhlLYrDIuELxF6srko6nLMwRbHKvn4g2EKOdB5F/dbIN7TyHEqpFsD33mfVD
KrDmn1bpJyuczi07deffwDIuWbitxRW4yIOp8WByZ2MDVOG/5+HKCdozyPEYQYOE
jmFRtGQqTGjGZrm/cZ6efkCtXfrJhuY8FafO2OnRXLYtsviKScB5EGVfT5Qu2Qrn
s2uctuhRTXbgYu6NoSipq+yG5khfxTpHWTez30wngdV+HK6nJ4nrR2mHRb7QelXM
HLfo7U9kD9Icwhd6RzSCiWgtDH1x9Pt0y9MlUqFrz99WhgdnRMYh/mryAGAwvK9a
wieAHtmzd/YYz0NKeB6o2feAMDpdALGxoqIeIM0b/w92fn/RNxFF2l5rT147b0wU
dk62wGU/rcbcRrwLMazrMmgQ1WKCL+I5C13/fwYammFBkq0ylAIpqMIIZWJkzqkF
F/kbcju20dtP960txs1V6HMBx56WzpN/YcdDMVamkMHpoV9vMWmAUw2RnOBQrAcx
4jrnnoTVyz0Pw5fSDJ4C6aadCmVgtEjlycWHQrRwCPym89qi5S46oGuw4L15HpA8
akpI0EugOotcPF7Axm1fQD32O1xGImK/4CBxkZGFi2nilJl+RG/+3t0VTWGsw0IS
zfC0Y6j+zo0jTZACx7RmrMimJDuOi+deJWDYGf/KybrQHWEVlwYp37CK1xKAyicd
SdPY2UkXSRQEk2XBVB0tN+YIBa1EFmK4a37LT/9h6KYusRediXfWGtuzVpESvclT
nDvMPgZ9WjLW546hCFId5Lp7QOSgJljvuXpsJ3JFyKvv2RqS/aovhL2jUHMn3N6W
hvvSXxtL15kQ2gCdGNLLaiFwR/bLmiAq46RjvW1wn62xsztiqHf54p+P8/whxsAy
uvsu6oFY9HCs8lQee3XsuFIo0KekfOpEgnOWrA2aQ9ukTJiwfcCl9hacX5A3opNN
GOyUQyU+qNv7GwGYoEEJr2r0vMFlpdQd5Vwwem5w6X7BfAOKUjo/SJrHCptSFoPv
t9qnYAoj0NEICUtQD4W5AVEEuiT1RQ9CLRHt7Fft2ht0CLt/Gxhx8jiEGQkfJ625
QSD11l81/JUGCJXwMZG7P5RNmpufWXix+pN0TneNiaAnVfTZJOSjVS5Qus8Ym8qW
p7TSDg8muu4uXxbVyyE6UHuPqV+5wPOW03PJ5BZO2KSJ3DDKSq+bS5PZSdxgPhmA
DUIYFiFvKOX6ycnklKvPK1DbmgL8k/nxWlmgXr+COKxzlkpUM0PzHD/LF5WSOfCN
DwufGc9R6jAGPU1Vmrs3K68ih/f1cLjBFhH/+QmW8naFK7KRiNrQ2ny4TxQ75JK6
O7RSAEwMsoFwQVvzuFvk/Vpfw/tIg/mbjCUr/VvMKwD0e/TVOslAaX6opjFvTouX
N0vWdXDedbHNoeTCoZ9JpfJkKuYbjQJkkABpWV3m366oQ5e4eXrLvPEIxVoSRU8j
vs9218388/ytyBs93THcPC1cTcfNO37DslfclzpVCI0UbP+nfuD1FUeZ6uJtBW/r
fuAm3iUnHyWsx+Q4LyL2XO1QG932+Gz1blfsFupi9F9g93ZWxFlUXRZ3sVghEtgN
kVAOmGXbszIM3X58kPB989SJbQcR+oV+Ieb1SwwLEsxo8NPJ6TlAt/6D6qhU6alW
qh1Fe3xmFInKsmeRlkWGHMP2oGzyJsCqJEbqVoXbHCIVSZ4QueAtAHt4ct3dPmyF
IA8o2E5ueFiLQ5Wm9V3dixV40+uaM0Z6ZR3N9eWpnuuvsuwLJJFOdPxFKOlfNPtF
wKOy/K3oie4+cWH+zmztdLBMpKMYEIf1Zj+wJDtnp4hzcf9v3BOn/l6PHzLpUoPX
5NGDG19cwmTW1zJvxQD8Zci+Hdq0eB/6aMfExIWCzep/lz+0QSQHRMdqB+GODP1f
Cfxi3ad1RSLOVt6IrqeWv3Cb/JVYVPTgerc4qnewuuie9iNo19TVIbFIcdJjzxZt
zXiAWbpNwV0rzkI8JLKtlIh6EpF9mrdElBYFp9zPfOtyh3BWqp0uA/eQB2POUaHf
004cxF87YuhDdv3GfTbkkCLxYGVDW7Rk6R88lOjxl0GK7iIfu3/+nctC25eTN0jE
D3x27T51jUK489gcppRIos85dldrjzvH1L0JXiT0TIQaEUGYePPFhDgBtbrdlvDU
y2aHMZECnWAyf354XiZmsHcBPXNs5fWAkpShjSIz/zw1CntweRY1cDYov3QGTVW1
TmaX1zXy6iqUsyP68EOQCHK1DZkd8QaqkClvLgG7Zsfl45to6DyrpEdPAm+IOopH
jVtfrA+0Ob4n63po5cz5zfx9rzoJhzW8sNf13Cmgn80m1BOUmiT/twyilJqb63cV
dJtHVe6eO3KxItoTIuxLBdkNz9p/IkJ564Yd5gQut0zluWLhTLQCufpVZEcQ5Slj
sOFiv8LK7Jf9hQ7oHNyxNRd7kTByRrnq4wdb3HWol+G+UW1fOvlK7/YcPGJzyw+B
FkskLjhWYGqqe4uTXsx6DyICnUfopeVIBGyvf3AcgjIKF5BRAwnQRS97FgQN/qMc
sXZl5ICivhLYnWlbSOpBLueNYPGF8WSAxxhL1hrl+m71Rj5M9ck9uHCq0AG13qI5
MqGwmFQtta1PtsDIY1cMf8bmT5aY5NCWVjeUJTztGwDPf7OW1AJ77Ys96i/KH0Im
bqTg4S5uaAeXk4PqKmnzuD1qwYTQFKTrvxSHfLGMNR6Ul3m5FpV8xzmBT0icVBIw
zbHg2ADSgkOQ1j+xBdASvfcJu3ZJbKPDHtZPsFxpyh7AfUAkD1+ssgmceCNxa9gp
I41QzsX30KqdGg/iuXuO5RubdU8VthzRqOdPyco+fzCw/v1DZK12O1ypZ6a5VPBt
fTl2VVaxI506LECvWYn0ofZ3rs+1teWSMzSfHjCKoA0ryrJifeA0uxG6he5p8AcZ
L3NWnBh00TN1hnLnA/lI3gqHqylZx0f+XR+HqdXne1xJlOXAYoPdTHoiWxFwZMHx
FN6zKiLdUionqJ5xLgkV6JnVMVm7Ai8YLjf857anpypD2qTIRge3miPWVnXX6PY8
c9WOYQMXvsDQGCH76bMlotZ7HOcsglsFRBzWUVXch48AzEyGcsD4blR1iZMwP67M
PH21A9xlSJ1rWiAJ6NDs2Tq7ZWj0sFM39TN1qzXKFWNuig/1OGcpas/boGygQLQF
tYltbEPQswf0i+k79NUlLbLJE7E8WiDYmzYyBj6coIY3mrsq6PSy0neTIBonHH+K
Qg+FYyrkX058niUsVrQQdzWUe5BPzCGw9m5Sd/JlSCERMToUujgXUyNCg1Y6kT65
Y4OR7TOTvbuPoRuc5S0/GALrKGSNaJPH9B6U49dbaiDUe2yXGRqH6qMR5gezQ0E/
+PIunmHzbd5o0gautBtkTipE7W26giIhyvZNzKIJtYWua8hfe6GAzITMLShjc8ac
Cm4fA0cm5UlVBkjvdALDlLFCCgaZsk63B/kjTMpk/S56QUyj4UX1ERuhtN32N0xM
GZQgOKb+LBwFErPn6NQ81R3OXRvNLNmNtmeOd2n8+1mmfOjNxF6Z0urJG7ingl7n
VOw4rxAeuPEJgiYXOjz6AAI2niO6zUppzNvCSj5olLc2x7X/xXlqFqZ1a1z2HRxK
T8QDYSzlNKn69szcRgpxBq7kL5kbHTJmpE5wEHxMb9zcy4/GESS3tlkO+ljQ6ZlE
eaNIv3kwAS/RMf2DqhJRVPMn12PCzBEG6IZDQBHgaiKjwowD74kFKdH2JI24B3d7
SFu6Fs9e8QCGFlouLN42J/fET9Eka92DM5gtReutB7oGQCDuC6ALwXKe+YpalqQc
+NS9pobugO/7JHZZQTjNEhYZPvNgkfuq8LZWXo7/3W6oUAO51Ke8CcbGU//uZtWj
h2M1w8e3eQxuSzq7phTe7F224wMJ1vgS73D2TssvMAuJLHh0yMhRxwEl5dEOXT4E
AttasgeLLtLyDzoQ8kARQj5YyEOmglPk3CzwoD1ipXEDeR0B9l1WxtHb9HqnJ+sx
gm3sgvpHpHnIeGeqOfvOsOcdb158cNNtXlUMpfv+lYcHHdH5cv/ALBVOOU4z+TzH
NUtUSnFGoA45KwtT5YIcdK1K19PiDREwqJZ4WMkJiW1bTFUxMYjAHVXmL9JgwvOW
jkpqgqwSEJ/z8NXXieQH4hrluFb3xKlhCtHgQFEy/rNpfYFjgxjSzFBwoMH4JfWh
EEH5JX2D1+vlc37MffJNVZfyQaBUcD44WMPEw9mRtUJaglR/hzgAV0eI2Ubw8DNr
zkUPveE518dZ1lSUpthWwNdYs/9SKQk8Q5zVmrRkNTapHWEA6xl6HazYk6y9lmE2
0ExELtlQ0lWXKV3u3OC8OFrQgVOGQjYc7hyE8EX9t+fjvxBRXZLxXYeo24G61V//
HLCI0Z/GCV7pG+Wc/4Gz7OytB/giZJL74SDPeZu4h4V3jwAyipASPd1C0hf0i6zE
3tUd7J2xw2yStVHHqOPPAqUW515XOaLom+dYUkhht4BbS2jUTZyl/fCoDXBmEka3
mk2/b7XtqN26txF1qFAM22yNzFliO1TvKsIqufwrwgvFU+oGSruQdz6hLWWmSp93
Ngxt5n9HYt1CKTcmAZjs1oRUN8NLVol5RPXdA0/IoapDGrUK0wwbG/2oWTQNhM20
Yvmp3DwRG+N/4g/zV3NjIDbAw4IMNMp342NpFW8Jpr9C7gTr6X5C0zHzPuxBCiHJ
fWvjpMnhsbFJi3fjXL/qZKtlkt53pZ+/uDmR4JEPgJV5N4GbxmrY/nDtN2ApKRDZ
jvjgEeLLkuI6AXGjVgVqUhOf5LPEMdAYxEPCeH4xwIS7+Mgmnziiz7Gdc47vrOOb
AOjNSz3tbf9hxg95XUCC5EKmAmzzq1hIxLjCW6PzO0OWpyUnw1ZX+SUsL+nf7gv+
opPkl8aBsIKis9k/HpXJ0raEdYNGBTsPSr3MxMP/x7IiAABuOeewZbGwaOlDOGMG
JkBIgv/cD8Ou/aW4PjSyyTqK7z+9wvtSJc0nT4HECHJCX6CVXa7lW6iWm0iSRGUz
zeXwf4DtqSJ+9TU91P+Hd1quKffpP1V2R5dmoFIVspHlty35KblUalbKiGMXy6DN
MEucS7SUxUfPc8reuCIQxLTZUSUFlvMy3P/p/3G1ejF1Qcx9yVq4TlN/E6mkTkEk
lckUWoySULKBv19xoFR+MBFVEcoiUE901zz06AsJWJzzi1nwYzz0VuV6kewq4RTt
keEfVZ88YpLofxwOybArbyF27PpjZ0nfYd4f8kdaQbi52YNtLsJCERq6XGTWMUJT
W38ThY5iRpj2VutuyBlPmXiTvg+nkFX3434R67cZ1Y/YHUpcoOJNSTQKaC76NYe5
4HEKSif/AR/laz4ofKAk2f9PhQjk3kjEy8NsQ+NSvzAy2JOgvjs70P1+upedggT/
1iRcH2vpkC5jYH1IocZU6tZqCMGdt1SgirhmYjrhBBD5XvD4iIAUSDZMpOCmpuv/
h1ZHkXIrKI83xXoFQ4cOkPc3hHP02P05+kFNDsTTj4lKU96eycqoBVLyQvb8gLyH
PwDah0uN0NNH/4TJMLftj3jqHX2D+LB5amcAV7EPBqFebZW2vDVcR8amxl0LU2wb
K97WxaAzjMINHetlSylG3H/2l5zHzHSKXOtKkKjXJbyxdOsOcYRtz7QE6mSSX5L0
7Nl3/qR6zR8/GtdkJ1Q2SUfdJo5lgOvmzpdrUTnOpsv9m93QfrVliAE/A6oOA2vM
Mu9m+ibQ1omZFccjQ/9RLrDEXMwtAxx5USeWJWOYKxxRqzQYOQCT7gP9/bDipAkr
tB8FZn6BUFG8DZhiwrUda8CXjADtnTm6MRVA+4/keHwiU8rpx2NoC07ZrpCYaQDu
7fDUj6+Li0BinJW6eX/IwYINrt1fhGwM3WF8cO1JKJoBSu7tWht5X0I6yjPvQOcw
7AjV2YtB2Qln1ZUzZdjqoElsLb5PXC8p8Eh9pnSuu2Oa1zoaaW5gkVGgvD3SWLNL
4Ug8acGPqRkGX7o4oikvuEbNk67vEAs9F8cwZavyCOnaP5BymT5iv9PX8TSKZ1Rs
6MDMjv4XSYeaeqmI/ihLJ2ze2HLar3qXsdsuvJzkZUwHfCkGPme2UVw163C0iC+q
3e8xayVLd86/XKSRWuwhHdncknrKE/XyN901uz8pdI7gZf4DXbYjQV1Mm9Y5O7rU
dR0DuiH4hIzZaANZcXl7aNgHO4o3pJZzTzHAnWLsl4utQULWSQqOjOolWyp3f2tL
15sKYfPw/BSm6sJ6TWJaKg0G1LqSs3wuiseJkMemYoY3ttB+Vbdua1zlvv/4DA8c
kUnTxVHBFTKnoIzA2PiKkjFuO9jTa5p2tAGeWW2dJqWFKkLPoK+hnQEPsW//H/jh
A0YgL3+78g4pRCmos6OG3rxmdG8879A1QgbqfOQKaaJ1fAH+NDZye2YEUun2MYPh
RRI73HqPyCZoWAUx12i82p0jaajBxrHVM3zuKDtYaAVb6e+Dk/nfbEfGU2yJpq8J
k/rt81E+FerIXIajFmsFU/c1L2VW78b3iSNI2xRO7t8dUmKfUwnA8ccEtZey8Yu0
AHJgTUBuWSnSGN7YY1gIFPJLwrjTdG6LhI21WI33v1qoO6CfKoRdtnxOAnl+4UGV
ZRXIS1nSvmRNRttiIfS9g1UkoA4QhPHlyAijqkDqY6iOMz9jb/GGmc2Y8UbPTtqw
o+zJeVo6ynrYbXqfzb6kRWquu47dvew4Dp7iUUHUyJpu6mHNx5JMFrZNU0H4lNJi
jldmUjs39zFD09eCS+Ol5khRCtNLhBWZzoAD84aoVtT9hfOl91oJH9U3kG7BWRsy
1WBEcDEeq0Ta8HdUjv7NWPRP2boEaaJ5gviXvVpJ6yEAkTf9k9YHoLTzfVeIQAlX
xUS3Ep00WDk/BM2QLh9cZLda2McTt6TRmmBTKzq7xtoPzHhCgLAlEZvzlEcO9U86
+Q3GMvyaJEVJs83hUaHK/0A2MQVeNVi4BsP36J/nydWAk3vEcC0GEh3WwGToHjkf
ZA2aiijwVveUOA4+GUzHs6wMiJ+TRIqQuEtTL7wPDh9MkUMXvR/HrIX4HflWNUH+
RyQvLWs0oFtYD+850+0UHTJji63XO0fCP6gJYy8/O5a5H//hKweQj1+4vkw++U4I
aphda7iM7iDWQWsANLNiPpufhu3elMDm5kY4rLK49ajGtVlo0JqOU/5tr7J3Kbi9
IUGUMmFPJnDBuv1PYhAJVoDVGfS6oHkejLkBaTXgrfMya418Cx8FEjETe7uWpLG0
HShImdOt4ThO52sXowJy10q6lfUeKHba/bYdEouG/XxMkESISJKFCEnIfk2HQuoP
pl0yFh655wVIUtl5GRcv1VAtQh4ixCs2z9Lfc5+CS9SahY1bML10gRyv8Tr0SyX1
MsEXueFKkXipIvEKqZAD2v3xOjEwqd5iTUbxpfErSQn7oHQsRbYtk3Mz8tq3LLOf
OpSFgAiUStNrJY2IlGwilNuELs8zplUg6TnWbu3kUwIqQYKfM1uf84kSDQzoB1NQ
o3W18AY8pucLGCHkq30P+z6AlzqiSqPEgE7gpP1MG3MepPf4nbB/nYNhFqtnpF4H
yooj71Np2Gvu/ldHkk5xv3IKrYcQEx9JdDCj31NOKs9cDhPV+QQ9KMVQ/Z+fSeSp
VNYU4E5sOHU3gLqkFdtOgsQYXydtjSJHJAM+Q7rlqDWpVy9tLDO/utEhtWy1DY+4
ADDQs+7IkbuTMNsVzIa/onmtEZrZoNekvvBUzvEX3nGeXM3znQDiVhS6QwmQRK5X
coaDaXUzvZGzaiWio6pFxTWb42xXTz7cF8nhTfwHBRGq1Vhc/fpvsNhjRObNXomE
OVSbfhcNJLTqQEVmjlAOZdbOffoXHfE2XAVLu7Lcc5/C7uiKYLIKWT0n5V08PA2M
urX3YWN2EFLP77RwaFzB9e6h74pDzraB5Gd3d2ToZ78Uk0302AeIW5ldCRMXCc7M
izgqMuKbrku5Etq3q57RX8zLBDxY3fT1z/NlQ55EJeXzhYwNkcmNjiOuR0el0xbd
spoMgoy6YlFP9URLJWeDqDpttwlfavhkf18BN3KI15Gkq+M4A5DTkTLVesoa8Gfi
TY00W3W6yQW9RYxQhtCuLOD9eyHgThs2F2Kol67lcdwjE26oQ0TY0RqsgW+OC/dw
C0e2bNT4M95YVFkWvJc2Aty0ZJHNiUY7pAjoPzYrRBdp+PX4ry7fh65T0DrQpN9p
612c+H5KBTzrZDAYZR4F7D2SociMd4pWqPJ1QkBA2hffLZzNsJ4omOcgC+gtdSmX
zDSwsm5YGczbmdA4kwczqfcLpYSqIEQKWFYXoqH6ey1V+X+z5kO1vAcw48Vj4AaC
gqGEPorXZVRLc1sAote1iB2thD6nwYuGBBzIDmIlWObhM092Rn43LtJF4pCeLPkA
8BDx0eeOe0SQ5kV96nv9PYTXhwjo4HXUAFa23ogAsy5s4v7tNaoZ7R0qKxq8B9U3
kJr9GU1f8DTJQRvsN2BmUint9KN7ZCBOc+OGWOfcH3nztIvOYxfDfqYnl6bXfqji
slM93FMCE7/lqxu3Y8+yycPrZwt6cWOQY2EzriINpRjMecd5DyN4eMQhkxt4U5G2
cwosulXwXCjbstoBdSYmecuZ5y0uUnuioqj0k27RMCuh31SZau/rdIbr5z6Y4qZk
Q15pf573svqoXQzSF2bD6blKRMP0CFjlSPI4n/CmNFI5rYO7v1d9iyS4TA0jrAHz
3P72MCv1+eyKLyshEFk1jFRtdB8kMa2oTtdZeyrKFPC4Wdj9T9UXPXQH/+IsA6Wr
UmZEFvVKyHYfV/KtDgCTEnS+en5B4drxI2RKkv60goYbNZvmdr5l81QL7q56vf2H
4gtFPaCtQdYR9ePYGLfJnpInYMCXE5mxL4wqgOy0VnLIMKYUdlOCT4t3R0t7LINp
GsxJQ6N1KTfPPQbrUdZRG4zavfjtK1msNLrlIjbzrNoopK8tu6p7vVs1YzpsHVi8
/VSZdQc7dKIQPV9Jq2QXXo7NpmozYvp7wxXc6xo/NixDBU97fOcK16e+qZKQQkqi
41VIVyhAI+JBP0FwnI7rZcAC8Rsyt35TppwtxJaB4T29ESFKso4dUHctDh+Mucrb
DKa3R5OGg0qX/MStpMSJm2assnmE+wLwV2r04Y2BQgDpHKDVANodSVeKHQfwAz6+
oX0T6xoJTEfwZzCJSomjAhKogrVccNtGv6okkFhTE9c8Xmw4o4mO0lVVNjHhPFKs
TQxaduQUCpnE+LAOodGo7gM+RY24PQSKY2EECLVLkF6SxJDPMmP/k9JNM5a4dx1t
rJeLRQdtFIbgWLN7LRbUzbbMclWjOaM9HsvOsaZoH3AxzyUv0mOotpp7KsM0iQEK
uAJ7K3vkuSpZkDgx8x7dytS7by3T/KQJvPjlcxaI1U2/EKz8C/SiPfdTSDKk9jWi
Ayy4XpgI9ZZEMFNQc5u65sw4d/uYO/gnOy4gaiH7sG0IPA+JUSeMChVZS4H2YAAT
IiF1/Y42Qm7eu7PjjgAO4k16xwvjrr57eyrkAtHPM51ma4WrerGEZ/A3TU3UZsO7
dL4ZTxnMB6oVtNeIrK4FJ/2ySn0I9Wp5pslrARsYUuFLPYS3JEBe1AUicpUgK7mm
HCkCHwLkZnxbA/fCb3ZHzmtbUZC9U2343QfT5LemP4cZVpzoDYWrlbBWgh+dRUGv
0ymf0aYRuzFMECs1NLhW4/eKtToHOA+W6vuwkxCHHEm4yJV83N9adjh9nOYH0Z+I
x/0oef4odq0yiVk2DTWOYx7kMP/fxJkrurMlJxBtYQZu/1CsF7/dR5ZEcQbqu5B7
M/erBHXNkHGZMp9Ia9HxAiefAj8fmOmyOWG+lnW3VxjjtStPB85iidqmsfef0uH2
VUsX0tUY+4sspG/N8Hfrfz10yj6kzggAwk7RYFNlbl4QPJE5b+mkG2seIDTE2cNg
CGkFi8WNNeNmbPM82kvcKCPfhMC1btWMhrvgq1MF47dFht9Yx8f3LqZc/fknk/Qz
PvXfb3KPuW3Mqp5WA/E7NCfVKnYL3zQNwALeVCfzvAW88kdXvDT4LeSYZzimGQZa
hsjd7d8edCfclRoHOHWcgaiv/dBPOZhSqQqpazlyLOpSle3sHfsYcxADz9oheI1Z
jiPpdkP02+Aew1nRq0a8uBtPD9UFVB7wXsQbflyBqkpA2He2e9GroqJn8/k2FYKv
UVFl0lw9WlrB/MMMU3Yyhe2vP0cEEc7BLfgoJdE2i+b3ZiynH+CjM4bg+lEifXhg
KhDv65+TN5Es2zyiqjzCcejMWDHM3x/jSkX7fkbKae4CN6mWph2EAVA2G4Ar1VE8
i5/hg3+XrHPIIyptpDn1E837OxBvcllmUnFiEA6MkBWnZIBrMJz2MAAZfHClo3Yc
TBk1AoneBKQBgdIGEkW1N1kB0Zr44gtLIDsJVGtiCUAQbEwkrh1ko6dYylJsVshJ
1nQotv22MfERT/v+eqEQbnCmmJYcEfUYN1aVG4i49oISYhBBUjNoml+m60idxBjB
2Z1TiqN3Zw8X2ajeWYzlN3lr1cVGUFJn231tbbHjuSYMxrgo7QXyhrU1SHXF4WpY
niD8cEFDn13A/FrUp4b8+jNoPB6Ta7pAoqTIMRqc2waxwODi51kzw3ajzWfKIiZG
bh/rL0hnVhS2PMV9CyOcuYTU8BGRF3tWaRBwMDhKJ62vgnWFD0dHuUuVBOGHM6Hh
cR74f/0pcJZnbs7avWUdccQo/TtgoRmKeov7Sz+wQuZUcS2l4volsDTWVPGSA2Fd
QvYotA8oOcgfXxUgsqjtRCQaqGk5rHDgGMrR074yLZ++qpmCn44qi8iuvBEyDD0R
4AvXipt7DVhUM5X1FjT6E1vNPbKTue7nig+1vTtrllLomFt6KF5EVIHwmesB//fB
H0PpdRogMDMq05lvrRMQCdjotGI0zO+bGNCtg97syCO4V2Od/faSERbtBrigBTDv
fyDlz1jR3sRJEHu5FxUXud+62VLzUIieIGQleP1aU1ymEefRnwlJygcAgNuvfuSO
xCgHgD0BILLnMrhFV2nHAlRT7WQBlj7cTCb3KLh1VErjiPXPO/rzEy0h26giJ8ov
nliFY11msDwnbzkwWfKHq4a3U8Dg4dMa8OCTVDz4D28twME6PTqDDvTXs+xwHMqL
2KT/jwaTi1RU1MG0AHXthuOjxPcb7BqD6wdnw9DFdJAAhvrrVJ2blqMhWFpXybO/
5MbQ4WfKaihR2pECsWrwjzKjd6KIRvOy8Hh83BZJaxTKSjbQgkDIOUpuTIAkP/29
jTI5kQScplXUsF2qj4qb9N4MR+3BdZHDntWuB0UhsbooE64k4obOr5DQlFD0FaR7
AvKI0ndaFAkIZPYVQL8N0l1RddLkw28kXHr5z9Dfcy6+TAKaIKpN1K6vBh+snUDu
Gn77NOXr0Wf6/s8N1nzvwWv4nq611qZmS068qy11oYIUU+JFPJy0pTsFFZCRrB4Y
oCkHyR6ktkWBF6UvCljNqS5ryYy7tZf91BG1e0OLbqH0omDVJd/0xeUs5hqCIAOF
EvPS1TCmlQz5necK+cEijZ2nCtsSPBBCOBPP1B1AXwdVKi8vbQTyxKCPWcLQGK/D
cK/9wTjYo/gu0rmtM2G93vVLZT+RT24WdigrOAyd2EWMvpDmUuP/P7quLquLY6gc
ZF67Z7UU4+o2sq7h8VKEdSwSMFLmboDhyqzcWmMs+tR2me0SyVCxLz9bI4jj2Dd0
r3D6/jzvN7nS76kWWT2SPxDT5AQib6uT1WcVQDcvLDPCo1/jpeOGuToRfYPsi1Z2
ujG3liMATlchtF/Ltatd2kNWfqSmwiT2zohB0edePA903z5vuptBW4BF7SX4eLl/
M9hcZYgqbyKoKCYUkD72/e3CtEQT5TCwJ6FpjR3/mSASx12CwANG3BkaaDGgC20y
Q2f74pavgND6cH/U9BBc2fmdYmbibU311nuFtZxrWMB48BSvMvKZp5qWamGr+BJb
jfNTf0EbsIEc3s0NmdBrWbSxf5wHGuvBWkDWIPHEEKQZPGB8g353GqiCXGwse7PU
zJtHoqjR6JwpDncSqChK/vCrbq4SfVERWs+9AL3utmhQ3qkr/8JNPlcpCJIO1T1B
8kbFmlyHk07K1oMFju1Nf07HfnDMISghcZfMdu/mMagRbXaY/+vZAyidTn8f4e/S
UK/Ax6fblehY084rU32Y4uKp443j6+efroxTyI2MqpRU73yeZemko7wn4WD8HBeq
nTZY5f0hMCcAY9nEB5OrImpDdbfaMlbqWHWtRZYf30ZepD3D0QbSAip9TX4RnWKN
hhCHl3uu07BcG2vR0ljykr/iWgsbpS0ZH+sfnITXKNsS2dGYXe160eQ0v4tMuHmx
uCi/3Csgauntxes/g3ycnqXYhZBfs0I8FhxeTcGbcE1VWpnn5D9IFbv3tYPPHeeD
9v+10PQZRvhx1Q2zheiQ/I47w/qG8gf5KM+RBAIZGi88GOZPZqNopALS9PpDHB1F
8W3w4emNaXGQ6yzJ4OmQR/75p59Z/2ACpnA1PhtyQAxCyzc7DV1OrZTuY7dJu5MB
1jDnrM9j3cRCN2TGHIKMVhr4NSle58CWpG3wdEayQAuMYIwd/c+2LnBX6E98ZaZi
TJzInssFDgmO7D0RzVjfqhWg0leaqkWEZj/1gdstPuGvkIvLKkYJ4jGpBpPYMHEW
hoEPw6TZJ7ypEOOn5JDe9Aht29G1tDKbz/Uf66VrvBUZPj/U5hVYbbGVO9bg3v9p
nEPMNW/DAKc/ARoUuJrE33rw9RthtTTW4e2WuYbXj3V+5lxjkOfrl/3xpME46SBH
wUTSfklbAXHxOEg07/DvC4Xb1UAX1aYDsOXm9TkM2H5ZewfStErt67GT3RTbN5TI
yl0OGCWbZboOkSp8MLByNJe8oEasRctUaponYuxgFsZngJ3R2ZrANgXFMy79VrH8
eq3DjIFWpGRIeZqfdQrduaPMSb30X7Vv6ci9iXYOSfJ+JLLpdXsiMkX5miPYDYuF
zbYUYUfljLfkgFS+o2Va5Fb81I6ZUuHyjr4airPQwyEvAQSNgqQ+Ax1ElswpRdMu
ibdPcWcggdbPS1fng1Ye9UnlZUEybsMp+xBoYVXKsSZalbPqpSYn5DVtEw7q3A/s
49P3/kcAp3+P+JZMvJdqT3cmC1Ti7KQ+t+/kbZKdffYhV4sKk4u1Rk0tXqlhrZtF
O/ZO+sFTUPyVJfta0tNMuh+xhHbR39YFFH+EqLEpKaLPpYATfMzUeF05OrYMDDKB
7ISGD0DJlzYpFO0hVxoXjHd2rILXCEN6t50uZK9of1mJVDmhbhUlApD30uGIuCab
n4sB+/oEh3VBSkz5vq2f1ChXeQdtzeCzqO+pxMeI3VXEs53U/+M+pLqYoa18ulJJ
ENQtW16/AUPcvCZbeNMgX/JqHUeIhAtALQv/2UBJWyLEWBFDE7eqCqCl6cASqwTn
3dcUKfFWgVa1ByKjXNoVjMi80pbjhz+fDuS2tWsYyKGSugZlf9XsNt7lhcddPbCg
nkIBYbH2dZ6VBV8NAppZYNZPS6Q6f/PzxpBapmnswjHio9xGO2AGCI2fFd8lLXc/
Za83f2B3hJEBgCp+ItNXbeBOTdH+BguH5l6PnAw0QgQWMromIRSDy2ElxuKpP+1i
kk0TxDAv1kiNLzbzOKOMx4ZKJgF403OekNOSHzmqH2wY+/81sJDIp3w7sRvsle9X
EuEeOOeiGUXDv0BDb+Jo4cQ4nQEnMiY411Ws9tLv4Yz6p4b5BlGCWENDf8bE+6vO
p/w8xToYytfN1ADr5EChz/q/rJhHH3Y8el1oITcFogZ4D4gHDUW0+itilMuCRDoo
pSk6tVuCvDZLlY+w+9m1rO9NEkstuQjXAyTwKxCc+zgfPKKX6DUf2LvqSM2k+QBI
7tKlwteXumAHtgQGH+63gCzWugl+CElsnMDpLsjKQR3looVg1WjNySSzN+fj9CIe
JLDkYuF/B8NwZZpDO/tcA755d8FWglETFkpy7ik+nMmtkg19r9ikahpFUEcHeXTX
S7XNYwgoPAhJwFNAbSS6qm5zrk7KJchW1QCTYTNSkgaynV74HFwfnOJkjwKEDhZp
e29mspmu6QAf43uBd4aR5L08fAQbhMIMXFu42qEA+itc1dZQtpWHiRPmFge6GcRT
KZHu8XCDWnyp9gooOxuOiDo/bCvOUav722r8+eOc8/j4Tj8CRFVHnf3Y/YbIcii9
QcLNMoLtflBOzMaq2Jf2B8X3sXhp5yNXlCJa0ychU2HCKbS8k6rdvrjhPNaltjcq
RYEb5fvu7WOGk7Sw7sjPbpcpD3mwqSGTQ0Fnfzbrtr8hbDOUGE2yBrKUUbqQNJ6z
+thY7JgChP1SznFJ9WzxgEexr56JfIgHL8Bz4XfQ+ePY1XpyebcZn/W/Z0NZoqJ4
TcOIGzrA0weMxz3h3fUobfRSHPRJvAy7npobIuzP5QCkR2RhOfwt/TWXs+rsiILp
iuv1mnAoU6uXstHoLxHuoxxDwkPCGjjHl0i5s53Fk4nqqKDw+gP8SgRhqsk47xaq
iol9or5dfF8eNClnnbeUPF8rxdWKo72TrLkpKSJ1YQ0DCyOepaRZHMlUEwgv+2/8
RLJ8t/pAlJDAcd2I3++v+1RfE2DytmmKTNgvFbU/5o+1bs8CVlv7uwfLQFzQmaaV
PfXAwtmPnTAQQ4Ar+Sd1FxCGdG5BBQjafZ+lwibNQnGY+uGKroDNlZH16MzHCQW1
bLFYRsApvppmYwwGhX90R/zsDt2wgdAx1GANeLEnnNx5+DNLVaGqSiJOfhuSSmNn
QGSj3Kox/6FhwBKlsh3v5L44ZDvLbENF3leBPvBoyzDDuYfZbFWU28UoyOlolvtT
LjNRH1hPq1+OHNsCcm6Nla5ZI0wN63s7YhdfJAwhEeIS2o1JRtP4D6yFnxRXqhs0
DAYxhCR2+yYsDf3b8/dsN3cdoz1SQlUV9SJTRTkjvd/+/HuW6/+MRq5Slq/EjsdN
LI7Lozk964TNtgD8D4yz1tWRx4kdmGWVzdfyOUk9oFWoQUa9d6oMVKNtJUYg0JmD
+BB+EHQgwcF05aCs7EtKIUMqAgobWiYgkEwB6YnFDwCLfG7DoMVKD113EXNlVVTo
SLtx/W6bTsZW8XMwiblLfavDa5cHTeZP+GDLoieEMghSfyt5XCRtZjQI7QeVJfXc
ycmNp23Ek6V+tPA1m4HH1lgeLbNdTeJfT7KXWm0e4neciR4Q6ZfbM7zsX4BnaDlQ
GGfmBtPeDv4xWZs2B4WOm0l3PHetbEZKKJlhkJP1x0z3Al9FuPTSqQWKlDslImEk
K1AfGo7YDD5fjN+fNneBviKi9YDsSP8Xw/C91+7DPqLFvwYrcbSphAHJZjGoDDcW
5uT9tbH1wPDFABMQA8OW+LKBK6Jic4VJyOZJdlQdFDKwM5RTZxs7U3/2LTQt/D8X
ZRC/1YNvw7fCowKdfZOiK+3AJR1178Ffrf7UE1OZ00+oTrI6rvsc+9v7+91s1SAz
4zkHNu6H9lw2/imlvHFIbNYI+/xJtgi5dg5DvGkspjs+ocHOr/BokPsk/p7T8uWC
U+VqxDyD0R72NdcZ05XqUCxVb1nCkH0PQ+tccDCRKrUV+on+kO30VLaVMCezneO1
a3YaphTW392DcL8NGbnHlVnJlYMQ48ahgEhYMb/dD8EtxR9+qd5dspDDU+Gy6Ign
IQBTvR7Ttm+g8mFP0fAZ+rlXO9hsGDoC9OckdKzMJrW1sS+LJVgycR+x+3bwmB4/
7TPSvbldd0NgYOl29YPQ9z2pJ4hn5GRMf+KRSzpszBIZdPy8az3F6dyX1LEkCY1s
fqvZdWOBzKNoHRa8EWqNrPtuXYI1RKy1gLkNaO3y0d4bkDMZVD+t1+KIbIdyqgaM
86e5U692uv2GDRsy9LlLiTLueUP26+kMVzvfA/uSTJxFBeMHEu2wFjcPDV0EcK8B
E8eXXdV5EoLXy+CXRjiKXv9Kp7H0IbZWJvilJkqoG9fmTRQDtjizOuqjf27YnRin
hv9JoypQqXBnEASbjf4c738BOkX8736L7lHqwq1T+LUuvBNYJ8LqMrIz1k8UIy0X
6ZBuNhzlI9lSsAknGTcEpMNDZILGc3z87AVfiDQdCgSQhv6BKoUM+BIMQ7xo+7b/
dl9T31xMqvEbtJVuvjxc3RVedJwiqi/9VYPhb2QTz27NQgepBnAfMCSox2sDuc5Q
kosx4AfnaX1IMF8nyBUW1RqD/JjMnV4V+xAT59i8XhD0XL7GCKh5dZFvRr+3GqoW
1U6B4mBf3DgKrLl4yo7D+e8kEQdO/dr4I6UZfeFh7jIyBc7Yk333eVyADUzj0oUr
Sh/rnZoN5xtZTwAkZLxTS8NsnBCCzBXHhp4ZpWsRxR1OnDuu2fZ9q6aY08VOC9cR
IDa60ag2kQayzejueQSYlNBOY0THzHdNtH7hGC+E+KSiYmkLRxK0TKaA784V1DS7
I90rGuCnW2ktVk3Z1AvUnhgY3ID2dP1PE0AVNau0/SRhgO/SDJ1p7JTNFYttNyHo
WyqYq8s1V+FVgyYG29C/oBbcH3gSbjtc8uLYINsuvL1h2K9UFzCdq3iK9DrKcOes
5gC+dNi207RYiUkT/QX5KxLmrc7UfpcVU6Pwfn5yzjXoW3iPNU5HK8pDIFWZ+JyI
53xoxOMH6xuJSYo/FJgs5FG2Z97qnJeVfUnEt0e8Vibl71EG66DVA64fDqWEIXKe
tY9rILt4aUebuiGj+VwQvWsti3xNQ8A69cBtmTOLFFJuwgsFJTBjHFElKj+lfEuI
uC+4poM/shwNwPSSIHrTjLcZNmzeQFcxV/zTMBKyRCB2SNqi18NDZLZWiJhMturH
77h5W1Fn7UIRx4hxgQv+QunZzDs2KuU8rqXnyi2j3gs+tzlFtwLval0D8iDnH+XX
48CTjDNy8vp+mTn+7my46H6F7UAKKdCP7qfIvqpG4LeA3lSMOSZRIO3w4uEOzHO7
CfwwP54iteyhwJTbZzUrZRXr9KOp5aszFo0aCkK0/YrvJIMA3z/QQu+DL+lGU4lr
Wec0KVipWCQKOE2JNxOA6pnyjKg9alvm/Aw9o84d7dJX9E5+OjtOwlFiWcYdTlX/
4bcUe+5rUY6cdp47fKy0h/4HS0XV6K5+ElNWrMGR7Kc8MVoMGewuMx89DRgBkzfK
yytU8vpRCNotW8MeBoaOFR7tEXHee0c/h6X87SyePNeaXzYxLniy5btDDK1x3LPn
SnTFHUbjfFDRTxjXAdi9kowLXsAnLf7FeCDENzv3awlou1nQgLj1tFmNVQyFl3MM
Ukk9AdGN1deWeF2JhIN0lpEMdDZjKZqkxrYIbArRkeoCpTmdAY462yQ4gd0ZKPfo
Cb7BdhAynHhZDn+wZmG3CA0KrxNfNiU8VyTT8lAEjPzjV5gYvpx6obYhiUiDqLeK
J0hCM/Ot7u8KY/GcnD8LG5eJRqtIIcseZ8FBWRsemXlWkENjmPRfT/yrmBBicBk4
1gchgOvgrMYyfO2VmP2FlFwxh6SCliXTjR5Lr874ZK76tIw7nJ+wbEamSMf/GtPQ
EXFKvYeyoiM8tX3M79GcBLHBXTGJVIbrTgj4w70dyZxR0FwqN4/S+d3QRllFedOs
rK6aNb37NCn6iXmBhlkrGMLphM9SNFubiJO/ymscjcBbUQ8ZbHOwSLhellnUFWIo
0y3zWTZos+wauEaQVhPKct+cMtnw+wdeiEAQtcNVoRmBZC+zisosYVZ2kabG/qz0
4GOrab1ZZA6Iq4Uj10RLdEFe2+UR3mISAuS+JCtvRYV2rH7gthiHm7VrKSoLUB0q
qpQumF35tTq7E2D5YyPTFSBbk1EHDgzJyCrWr5xl1bmkMLCX09d4Q7ELNE8MnsD3
xgdNT3bEaPyj/GVskQs7ybTJ/evU8AuHO8CNZgqHQFoGQLZqjY+ihWCmW55kFi2a
SRSgtrUpOgvwN0QOQBJk2Bme/YCQ3Hj+0MbNq06ODuhHHSVpFZDDyR/EJ1zmtwEp
bpNa5R6WJXuDU9cTOTwxa/uZ/7aQpfx81RKY0QZ+Z1BoPb0xjWqAo5CP/VnHimEX
M4Spje+VSpVv7y9h1LMxLowFuawrqYOP5+YDR32dEy3OwdrNUviw4euQgNySPOiC
5NhPkBwYpYcUGoZSG1tdtpjrT4VV6hRqajvwHWVaYEY/RIrZlzGbrrTZ4YxwK3UT
LSPjhkwI8Yv/xvsKa9zZipCQRuuKg3HgYZhO3cWTa3CYilVWbm1jICB6YUDiBuED
l3iGze98ibXib4yVBmvfAQV1/zpCXnaE8wczx/AncUoCXetellfhxAOWa3RzV35k
ApxeKUfsbuT1jXhVC/DjsG1KilFlhkci0cs9fP5Jd9BUawsnqYlDktACKagT3+oW
ytaDRwQbv0YzH208QALt/lca+JRvXZ8yX8kdhp2XRVxNREUFQz9PPGa6EEaeQWaG
7NLXu6QfSJkTCS783lIA389WyatIH1kGmpbNYVrucmwyKAxElOC1UgOyC4uFx+9g
fxq3MdS9GxEBKDpZG6bzWrEe6XfdR/s1wqY6MQODBUWE3AI9uZWqi1hpFbyzZtcY
x4JUtGAXQHd8npFs4Wi2rDJtD3hTDqw0Yd0EmrC0Zwef7Jf5V+pJ7OsBnJaTkb+6
XadTprp9m03rxUThdLcpUfYagTcR+95OApdp+ZEUm5UfHIyBNcaYY5ixBuRBr6PW
Uke3jibBhc+DDggoHqp5/8sOhzzRg0lwfZenpTBLeNPvKyWDlYoU8b9WP07fpPf6
1/zVkP4zqhr0XRtlo9nfv2mnAwT/hBhlvX0DqALeTv92walA5uxH1pCBLcpaAkYM
eFwoSXi74G7DUdjtYAoQ8kLsJzXu+zYWEGyOg6ub1JLybtQ4YofeLc5+qL1KCWWz
npbx0Gt0iXhrQ0lfysJLMomsRKLpxMNbjT9qWoY/IpuPCE3dODKMkPkQxc6A+Iht
L1QiLqt9OwX+2Xn3zPV+SW4f0a38yzs+S0MNT2aWev6L2TQUF6YGuoEzt2OGvpgp
Uar6kRSS6KHkL6mSW8F+hjyROH2A9EhbiEyqgh7n4OgCunKXBCIJOXTsAQT90udi
h3JgBMlPwm87yJrRDTfSummdAIpF9Er4/w64Ob+wCpw6gdL6Q5Otc1Eljb0m5EoQ
oyhBxfj/j3zaN1yHvmQxfbExZVhzYWR0n3YFvBPSbOHrzw5x34poDovypA4xXVkL
iWTtcXiUuxACQCFppRp6sJPJZC3R2GhvrdSm/BTdjcHGRA+TDuCkC6rcD1fKoF0h
/hF+jVkwgScBi7TgfH2X1i+zH3TwNrvF1bp98SeqdcxcApmCo016yrEt/nZya4pf
0q3vraifo+z5UTR7t8pYNciQkgf7yg9iz6+Ovo36LDUxHQW/SfsnDxYbhczPmNG0
1r9EthO0mR34U5MSqrTab5sPQgbA3W3NDBikIffNMjXHm65YMmAFvoFpzPpNUDQ8
pX8TZFJGZsfY5OP9CX4d8m5lwKRclVy5JLFWtGcF0uoQ56kiVR2xL3++hKjPj5QZ
IXAaEliZGmbakCbs79gkjX4YcE2i5YZDpPdoiuq//lynr/1zH85FDTGGcSMTb++4
O2prqglmDs5QrsNraxAVuP7bcj09agevxGqznlrW0j3SI2vaklAUffV9r+Hy1Ess
HrLyNR0IvbQ/TsCvXe3ETInbk6T9QlNOURe52JaNhNHk82OZv0ESFlFW3RJ7lmbU
PcVHO2DwckDCMBDrMn4GYUKyflVoZN4dM4mtdPdlvrOfRXY0nB61o0lMtIHooxo4
YE49/Yu+q0/hHfKzrVfPvCUZRvHlSASRcII2QqKjvyNy/MMHixt4GJS3rNE5TS36
hSdC8wdiqlwn571Z+0hzCKMsgnYdwWGb7yFxiu2uVrFEU6RDSVIERgkU5JXnYT7Y
4YrGxFvQrtjrf85Kh6yGLrZJkJS2MMRFy8sSVZdM32ALvHb8jNIhEzTFWvb0YF2L
pwqxuN0eexJXb9DADqXVtZSuCscM06lVqxlxXsJK8xVJ4/cCvZPmok4n8KAsSJzA
rJI2CK1kr9w6KFCFKZZpf5DGmYVYA6gS4X8okdnF5z8uDU9scHrKOJWvaXrIdAR3
cNmre5XOIZvg7vCUpMvQxANq2aEM9ZJSteKW8tcRngWnw6kI66IdN+rFEgoUKoQ4
SWV+4TeYGzQuUTW86j4YNhLZEtHk8HDMtCMlZiCOnDDPlyB19pJqf2ErXZw3s/EJ
H1DUBa4wDxho+AAQKqqUBUgD3U6H8OuV+hnD/TlHEmQCQWpuD7hdq19qLA+W/WjN
+zllhsLV+IzSOU4Q6tiUxXkwHDSq0ED6ZOQ6Hvd7fEeGrBoikrzL3bWGsJN+Zt7o
OaQV0TxENlkLZKmjlSkESgZQ1DhgUWHY3lER0wsD7+9QWc4fxfBEo/5srs0pTT2O
jVP+ASalyo/WbosuoX8Pp7r/rwYNcfSVHLF116jqsQ/nU6JXLgijVYn/hrwj2YG3
GgK8LZt1LTJOc4yB3hNVAazeX8u7oDvk7J9MkNRpKOhHl2nYk376o81WZO5ZKApM
EvM93z1UEq4LrgiaMTv8iywh4DgTIr3C2e9rgOzA5HS386VH8EdgKKDSBT7UBaPh
0DhcuF3ftKPKBgCqOZtdIRcd7/y5QHMicN2WZ63xCvYdUWlDT9ses4FT3RisdI8O
ubG4S2vxs5v5N8hyM4jXNgP41Cjjau754WzIAr8925ywHykmYvvUvRqRK9nHArr1
2eoS7fS+nlCBV5VVNqdnVker0NUdsCt4OMLsCFqM/Pwyfu4RCQYJw+cg+0kfoQ6t
Ssa9iVhpSYzV2om/5grEZzpQE4cntEFByebidOWPSW99nV6nIeetopFXhZYfrgPw
NKJK7SLLXBDIp3GzvKDlXCwO/PGCPCF48MmANLEKMlI1V/AU+QKYodHU+Gr8OJH8
SukPkLsBS2U43sv1gzIB8IIqPXwIPKgZut0w/pz6TkeRhCwMUR1yfYbyZIOggF31
/i7I2GuYr5Hnql+u1vRTa0bA6qRJnYvOt4/p5CPgWv3nd1RhQt1+ffzAwZds9Eym
6USQnplOgLzLGAyFf7ynnsWVNtPXQP5BEWyxkVHqo2kM4oDXqw6YXav9XTG4GSfb
smM63/3aEkBjYON/q7mfxSHj/gBBfJnrrL/7l/Gee34qWGe7uIMrdp3XKCtGPgTE
GPK11dSGSv1yA9ajKMp2KczkuSD/PWhX2OnSx1TKMOYNb/iFZ/wqMDJ0dlcPpnZv
KnB+JSXrpCUzBB/SOSXpzrnahJcWQ5CKwV8vt3Tgm9HkLW+tBm/9nxcBFB3UARVy
NmHQ0F0yGESfZ8DPUUtWEj4TUGWTLoqBt1rm55RJXjVlSkR78RBvP+gfStriq4RR
ovNo0YM+n8LF+5aEhIPBAR6xWQ7Qe2DqFO1/0nhby0HkPxpE5rDtXx41NLJZOXH7
+TO1vQgXRJ1QVPEaiCTQ2u9D3pG2bDQ5qBP4O+JZXScydTCZfhtJgWk5QKmRcWQ1
wUcZxE2aFZf+YSIDFyVvTnrI1I1o6xKtyDgYtQBtSBNoU37jUTZ3yDIfKvIQcWgV
TCiNnxE4cxlfZIWx4I7sM9nWKsLZTe42P4p9OGZUyRoYznKVsLrbxHfohj1xssMD
0Rdwb7wJM2HETeKZ71dHEqoGa055qvOD47alHe5pAIIn6lxFapuZqb7EGMXB1Qyw
kc2vq0mHbZgM2J8AG5S/LwqKX6Va+HAfZeTVMTS05ZVI7bLmFWJ0lKnsLTDgfVBv
8ED7vdSwHYMkddndBICygEZjTlkF+J4l9vhMvVU34QayjYHg7zfqRSiB509LDTTp
DvzExZixqLqo22ZKSh2Cg0VatR5axQa8hnQPBmK7uxj7xpcjXsG+OIjJl0v9Wh0j
EYPrTG78I+pmAMEBlKAL2ZY4g+HSfx1KjZwpxzjKFZYpgbangheBFTisYNPoJuTb
6AJKG8XTIS4YDk95OoFj35wTNmkTafttq29uECNWneIbxM2+NSs+AwbN0cKfGw33
Ajy2bKxWr/c6bWvwkF0f2swzFO/aaEChrDyaV3wqJ9EykUl9e9kNtZpPuHFIpC8C
E76hT8rlvuIszRGopbjmEHvu/Werivbs7BkRm/OAPDFmjNsRFSSDXJzRmhmCEOvV
MnYkcA0oDkxDAe0hjQwM4PaC55mXwyLb7wLMewSN/hE5QXweQ59FQnY6Eyl6KrYv
EIUES4gjGUnMyTyK22gofZuJMRrdvy2GcLTIJ8lzRdIokUkOHFsfULg2bNmVatdL
rJrBz0xdz0jSlXcMkaosMuCItZtnwI0v5uAxPlMiOuco7aOJKTkdGu++boEurycp
mGNbm7J2EcnjC1c1Hv5oi/o0znpXlyNYXlsksWvtHeI+Lwuvv66/TJvQrfISTx1e
EFxhlAOGRm1rbnVx8PZ/cOXE+F2U2HkQdaJVD3ot7KAgxWhlpFRaBDzAhA2Nhzti
PlIlelk22+H9ZYQsq4AZOlGQeHV3vHmXQPRmbPiHO6h7gWUjXz0VhaEYzxBZR5xs
LybXs5dBp+y4eBi4cqv2lUs1e+Iq2UXR17DXCpPOy4pRkLgAlgGMkXJFTwU2/YWC
LI87noiUSONpUH+mEKXwn8SuegE92fM9OKFtsQcXy4YK3fqCd6BB5fMlBs8KTEo5
QXjCKa9YsGPx3PtNbYJz1k0DaDNP5KQoJG7tH0ATAx6s05fS2k/PEYTJb3DJ6ipg
8t/ow+LsSkhdWC/SIAjvIOnb92lk0++vpjD02aAti8EGR2Sh6e5tdYjGpBjpqhfP
gJ2poIFkNCTPu7hnyIEF6bj5Eg1XbANMDnIXFKy+bvIGagotGFNlpIYZWyDG1rke
Lswav+GmGuLiWj5dbukYpeh+PJgEfINmfvTlkTKgwKHLQxNrJJmfAyNDUr4x/5FW
b/ah8nabklhYfBuaUn05sYYEpqRwC/2hTNzki2uER4Pbp47h9aV1fIN4EbZxDdzI
Au2Em8VwU0wJYcIrHs27FsqpnEO5bRowI6W78dREx+mGrUeVCMWbwYPeqjzeaVTY
BXANpZwF4gaj+xR53Qe5gR9CCYjhVWmGu/YfG/js8AJXMcCat2XzXBESUruDm0wt
h6fyA5pGxlyTxYIfT5ek4xiVuUoPbyHxy24NdsqcJl/w6Bhaja9V2OyH1HkxdTBA
KC2hjkS5ByDFYvslxGSXcBLvHTUh/ykYgq+lc+btUExnZsj0A/zZP8GEhyoT9rWj
OUGULfo9LA+/UkPonGkAQMf1wNEEtiwpiLL5fd1hRG/lIXqPhRqTxn6fBZ6QXc/q
9QQvWgHK4m5Bmz0AjP/szxCP9RbyH/lIFyrBsMaqzGDKie1Yjrd3vZUnCfShxQMh
GMJmbN1YnhAjm5zHyoQKt/PVtEvaczAthCzmSSLZ0Zgp0KHnzOd7glB+6Z5MMmeY
Smu2h8J8iMUa9X0zxXq7IgzQtpFUZjZzfAbYakGYg9SRBX2c57An8P0pu3JPS1nf
dVOp/DAF+ooxuf9a+YrbyyVWnOWgSvdCW1dXvO6uLjFhzxtTZjLaUZe/4gu22Ao9
ZSzAx86Oq3tUfTTvMIOvj5eW3jQYjJGc+6fL0daOIriWdGRMe74UATOT2eBDom7J
6MfDcJmYoXmyhYHpCLxCDfiKBFre43BzYUEaE3C3U1YaQoQhPiq8YpdU+UXMIFf8
sguGV+wdGSHRYVKTpqGnALfn4xRFBFmGC9dFApbOc1z3T3MCdnatcByYpTWAC/e9
c4hz88Zi6QFGoWS7m0DyIhSVnIPUVYheDZmkaOpScCPCTEzPNa5d0P82hltOQIOp
lBqCMpb48t60QbbH6L2ZONYIgWNj2SOLKvqfDUpZw2jpuxjQVQstB8rfmwGAQOzP
JurPVmiZC4tRaSOtFi6d/CtAIzVK19OZ+QhLxJsCkEJ9/mV0FgvQnyANT9LfHOJa
oh6phbVTeHwK33lBz4vvUXmF0Md5HqJ+CD+AX1ziX7ubcyrLJRLTm5nnFp3TxEPL
+AfDtDC9EasRetHku2J2Yi4vTVsU3i/HQQJmTibCxvhvxpN3yqHj18GXRWOTcbxr
1WtboqRPDPYV5tF/LkazNzZg6MTBvXh5zLf4seXCnsyyyt9wUm4aNm/gGhntePEq
I4O7QyGyDp54BM/d51ghPYWEkv7Ywlz541pV8i++5ars3PV6K+xRySK86IdZX+U0
lutfn9fD/iq2RKl3AE5F8D5aqgxC+iVMrLpTLHezEnlUe5EqeZUXvS+l049cefew
7xjQCKyBp9zlhazv8Q0JED4KKnpx8FhIeg0toOU2byHT5oOQ6Xk3/2opMoOUn9xs
SjitoAFFY3wsjQ6D0hLvrTuAOBjDqPzx1hmVrdmz9MNANfrFGjFjy7WGN+KQCsEo
/dOstgGoH5IHbYSqkTL5dAbwWU6WtNzk014eMqnvHOh4S59kfHzmSkzVdttBFOse
im1R8IfjeM6jdDqh79iOlbbmdbBuPFWSfDE84mJt+WgAw0nxofQJxmOoLUDQVxqJ
XPP9wMdt3aQCopIpXYF4zQuEEGF74nGUVeegs/adB2H5TyTSaBbN8eOWKtoi35q0
lBjXuUu0lYvStZoCU0OOyW5BrO1JJkuZKaQ8XURFtpSB45K77Vd9uurQ3IelVOVs
HUELSp+/ctjpSnuo9oCwxNcpyRheMy1ZYuDcgFVKMIduIysdYdUa+di7+76A6dad
v/vGFbYY8QmGNmRO92NXFLwNH7unpZfTJKWh11aXNsqM3QBzZgKqqXwI1YSQGyjk
ZJgilu1zN78SmBmTgaXJbjBIOj3GlNNR9Ugb9jpQsOkATeCkHNM0XA09ueENijsN
GtwxZCj7/SlITaNJaQEdCrKWDwGLm1jCI8S0YwdPvLFKUo9IG9bgZxHGmI+j0+Rr
WFlqGg3eQ90+FBQIY16r6BL7pXHIaEVWJLL5dMzW+ib01D6MsdJlm666lfupzQCD
K/q1gqkA8G7CwjGoVLZz/rQbYZmbHDj4KMaMwinMAVdVL+8Sn+TtUtIDHk1LZHH3
oUblocC6TxB0I3ygMmXJX5RmHRFa4YO5l7yG5vlPTGMktK0tkR5AUwiZ157NgaXL
+JOMNzLLGgpfNyc9MQPm7iyY+alCBsvIjbqH3JP8D2syU8Zu5IiUaANO+nAvEvIK
j1OqNMonZaQMA9ugwz36SdcDZCKNOahs16TWm5ED9qBW+G7iYibTbX0DzFl//bTO
bXW+IbKaqrhGFJuu2gjbJ3VaO2HmbU3BYIYgDVMVa83h987VO4VJZOJVVMqFreAQ
xLh+UoSdbafi06QPLNpNjcwqtYhgdIR460aEP+YH7HnZb2+hCT1lWdtuObBdYDaP
vaDQmXQUsM6N80vGkg3ApaiQRtIUstZUz3vjquzDGiMM6y8+G8HZQqL2mmPr4aoo
NtS1RMm52CBss6a94OM5RwYCl3M6XShLDecVJfweIVs2EImP0UxRD60SNpnxii/L
KuO6ThJ/aJj/FTantUi6Y1+rUUZzBCzwbadn43QG25pHaAw3daR5xmOZykS6FnaT
OjJ4BUEslu/IfYQypwT7MaMtevOCYKFL7HhfmllnDQNCxldxNpZTfSXs7Ud4s5vx
z2x8wNbpEuaHFyezticUCQziTsbXD072SpLAU6m9NOhKpdVTex18Pk8jYl1sDy/v
Ft19al3tIuryeCqf6w9mlnq0BWf4RtvhjbYhXRit8sOoH+ew5irsaEpx9Puh2zN1
xZKr+p7WF5cyVbxqf7aev5xxwcWUvipgjIi6Y7d5V7s8YA/ir/BkOqy54AsrCoST
TkEr7AeMYFjgwNW6enCEXk0ihl+to7q+y3n78OGmyMbtOGBD5SHQkFI6v9fOYYC4
sEvSTpfMSK/9en+TZfQ63hnimE8vjHlukk+fuCxN3UKRv1+cVkmuf3OEYcYooyCL
FU93XKypEjwquAacg6Nqj7uw9SwAfN6yunkKj92KUaAlIErJXDhCyhcJfgRQJvmC
6RPSFt0EIWo0K20Je/nQTGiVRP1Q8MkCzLZVsK8wb0ix6Re1eZcJJGciubhIS7AL
XTRfPD/8XfJvktfYquN/uOgNV7T/uqcNjfXeq4k07mZ0gGd5vCF0o2tjSS+M0AeZ
knMsGlNiPre3aYeNmZzptRuon5VXXyQlDH3NvxyDEGLAQHoFAwJd5gdGloGmwnCW
idHwEjgpPp22wClodelNnvyjMBsq2gngv/59W/560bPxchIO2f7ftGmLjgjt7Gqe
GzmdjiTadZ1FM/QN8cZ4+DiPgJuqwMfHbfYg+5PHGI8UeqORKwVjvQU18EEHONfi
wJNtb6ChFXd/ZrlQylvcgKjnyCiAgi+PiXfY9PQsshf1hGPLyRwKI42KWU/Fv69n
EKKaR3ZB1PmFiIgMy8Q3rmx/qj4s4jUUKCXREL5db3/sW1EYSJ2omFtxE46FdL0g
oOtdYLYjcP8tzDcmLpCHHvgejJ+Hd8L7QONtO9eRY5Bn3OC3RY/CZqb+bBDF1YSh
JGnOviUT8y9rT7KEJCj7z39Kcw4LyjkPqMzovxm3vqDCUF79IZqpy2iqcDMIdylp
KDzuOhBAo+pdxgnHmoYb9V8RUKGOg0W4Qj8shu577VTvscc12RckmCVBWWY6d46F
x4/216m3+sd3igV5TqMC072K/EScu2E/IjQLWX3zu7VcqIWQaGZbnIYerpzsXL+/
GnMH6tb1N8BX0nj3gvgq+w6kjdmJ38yahMxJngOpPq7fXrdWRLiUlSn25Q+c6Ft2
ptxqtc0sXiMn4HznpROz8w4zMK1OeO3/Yj+mU9+ccTmmxiutM+LHZFavrdCqPGON
dxMSp1FHWwV1XUBZWuXBDaKPvP8qvrzVwyd1SMbHdQY9odC59fetGUiKaGyoHIS8
trXEZWJ50fM4aH+Y4fOm06/Y20XXFwGdo2QF+W4X0OQQx+APfXanLHsNBIsz552I
G9xTqOZP4HuP/fQyvAmqNLZBNlMYLPVUwscB0w+UugKZGz7axiku4NLVHJdR6l35
9IK5DrAvF9RnUGy6t2VkOE2uyZLSMgPwW8zQGQ+/fviFN1+BEFV1roC9JBH4gOWJ
Inf8xtHuLndpBcP7jqnVV9kSVkY01soaGW12MMWsRgm6HEkBWrH8s9HnIa3QEWKm
MHb0ed/FRo5RTgfddXoNv7ImNniiaz2+peRUVZptPUKLyFvN0tLAJ3EG/YQwbaSh
XysjbuFBxvH7V2EnQjNEbyX+bs56mySZLM8HkqNn4ZB9jbD/50ruaV9qjJMkOECb
vGCZsX3zzq2YcSnvBqVhgV7wxvomh9YvKwbJ9pRudpE4NY/8nbgUF7lUE5x0jmAB
efg2TzS4gBMDc1ou3MGSQIxwCmt/1HPs0afn1qwnWcBzP0lR6bHlCTXkklbhSZza
d5mvGKe/1+v36I0s0YRf7UzWu2mNyHEwX0Rs4k7nPfvQQ7ucIufr5OblSJGIGzWJ
/jeZQiF1Ryt+R6rWpYeCKqV35AEsu74yRkqyofOuWWEqKuUkJeLh28ty6hLi/WPV
VQqfFNC77T4Fq5fhowA6WgyUYWAqV/XtEe7+6nhbQNRXLXXNC7L9LT6x5yR09rp2
lJR3ujpVPxK1u7vNCMSUzTc9XwUIMgKUJe4o6dr5tt2SFJQv/x2UnK27f2XeQk3y
oSGSoracKqclgCz/DAMfMMjFVnx08zjdTAT9mhgoDSWtCmjvUDHStbllt6hZsoR4
F5p7vsYUUQzN9qlCIEzXBkXfehxZ4Gg2Hlv3hJ7tG7azNwByzBRFy1DBQUAcbpp+
dVJc56GS5IOXnnQosDqTK7Qd/GLQie0jZ5JdPQt22ZOzcIQPS+cJNEchljGY6Lg2
YUi5ZH/yDCJhMpT6lM0y72mh9XhD1UHLO9yZrzQMikvF0VH3vM/BcM3Bp8LJDQvM
Qwz69KUWSZjc55UzzQoqI++2m0ZWzJBK9ZJCQMLEll1cYPkrMs2otPeTjtiT/vQX
fRIghcLf9CHeKGxKfWbc+pv8WpupkrDVQoXYKlT1V8zv1d2C1ZMj/VHOmxa93BnL
eWxdXAVxTEQWd0r4y3xCbxozV6CAWOSZ+IJCf4u6xR4gXOgL15JqvYpPHdhFJ8Qn
N4qvUzHYMcB5vgorLSYHuVAxJPs9SWQMuT4zSRMtVUdDY1yABeRxOtZxLRWB/LRL
xKwOb19IQbOBac7jS77euMvVSkrVF5Cl+2XwmCnjEimS6OH8pbmzFLKAmsruB44t
r1VIdO5TPxiUbnKPEPQ6yB8nSeSzkNoL9JfwBnKXj2djgi2WYEWC4WIHXIdGt1TU
npZFBh2Prrh8UWFlvnuos0S7vBoMx5Q/KvhT1HarGq1xcDm5Yten5E1kYKS0wauS
b0/+hI7YxZEj/yNN/DYhUOnWHEruh9HOwVNZwY+pCKkPMbtnLNTkN6AO97aQjWsl
acGw/HDUafYsIWPaOPeh3ytQAhcX2cW0NmPhR2zPXjnsdZCpULZIdrBkaT809jPv
T7WOFa+Hqi93M8lmutKHpuRHEay6zRtbqR4c54qTWiTf/1IiuOwHSMq5AoRx4DKh
O/Qa0UvparsdXdPRklYXVaxswxrEjcTFp7AG1OikYUiDD24gYgbo8V9jl6BLxZyF
pEuetmtnKqih1lAFZD4MXkWf8O6Ud+zjOsf26yvDxcubItWonYbdcheczjP4zFV6
uQpfuZ7f6PIAe84t5WC1HH9trBJUoArNC31fuLs4kFdB/38g5hws6GnNj1Qdd9Dg
gGaKHyUPuBQYN3QQ4L3+V07M6+F8mjcHrgFFwOVy0baA+VrP+4YiTRB4xOYAEmND
80wOPZZual21vinvx9FDDbyVBuhJ3WmnjVVPvgXWFm/V/kprEZ3Ea4rabKYIhH/I
dyYmSYPYJ5X/JxhcDmYpxaVl9ewz4359sVeZKdaS3XIh4zsZuTmdMT8sLIcXu1dN
Y1MahvplGOTir3hXq7iKqsc/1PgwPl4FodFLyrNwrk1kSOSYlM618n/Jykz2rKJD
aJVQjMonJBmXzS9JqPeDTVCCoE05uaiQ3c3XNNOq8aBdipNbX4E2TbzHTlf/o5kc
s024CrVOX9ZrnVqjgP0MQ+H6HpAZ2hv4UCB9uEWIKFk48tkUIvIQp8B28uS26csu
1bX3SNB7cTi4QBf3496CZLealgwLEl2+/gtn3G2y+mKF3l6fdBFCRifYiP9NeGxu
7r/A0IYZzEnEpGR0WXrbfr/+fTVjOAyRzJ+6vaGsaiW2ntkX+LfJg5AHaei2SOVX
Hwqmgso7B/r/WlJvCTw8m82zUusX+z66pFwHQVBL0kAUqfpbX1mZb0oqQMYyXsOa
y9mVI7RcaRrsyUHcdXTNI3n6tI+uqbM6yZlI1JAtwAj17eEFyHVbraDSHXIRLJg5
NShfhxQYMXNg+6SqK2ATGh+8WODLIAcwN/5iDKdd29DjFXvpsxDZ02cRUcSKVFVE
szx1Z4mcL7R5B5yebpZ6Qq8kOsZ8R9PITAo5oIDcf3fiFxO4T5hE6hsVZTaQpQ0X
PPn6+8xmgV3+xxqA/XR//J3Dp7cHxvdWlKMNDNuxqOll7ydQzt3Ab+6eOKtw3LbF
CfpzWpsyqqEBJ1om5/pOUc+MUbB/tARtx7vMXDT+Zd0rqxlWtOyw7IzxnkcmXe0Q
SW+Ujhb2odojN3M/ySwpufFuMOaPvBSrvIlhveqCxd5e0C1PeFghDJNOt+8X+3q1
iCOLxXn+7W0X+Fo81J09Gyq3EibpNUjN626LGZ7VPO0+r+6nveL8p04GZvUCBeSS
untM0lA/BdTFHnMXT2GZdgUclgVKQX+PmbnE0UmO0kX08uhx3cXOKS99RTSmxs1I
hzGwO8y65cyVZF4KY9kjaDQoUqiIhirXraUQH36bdSF0q/t9QZNdBjZivobOjEZy
fyfTRcLL/Mo5iqz65hCGnHe7oRYuZWwlLPKy9ErCtf8s34Z7GLmISyWH5fruEh2u
FhJSLV5n5zQ+dPumTaErQGBYV+WD8JgNIJUlqEPz11UYVenKWfyWZAGkdxJ4ZfCw
tfL+qqyvUTAYQ2sdxuQz23C6rJXpyZ96cuMhF7jY50K9+kiyC7125M0U1preaUb3
MS1pDqbhirHAC5+xzfGEatCagrtuZ4CvUONHg9CqO50H4MerL/plQrRjKERuZ0xO
eE00UDfjCddFRXV6to6Lts1+yFlmpBl2FwsO7x60ODRezkfuqBkR6kWyAAR9IxUd
RcQinuCHWS8NMMJPvW4VEIPEy7wGO6wpQ0lEcjVGR88fKSf99r7h/r142/slo1NJ
ue0M9v++gNih/rm0v9GR8dxihtOd9YBhqHPxtc5vk+0enouI37lSSA04FmOnf+sf
IlZJbSEYYmjEBGrOD+UEJq8+kYtp3E/8UCBVltSvIXIjFltNqz8WPhsTDl1VPRzT
qLxSt0Ss8j8zfwYfzUQocvnr4WCDfvbkqFy5rRveDdenkHyfE32kedsuNTqlqxSw
f+qOcUeLEajqZUCnI/xmnzJ0DVuKKZQk6GZQyeJ4Gx5RVU/eN04AF1FEykHjGPdc
3MrDUNijknMwICljy/a9whSTm8QBOB1J7/bJ/tpLqGq3Ta4WcONExiy1PAnGZtKA
i09jDqOXO+zU7IQKvP52jTWV6Hdx1lNg/sTe1oFxg4CyNOiCb6oL2OgrhVZBgYFs
RheE9ydL77EAXTrKd3COhpk8m/jnCNidjHfsiz7NK655y+w1cNa2/E1ubqvhXAss
sk+aNmdFXhROiH5aGHpccwoM/qlmVDNHcjOMrKgYLzGcB95mDj7JMFXPLLyc3y0S
+9yS0gN0bmDohJWMYFtESvpnhCaTKCojcGN6PDEPGtiJ71wDeqAsGDP2WB1rK4nh
/BkZt3n+DQHNXBfd7DmrJSQDR/DUX02TfDCxR/zLFqYedkXSl3eE3CTtFOwQaOK+
mr4+pQeeSjqJcaaMnGF8/1RsLeJMIOc+JQU6d7K8wZrCXcovz3wKhnIE1gd2cuMY
tFSGlnDCHLGFamhev1KIr1tgVIcsV4ZQhp5ZimkWAZnDdR4S6WCXgbp7oici3Aot
DolimolP/ZdYztcQrkjj/csgDPAHXhR4kerChYU6L48XqDzxMI4w4jkg29itoL30
y7VrgfGQDpXjk86i/BmqIkKAbRA/Cof6lDRVeKKxOM5exjWPcIrAAbrPJIWyQrUy
toG9IEVhVVZfiekgQ04feFfoiM4/+ls3CrtbF3Z+GpMBUTtFbu80UPnmod611yCe
lK0CDgrx8AoJHs/8f7iLQLqJQEwVNvRWCjpikZ0OoOgRh5DrXdiWlXMC3ckZzpAC
egyMvyZed2iW7SblV3NmYH9QllWpB4sE75fT8ZcjJYGrk+5HNqykeGP2Wh6MdMGN
suO7sw2/BRVDfHW00e322QR6ssTHJSbYALWIMnZi48UGLu3r9/9BEfOT8fOgwvtJ
JfAdy32GxMfvLUfbqpMOKXQkDmdnvnns4RPUbNvjdjIhQU0usz8RTQHjUZjIaQ/y
P1v0Qn1wCNmley8+ouMSZXlonLwkUSq5dYyK72DRSxEBUNe21V7OuCH+/iL377Tj
gC9W7AjBUx2zc9RVtRHb2+VgxcHzh6B/5WRT6v6GGcXog6ndLPTO2dTrU1N+Ryjt
Hwmo3dzaTg2PeH2DjVzxncdOtAtm9e8HThM1JIQZy27fhe6JiC6VQoxKN/cVs19m
1Pk6mcgf+bosB8QgrlKXU4Xzy/g5pA/CbOxMpOqr38WRJikGe5gKakJ27ovDWAgN
E+dQ/DlGtGLcNbYsgUc/Jpg0VSy3r/1ZeNDv9rZc1mAq25x0h4DJ4BfLiY01Rrsu
1cD0JfcqLiq2TDqf0ecpyXqrf+E5AwuO2TWAPbS9vedk4pMaNAl107Kln9zmds3J
+8xSjBwBfhPNbMcTGJ+pqvTOHx4N2Dp+8xol23JOUz4tDMAndhMIt69mIpqZMLRJ
XX9ghU6zGoeh6STjMTcDsZ/jh4YbVkzsJ6DsJvM8dAZICpuc8l2mSMp11lmS2Paz
8P0Qf/L4QrTo8iaSampg3FgknavkTqzDaTn2G1wbMgqJKmRgualCajaZRyMOJEpB
plzYmCaqBLqNwtlizMhxRqQ2x67Td0Z9hdI6JXLHQJH65QH0tQn3AdrEAzLUJBkR
kvMuzuUdFP9y9FmONrT6WloDbt2yG9tHGfH7ymOFzAfKnIjWnolpKQTJsAANIGqV
ht2cBi3OV1dDZ9DpYnIc0L7xo5qNiKRPEJGxVtNgkFZ1PGc6fsL7JCenL625kDQa
lerD/ByNm93q+3j7g3MfpqFoum0L8W2VsYjFJw/5VkuVLj6cuyKTqQ4y5I4gA/Z9
Yzl/6De8ixBTh5k4mzJsWXFkQon+JB7ZJSmp9sryNkIokQqYv46mr2+KwG9V/zJd
rSCbZ1aCx1RTphf1GpGQALXiXpuhHdKQJ23e02FHsH3TnIT0p+yaYVvmd5E5v2o1
Rrowr4xh9Nqsma9kZtAEdwKa5I24bIfBSv4CtDjkf/d5ckyTDlMJs9qD3wzMJu+c
tYaTG8pSGyN15VJsOo02tA/Zdkxrrog2iQsmxlmBVh6R3m9N0pbtVLfbvUe0LCV6
4CKutsbgHsRuU/IECYqQbCLUkmjEMUmeFJawmTkzGG5Vel0AYX5JQH3u4DUuTaNF
ByUT1YN28hO2ziMxpGEIk15AYp3CDnQ9enieUE1StZP8YYflW96Xu9x341TTY3rI
ioUIADq8YU9CfkIcYwLYpEwp6iuh8P3HeXrmH+HX6jFCGdO5KCrkV2UptynPvEb1
cjKHxIC7NFksVCcE4k/P9JhahkNC7GeMjIF+c9vIQBQ57x5RG7Sd6yN7Ygvko2H3
/fQcwWhgSWgzgVJYiATe11VKLAFoEfvmIIrInhqjaQA1jH3Xln/bRfPrJk65dfio
N4nQeXm9OgD+gBC3VG4QtFpzJ/riS5ImF8sh8w9QEV4sI1JALZcRD4NqDqB04Oic
2ZG5rC6gC9EKU6IR6CnizfWeaq/0tXry5PcgHAuQUHZvkGZPUxOcNJCE+2IxSNBi
Tp+Jt47yN9zMrs/vYCvXjObHP1JyV37i8IayLM2YoQPU6ifBWruotAj0tQ/GYU/G
wY8hpn5GBHvQAAEZTjjhOWGoDFH77XDP+Gv3kHJP+evkr3ZyzBJbvO1gM/3g73OS
2iKA7kVe1xvzfXgqCp5NLXQKj1R5xjoow4/jgSb66VCKc/rc05G8h/knp4LcchUu
5BDPqMRRhj5qOFpJzybW/mUAqPwKYuxGkP2B2f01HoUgP5axhnWas4KlOdlaM8SG
WWcTnQoX/3SvWenMKVLxrGbIpNMoHCuwer+nl0C3bgj69FEwd90mkiPS/AEPGQuY
q29k8vcPZ8YbfgDgw2iAEb5e7GLubCzRFlEX2Ecytjx3LtHnvc8q5c2MpxrteMdS
qqtvAAtd+A3Km2s42rHDV+oW1bWHIIr7/IdtkJmM4W7Kdj0fw9mzycAHc57+MWyP
tcqwT0h1SHeCSWBnbKkf8lNMcWerJ0yT5sRUJfdl6C3XDoBDA1+2vf8tTuAjvunQ
YZGeCMBR1rITAyaLT4kzt0uqqRmmn0maYZbG/4wZScpxytsPE8gD0vByecJCRLqq
8D8vN9z1CIXpAgoWOLG3QUiBfwViR9mcCxJv3M0lmv4lmaeH1SUBeRNE8Za706Lg
YpshkaH03JeMDKpej0YctD2g5u01H92GhG5usHysTOFgCKWj/3facPqMGssKLqmM
xjuRoUJ4str1gDRsVM4eaphitl+SzPzxpR7/WkFFC2mwtG1PHkXcJsmtfkXHAngA
LTVBZfRKWtSy5dEK7ErsUMTTSNzT6+9Pxn5M9w3SImn2P1qpP45JvXw+yKJsG1Ye
E7uHcYdfR3JeNW3TxV6nDF0m6yYxxTz/vp5U9fyzbkIBhgy9gwJpbWiPpCN4ZKin
ju+ARuRAJ5PYlu56EhXLdgr/6AxVIwXFFvwfo9ZA3o4BvE63vfb9PLNM9hawnBcH
XOMWaKC1JnG4s111NIw+i4J8wkSl6KYS4T9xb7SqeO/21F7lncuO+HGn/0PAYSOc
0Ql8Ual9N6mpK9Sk5FeYCaBE1eNJa5xgSY6Or0fHlxqCMByjnttLpL2k+hJj32QY
mNfudT8VYVAyNtvWuNGmIHUsigH2MLai+gr6TsD/945MkwhwsQQ6jAhDDHk4Pww3
mvXlwGLn74EqzRc9YKXIhcdiY86v7Kqfs836m1c/YIm+Mn0+036xiqYhNFqkHfUN
l04d7k20SmHalovKS81+8JbfsdtqxKMNRaB3N+yi4HlimpSci171Di+ALFFcZpzW
yo/CvwWgrIua37TjIDPkNthRGEOvCrNJcSAf9poJxtI652TPSOnEbW449973137M
NgQy4SYg+dsP8hW7PeCw8wl0HUYbNnJd474RNSoKwqzmF3BGdzpITwGpw8YL8WbY
OzPJESrQBvOk/m2P/3MRbfbRWuxyZWopGnnnG5+FK38y2kq/pXvXwyKFC6qhxddp
5ArEwQ/vJ7ceefSWFggaf3jK6KnMxOUC5iMVANEjdod14l9/NXEZW2xh7UGT5qV8
6Q+FjcmuqbEYDfadHGoN0AUFefETnZG24BJIpl1AosgZlG4w+fqI8n4K3OhZ/p48
pH3woO8Gy7v1J+7ykNdF+mQRAGkArIgwFkGDQ4/XEwoclnGv+g0lgpBS/py/ZxAW
P/Xsm1QVndrfU8DlbksDpERZk97JiAQLI8/M0y/OoOOOpqRffkc2Xb4+ybhhqDLb
U92bgmhtQB/LV+ijfrAscg95tgGS9aNroonMdFKCnVh8WCYVxFBuuxnBxd1Oj0J9
HFyktwPHnH2aWICGh9zqRJ3zUHIuMD/X8h/cfEpkY9Hj3Cjx7DcBPsUh5Qt7N5lc
8ZHeC0nxpamRn+e5zjX/QfjWGc3W0a5HAjv95VqJpqjw6q560PkIIMLP3gqXq3rC
wxNRzxVtK57K5x4b4Jm+bWxnwyMljhlGk5kryKUPt1YQ2QTZzFuoidhzkI24o1zq
YN35cqnlP0bGB/sA7sHrGTPR5KHEXdklVS9XfVLSBHPCLZB/9MkelLTPMCpixeGP
TvrTq7G0Y+TBObSEda9G5+qckvqa+6BjTzvDYChyFjYLAuRYVpUedVpWRWkS93ej
WMxH9dbuM7DkI9/srHboN9l3vt6S4OB2rV0NqL0W1l/gUPRyLXvnBTMx9TfabYXW
ebEs1sNBTGkzh8rW33WQdDDOkpA/4pS1xmNPJPreB8m8GCoFfb+0jPcZ2R4B9qF6
gjKMFiwEMA7X4g5uKipHoxQMceXsSMaKuUQtl+2mJsg+WI8AwXDqN17GUgJtDB4F
xI4xzm5HDlDqm24vLfjOMwR1GwaTpCja9/4vjC17Ps8N40N4FK3abF3HBqJttTJL
qyYb6JP11TfyrHkmHkuAmOzl7gyw93lVJSN8eSnK0kGvUtbRF+KoLjslSP+HP9E9
tLtHqj4U9fvDqq2lgJi3ofOknAHVD9Xvm6ivZdeA4D9mxMaFgLGAlQONsGnyOybS
WAVuSbUDr/Xury5G4XHztsiDumh32P1GBOqJ2VioKIAL+hZC8xzi8e6rv9pdufIN
5VrGuW775HtNBUw6UtNokDASWJDkbBEiNgAGJCwKrRKEc+nzkD3Ujx7NqOcHZD59
TNAgTpqVTt27nR4a9RUzVHCl8E0Y6b4cj0KO2MjzLcbJo4FV8NsjnnNqUo92xMeM
E9W/DgJfgdGkeoToVXVQ2WbTzZJvKOTkCo2Adgi41mEt148zxg+5pgPA6eG8xkMT
63oT0VKWBUV/+Ybv9DCjYKC+bYLehXrjT65FnpRPjtyMNu4N+GzOQjcjh5RapYEz
utg4vd1L31ogOAKPGdkJY0WjJNa3FklMPIRqnJCOk9OmtbGtPmHjee1KJd6qL7BM
w8dmizr0LuZOLbYQoQMaNnigMeC4CZCgM9cYOYSTawHf/X64PWV+2VxG/fdfb/XR
wiFEUj5ZU+lcbKxC4l4zMUrNHzdQNNfaemnjt3ERQ6lj1SDD9ZhEmNQAnidlji3u
A4OTPqJHNN9ZKnTQWKvkOBu5kIobOuomkg34OrisZuK2NOqLJMSYmKX2TBXmtxtn
evYas1HSKpLF2fvdojiwMKhdILblnliKZt95gtAJmg9fV5DuUpvTVtiFumM0cAi/
1sYUWvIjuBV3upREbIWLCTLvJQvOrBzZAmbHI6NfkLzd+SX4qAiJOf7DIpiFdOZc
Kg4oWquHEIBAaSrbKX7i+IxtD1W38adsTaGXnkWriCV+H9rLSv5H0DaByKUOGmCi
KcSdB3KHUUEx+GYkLBMoFHTwKMvdW+ybA9elsauF3h6M0+2B3e0nzwHczOAaQ+y2
iADvDp5RvDt2E0y7MdIe37j6vA+bJPTDd9O/mP+RRWAN+KOPShaY2ILu834xIWTe
mlNZ1Nq30R4Rl8N4lqDPxqt8IQfNeTEXs1SJuwz2Htm+6U6c2TQwIuiO2ucs3sGi
J/XXBa3kMVE8gqom9YaGv9jJfI33e5ArmrsDWVFUalLhCpVmCuuMf/mBPHPtQXcD
oiVtB0zPWK4LO/2RAnTKFr7tFkw458U5cSJZCHisvCAh3KBpT095B7nENZGX6vt/
Mhk1v7Mp30JvWB6XNsXwOnzk/rPvUVZUki9QbtOf59Jsh2Qe2AIkVc50euBSe5+6
0GiVvMPZE9eoEMNTgFxcCVIcHHzmPt8NeWjCRrC+ggMXbxRnOQ9yYCEhrExgKFee
0OLxskfmvGtdC/ZHBrmSBHE+emwfB5y4xn49SC2rpkgQxGrucjkaFFFPOSbaDQto
eLlIDNLSJvwJ5Zttu+P9ztRRoyOpKo1HFkKtqU3VTqy59va+XVps+99Vz0bTR7T1
krbHG8yS+men1X1w6kUB9iTlkz508YjehQjExxMbgzNK7HW1QXUmVsgfHc9Gw3j3
oC+MFj1nxedpjosEvD++HWcWGWeOjzOHzHT3D2opX+Ovs9Dh3ZsyBnHsXHYf2OjN
UVy9L+i84GJOXiKkYzgPjAJP6JbeyUD83Fm3/8v7acvK8n93dGW4kXApPnFM8kxz
Lg9nJyFv9r2KBjbvPDW8V58ZKE+yQos4YdZbOoqSLEnnxfwI6u7vAunC+6stXsSU
6U09m5LIWXvLTo2JvMYxw5OIRf8fVIuy8mnd6IM4IVHTNxIlVLxgeBr4btYUHnr3
I36lumt3gTTdEbOuCTasLZWZUdso9dt1pCw3HcUV29ThQUp4pgwjgF8uyEtaZTL6
XsoVOvYJZ5d+eXgSOSTTYFs6V5l7JfOuyTs0QfYoVLyiRBK+sdxjCjub8PLgdjJ4
dG/EsX7vsuHROyfF1lQtpV7lPXb4D/Tt6Mfol8ZaL2vZpZta9R6gkzz83h2Fj0S0
VLB5uH9Z+O/CnoC8199UFhQ5M4BA0Bl+0qCYNFyXfxQi7DYQ9MEPUQTNznyRUPZZ
a5g+hTTA+p/r7kLqvvua5WySDYXBJ7xfRh5r1a0qxi6xio+NpdtgrijAjxeeeejy
U3rOrwli0XUvVS/segcEzsOfHiI0lBvl/Oq0BAr5XQL8hJWcqPPkXSbLWp3SYeU7
/MxhNyiarCCkBYTF+0xwb/K0czK3G1dhoSfEFT/2AV7zcyKPjjazteWMAZlBwMYT
bD6GxwKo3g5YrU6wXr7IZvTFBhi8v5ZeHbwjS7DJPB6Z/Mnjy3ChTz1EI4//YvdC
0L7Io9XvE8r3/Hphi9X/jBdvIckfD96AQ7mf5AGKAkwyorQLQHJxn/ylACWRlbW8
Ht/ljINLU3SBkJvsBBBpB+upngIxxk4BulD2N0LM0e2UQpd6XpAGR3Yh3bHXqH7y
w/675uVV4H7TCHesuZ3m4O6H1PYcyteP/BbTw9htM2juBG5DNBC39PETZC69opWy
MSpJHDsnzW1rRLdWEgHnvUVTvEwPY90wxWWFrCV1CnrXpikigCdYgTk9PsgPxzsT
3eZykcszC9Oc8ioKDNiUBI2bh7o/AHC3qGkR1rbO7sdZw+cGs36DTknkopdTE8En
Av5MWokhY3yRmYs6AAIJY4BC5XabcKgx/1r4/VJ4AJELtcbw07rdGohuaUGE7TNz
EzuWL5JnbIbvYb9zInytwwLWdP2w0ZOtSuLqdu5D1IxeTCsCPmpRJQMNpYs0wHkd
XSrapDdROhNh7qSOxWVC8a3GtWWkreAZpcEvEVv4AqQTW0FiUsc/FF0VNUZaXFMg
TDbOOiY89ssaY4l19mik9FC5ereYeCmwP5fqUmbQ6cEYIOi+T0nVAHAKk2/xvuN7
1sp9qfYPGteYpRAFe1fDd7aQn1EZij1j4ZalEf6bi+jVaDxsN9nRvV1GO0Ao5yR4
9NJrXhKIdw9Qr5+B5bIaG8JnfnS5M7TiaV2qyYVvmSeXkdhC2oSQm7Ull6llmubv
0s+/QQGHb95VDwokkr+iRSWpWIj8SK4AHe9jrvjddc9ubxcsXVXbbTYzOyxzvPfd
tacH7/gzGBRm9CEIXST3JNIcbktJefwpTSGyAUH9j0AjVEjwhilDEL33GpPoN03i
vA/R/l+2/csm5WOL0AGaR8Wa3UYLQunqo9FZDs1yd4a7kdkOBwPtCYgZaCtXxaPu
loOrITzBCd09TZDd8q0KRdyx2s9bq6VD7QA3jOoluaevStoWSmAkhrmvvMtia5gi
B6cIMRnGNXJ8TZviXcfIeZWQPfk/p/SNGQWdj6Sa28EjZ46nWAdy57pvU+Yqqr+B
2/wqF8njw5NhxKna0gmuZ1/4mNW1KmfR18nxIL9wmVF0taPN7gxJXngh8PYD1w57
pPqjV9BTJjkgQuuMp2w7/m8swKD+1Zft9B9ijwN5uibQPmbQXHrrWQkj7M7nddFe
CxZJ1letVUJtIcOt4UfU1V2JiSAMd1m96/iI0gLoOkAiSNILRFKiZTBoMAr+YYUS
Ab8J1LTvP0wSbttLm9oCJ4AcBQ9UTUvsrhFXl5WxHCm4MG36kLsPpRPh6+9sBmEV
Wg2kKc0aGm3DBNiiBeajf973MbQ6O5ZOZXvr9gLfCr2mHfO4i3woLvDyNGK2rIgW
RA3IqmGpgM3XrrEtwW2p8i+wauyOvKYop8DxsygldPA9vR2GYdjOu3+EdXmzTsX6
1ubbPl/ceru4e6vDVBs1PlGRF72c2Trqp8gRANM3QObMBvJgXYCdNJU03A5vpZrh
`pragma protect end_protected
