// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:09 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B/0KTZleMYYecx4HgEHlaz+kWcFDozg2gz9nZ2WLoq8djRBcd125iSLkJI8QGID4
1tl43CGVLISaX4MMdA7NDzwQQovejbK5Crw+eL+BL49r3lOLwTqfXqgYqmTnAXv6
LCi5lByuSUyTaPn4Qz5DPIFK37BNvK/4D2Xlw1sOgRU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 51232)
rmJ5a8Lxo5ewZPkkuiOKeecJ9tt8q5oXXr8Xw2pUv4yZAbLZ31M+Ug5JbUn3GUbG
ZQ9yRVQbn7pZfDCx7HbDeB9NX1GTgATkQDZPFG6LREDptm20GbDcq7vV7gat0qJt
ghUGqQqJQDw+F2wr7FTX0ZLy+HnZWN4ACsypr43mD8mRv3KYOg0zqBs8QaGHoR+c
h64jFOwOnOO+6veePpCyBoR9cPUfqf7SxQA5zikjas6oGGKHkZqBqduiDBfTYVnU
43XxX0muxfUw9H6iDdoBXeZrcJI/TlyhEQH1G9SwpTukdGHB75sMrCP79KbdZ3/Z
28AXAM777P1/25MRiBedFM006nJl/lS19D+HEMwav6FKrxs/tVPejtVsUzaplXLT
YM9fj3IDedVcc6MIRTfiPc7fxMtDRQLAUZfuwMp62YWV/afic9fqmcu68ombf6Lc
rQF7eqMAbpTedsw4b9HaBOdizNlw9wgLjdVvsY3wNJT+pseCJbG5gJNe3al3Q305
pdU5i/BETmeBit9VAUCoJEHWvKkk1AHHtWkhQC9V7LGflK9axHdVkleg/lzIo8Fn
d2BbiiVGMvFzbGJ0VoYDFd5u0gshDwwoARsTdYoQS//Dts5jRtnU6+pFCM+Tyk6x
Bcmg4B9EP5fJ1dr1WPXkajvHGN9oYBdWEw6gvGwhV53WL321cSwl6Ec1c4yBTULt
dA+L97PLalcvDjWmVgWYjS1c0HgAq0MOq2E6KD9HSitCauoh7B3LlQLMO0TWij+g
8dFs8fbZT/ODnqKzaWe/z4AdXQGFUOcFNXocmOZyGHdWEaYFK7DgE9HqcSrjADyN
171s/xxJY5f9fFfGGdt184+tDcVbtRiyY7+xvrvtHGoztgVS/81qbgD4KRruL/mf
18I9HmCvM6aff2YHZYhYAiBXqRSQ9nvVFgAz6J8RASNDqvWDbnM0UjiBSO27BTpZ
cZLix2IQfb5THL3wEYZ7zPTLSsXpbjppNVm/N8Bl9A6R/oKtmvz6Coc6WXSJgrql
gy3zHcf/3EbaxoBrqnkfUrUd/2UrzlTkYsX+HXrkjc23TckneY7a4PV0nlPgZQzZ
CD0XfTUw4Up8NYTzdzxbMUhwrK0mPoZ3lwt1tayYYWuyF07ThGF33Zg5WaMN8+HW
cKnH3cMxEyg8JtLbhpQIjz8teEw8CvLuHyxavp5D6CfmTDPOPQMu1jRodmEy+xCH
YJdU/03zmd4xPCQua/rJbdBMJ5y0EwNx99sVG+D1bj0ZUVh2UDx/iXB3yEZQ8EU3
DxOJXcv/P7950qfDGXb6y6kysvEurJDcIsEy4+YwOD39u/E7/Y21/eJye4URKfEn
2OuQ6CuOc8rtftDjs63cU90OyEAdd0OK7hLkpiQuQVP2W32yriZCoH6fqHsEgENr
oXDTgszyrAaXMrUksPswAqSQK+Ar2cXjPz9o4BBKaUdlfTvUdH7TCqRUDKVctY1j
ero3B/CKbNPQr5wU3hWiCZ8X2FC/SbVriettoJS5Mui88rZLdtuWdi6y0MA55DN8
wuYCVXmC5h1xdBKN9uX2BqLiNy2TE9bY41qYnVKZbsCP/TTtD2rBouOtP/BTsyBI
/ufJmnyJnngxshzYIrDAGIxRXqX5s8M0mwtMh+6MQf88ZY6jCxwgU9CHVqpkTTV4
Gy3c1VHHfZ5+88HCS+xEDxZasdxzX00sdyWDkIyD3WvBbjXQhVQ4JX6gvowcXasB
XjH+aXlwNDwiii+7ALKWvfrevhn0VObNPoJS9lvM3OB98iTdfL+42FHiMcHXzmzp
U5LhF2W8Jme1xbJkUgxfjaJkZpcIFji5f4V0T4yI7xczg5e3WsyDCc8WIuElBtfn
kdahiidFmv9VxWPPPYNs023DfJvOay1Yp9Oj79rU+AOJZHMNX36VeaCUa9GQ6W8H
rBDeXFyp7yVm7jMWAJOOmFX0kiviWbFdcBq+ev6ErIF+EvxEYr1MsaOE7XGE9MEV
qqrkZ+t7iJ2bj2fekVTw2ftEF8VqZmwPC3JzHhW4q3Ey33X0p926/HhqOZvjPk1W
F7iEAjpqjoFV+Bs0tCI05CqCBLxeWRizsRWI+MuvVU2zhzxSftD1dV9XA3eU/kLH
ZLPtsJHivsS4NjOpdgWMgsFgzXHrf0Y2dZ7H5J7IrDimlRK6cX4xQ7caRx7ioija
aPpTPHaC+AWHr+QjrdjUtOWvSNkn9s2JRshQuZzEr+M/WjinmJ6FSJP2Hg+TH5PO
tj1gpYf6OQBW1kW403qElVhE6YI+HWGxYfskAmKy5rKwD1aodVevmI7KN5+1jcOw
UoPzVzUQQbgP7QlG65LoLt387mDsD750/rbe9GESvec6Oup9Cdzj3Iowhuz/OHng
MmrYlWnIhU3gGQ39OJNi4tWSH9FImjiZyP27fntEt2rzDg/fm5Jr6OoGo2+xWhyF
ClOJBVxvzAalleYFClzWkLjCO+P0AMdYOWuxX/5kU8bvOPf70WLTQK2MUZVdTRTS
SgNSyWi69GhkyHb8gHP28JPyMSNQGcxLkPPRwyCYTAatpgZ3U+aFhIXBlPx91o12
K5vN/WeUda1WMJMyXVhmZb5gJrpdPsEJYgfegk2ytLJXtQQsnefn+ZpWvjAWx4fH
0qMiIi2o7T4jIFriyEmBQsjtMXNOL/UjJ7sMZTQQ8Gt3KQhdm4VqzokZiXnwMdyb
n5T9on/SVt8aWJ+GlYY7TyarmQKHiVLxen+k1AKudJ5A6Z9BKeVn1Wje8B1qFAku
Zk+QmoTOex1NstgPpQRsR5v8Z6pTDzcbABDUAHlnTZD7DRu1oiOGPHrmm3PbnlM5
CwbWFpWCIrvOq6zbaKtjY1rKlKaskEt5NHoRALPnQFH5XVeoFljp7U8GBJmotfAY
VHOtUsAHy/CJPKqsy/Jl05diaoucqjhGiLJvxah2NXtw/uMCIf9w5TPw+fPtLzB1
C1otWVFT8N+ltLAy8Q0E/I/hSEhBPyeu3Df1QG6Zv+y7kLHEL2Joj3/TsOQM8LXg
QXMj0gVLiVz4kdn7LCqKHEv6AvalvrR4jG9h8chjdYHQsbuYMCzMFqwR6xSw/jlf
Pjf+npzTxkGMq5Lr1tOZ9l0ZHz1kaJmp5536Oh6xxzT+ahiqsk4+5ADo9RNWD7Uh
caKrdCqQaNNN7nfm18T0oGNNNXcIeBPdmFw84NuIQehDU8qQgqGUGr7dnoaLk1uX
SLUn4MPoEte6cVyHeZE2sWWHIK3cHualE4HU75CYBP4NlcvVYq0ISaYE+z3felQG
mo5x/ddexTen164ihyTCnsywmPnSf/IBacpgXNn71+5cP/JvQKDBfWWg4e9pPy/m
tDxZASr//LpH3EeUvkI6ytgN1+m11OKTP15JELtIVpkjW2OSrw/0vqZk8lU7PYKK
ftE+7h4KpHmmRgwznnVeFsOdn+jNJ3idMplyqUoSTbEV0YGrS0IsC7W2Eyi+dl5B
ZUnwa6heYTeRWDIG/C/DEvmuxnGnQMr59Dn7rLGs3wfoWDGAJUoJUJkYF2+foKo2
j+jltrlTPAKiBn9KF0uQVEv4cwfZU8z8NVnCzjoEMwCv9yHvnVNoSfXK+4b1vN22
gWRAkdwJdBMiQnggyzHJ5Atwf1e1+5x7hOhntt+glWGtVVCrhhe+JrwC3rpovbcJ
aS0z0ALh9FyssDsZMcoxQJbVnSYikl3ADHX0qbEx6zRS6XD1ZC9yGFqLb9Ldu3Vt
00g2q1tN4LCN92wUORJrgBMrd6KRrI8YlC+GP9e4F9C3oRN4889IL2l+Eqw74Ke5
gX7zSrMlZ3k2a0Y8Qtrshu4UIYmJn/HHAvNhtBHEgg5vMkt/xrpfJ4bjQFV2uFlw
0o+BJg36mkvfv46Ba1otlTRAQlT13ZkhbGcHU8DKw91cy935fjM9YsCLqsFooWbM
nHP7Noy+JyLuR6iMp5+UazHFyF8ExAN0RYwlfXQiymXquuIRS+88JbbmeMYWifTe
W02u7+VBSUf29x5dTY96toEAkGCXOBwZyCO0q5BCmt6spIDOkci5JmqEt5aH3OIw
EXK1waWQqruim3g6VmjNJnKysPHldxBtdvkQ3ZLMAVeSMcRCSJUYp7gofwd6eSO2
ffT+rBm3dIcMZP0Sah76l4EaVRif4/o63C6yb9J97sEFt+qYA9zAmuN+iC2l1cWI
rgU8bShqDpF6GZZyzhWUn0Jc9RTJ5EJNhnk/tLa7vSrcUR/e6a5bix+FEhqQ20Tj
6nlRHOUlC2SdGxVmgnL8eq1WoQMJI2ZRB751gh/o6zuse/mui6oU6LLgtvT2hpzh
0j5NYQpITGHvSa3J/KqrwrY9tugar+igqpIUAQokb7RCELeT7hCxWpxROvq8nhu/
l/VFdCti1VgCPQimWU1dyHcHuET8gQucb1JtSl/WRuTtQDezzwgTuudH8xZIdyz5
gJoA5De4IhwQHovIglrJi5ckRDwbr84nXX+HQOzpTf87PGcLDyejK0h4dPbeJwYr
5uJDaZGYn9jdfrMWEG5Wt2RLVorGDLVu/+XgmOxM16LC7IjReI+6UdFuOvBV5fgf
1FFbUXeaPLEuYVi7usOGF+wRMqFoQte9WpBjeyUMZYLCnnqwH4Q4Bd2w5iyar+8Y
gwrBJjWT5QfdO8W0bLtwJho6UT+s9dzbtBTbE8U6a2QgATcPMAFyqTfXO9O+QK3p
06r12KpH22zRMrVlSBm9ZyRkeS+bckwVJQjKXp027fgQJCTAPr6+rfbRZGzTeg0E
4pdXLdzP8mIDzi/dK6e8GR1aw5XxIc5Mh/Vwj5sKn39alKDPeQxE1LHZXjwVR3m9
QwcRGho0uNBVOjGYHSW/sYmDqyMs3SQBbhEooZGRTdE6duIZz1ZJzrIO2lsbk26l
SaZD+nFUbKvIfxHbZbYZDLTUGi56I6/Z60mm4104oVCLsJmzaTBt6paD0RuTjAvH
2EdPKmpArdHIXFBECTlCG4WACRmJ20NhzwzOkQWnqssiTIBrxsvb9a0gZx7mzLE6
5i/+8h4nX6JeQZgpJEVBROWn2yDwSfELlfCOvvX31SkgW2Dsu69aCwLVy4/DiSm0
sLFLkqVlYWM9OdnP5i0yUj1gU1db/SvcYn2rJoevWxJb8WzfKaqN9Eh44+aS/H1P
QPnSweaqBJayvAdM+AleDg5nBdNMeOp52wIDc+RSy/TQHu+TW12eMPetkaE40Pr3
/LipofTxMX85HKRu7WjmbOdDn71rAwl0QEluuc5YqFpl2X05S3IfI0y3ZrZywqWj
4VxKoh0G6e7Sp1wf2nAMU/fI9Xb7Vzn5gOofVcugkyQ7TC6tR9rZIPzT/LRa4YZU
fupHowfnbYA3tfzRhC4MDgePkRKtbQi2sYdrAUEAH3uNKOxn9ugjBmvXnYABKme4
FR+wvlDy/gYDPf+rLI3v3RB34Hn/USywlS5qTwwck7b75iJ6/P1KfC8FFdTRM6Jn
YVzHWMvz8DhmZ75f0n4T7D5a9B4Dagwpv0Nns8NJ6VtbNEdBtVO9VEh9FAIZjapw
JCtGipHaUU5PKjxUSMCJTr5nFRDGDtBlYhrSAhcYs9BFnNN4nduzRUrc2d8G99/P
u7mNryoMmkR7YGuWuRPWsyOrF4Z7MdPbjLiYtuVGcdRMpcvEQBxm3KlY6CxkafT5
isHaA8wrA8HsINWOFxRIkIcLGNY7N9dga6cepdN0jxQ0nMnLIEgAqI5Q60eyYf+l
127Y/VA7RcX3tUuj+Emj3GsQD9S6+MDvgyvbRnF1YKVDl6yoPnsX6rWSGtsnIljl
5c5WLyKhKf7s6okc0W9/QfW04zyHTL00h2E4Yt9QuXVGsAxBz8dN1VpFxPe8MO0k
crcvcbaHJriakqngiOu3tDTqEkLRHFaBAct0G7LtqUrF0RrES6iWyxbcEFFY+1e5
9in8r5DQRxv0JAe7AnWX5aKYakeWc9c2L6JRcm6TAxQgBFBRfdhnjLrzqJBozWtd
3PvIGa+L6TRrPl/XGZ9L3wpDSDw0z6Yp1Q5SwyDRR1L9YOcUfNL4LGyr/j3aZuNj
Y+0y/+4AeGfETAIdWSg82KjzILxtJsiNLpA9NAKEtPGvL42UYjMy5g0M+xW/ZNkH
un6oHW/MWaz51PqSex04iA+D/3SQ9e//2sxV/jCDc72X62fQJZidB8J82gp3a+/u
MZJNwznje4aDF7VC7NZKRd96xs1teQ862q4i5mv6KfzH2/y7yov5D7Kkwv6Ntjfn
yzOVClt8dnQOYZFFIckM4KzoWRsnsML5eP8zlRZ74tMXDACowL3/fqzy/mf3/94g
M02z2RoOe3+mpt5yxCjIDfOd0YuC1GB3hpYX67rHWJ4svHerog/kMiuIuixbPa5K
Dr/30qpDFEXvJLYne7mMBukuLbtoaKuivgviYN5/FL0SjgeHTsAOgCESSyyxJLbx
JU1FEf6T56pcz9zmq2hi9vVUJAlEOCuqSXYh8O9A+zqmFRybpbARCsAjogJt4vky
FheFoRp0DQdk5l4URYEnLebhc6LkwBwjznG9bRA2jGKrO7cDkNXgD4gd1UoqM1/X
FDKyvgLU+RcTFDpIgPXzq5EEj4SyP4e3/fofvoA+WI8mTXF4yEAGawA61GqsmbkH
iFTWmW+c6w9vZn+zv9VFt8TD470nd47AvH01FiYNNa7FOZ49Gy0Md+2H2O9P1uQk
nbsjeAYdeqF3eCk7OoQiFqDIZOcoX0p+buvZCrHZoUIRCRxDXaVZvt+XXIwFWN9n
/Bam3BarQAsCuyRZQA27Zx/MGEsmnUbWpONlndw8GfhORyhpkHAJGcL/Hckag0F3
YdgYsiKb44fgfIsiGGseafYS9D7nUMHZcWIjB9ojCglM7psYpFwoN/Pi/UI7YXHS
4++hjilOm3yXbZi7/Uy3nxwhLuSlhBrE508T2rrhLYxSnIPJS/dqhTSkXayKIGvV
43HoAESH/iJ+JjSL3Jo3uL/G94Y7fLXCLe0pbsZv01dDIHWiMaAJrn81Y34aEexl
9wXzcJRkrW2LGxnSOzZM84JlQm/Ntl3APBbkZYGEZPczQcXvi+Iz8YNIsya1D8An
XAAucrFZK/7+mIzSlN2y7x1SsF7kmN7cWCEg1iD0a/6/1HbcRuZJQaMJZFUDJu3v
8BqYigr04rMCFSKzveYsjidy/xywmGg9lAnv4gBSOD58tIj5kHrwrf+HfL5EBBja
Jr35nZLQ3O4MGxLbAZ8CyRXUHHHNDDp6WLqjHuA0oQQ8JpIW3lfMDS66yo4i85AN
AziT0Cx/3r6HK3XsFY1MubWRdOP3YumBKk8OIjnccjoybGMuH6UQIePdyzmhGLQs
5585mp0V2r90hI6oBJUPpECC8Pyq9yEEcnY4aE+7dmwbiMcqT/9YThNHUVyKFY+m
k+2QFNzPLmPUIeTJNXv/jN33XPRHeLF+oqJBCgXGC2jQMM1r1T7cSW3rAOIWTstR
HXvbaOefqd06T+TSfVbcudB+roIIUkZARagorMV8Mqiff0SpCfbg2aadutOde+mb
SIszAmnB6lJtS4ziiSPEYI4zcqMo67pK5Jc/JrBR1jenA9Yp4y0GRv6XL4Zx4xnM
SJbxNyh7HI8heyk3FtLiRl2/hE5CcdzJh/M1CTKujlT6jIPIPAWkl7eXZHbnyc0Z
Jc9RBu48gdTrWosEgkuHVI0jSkNGnjok0XRPZ/olbr2/SoswquZSU6B1/W3JGQah
IMUNzhEaP2XFliECtgCOYAw03bVy2kU01x2SbPyc2r3/Fww7UQ0MlxKwbtVquIBb
cW57vIIy4dJLqR4jct7IroH/6HusRIkKR2dgui6OOJBSghVoYdhEI3iaRZ2Wfp2c
gv26GuCcXiK0jC0AfZdlYxC0cJcXe08J7hTI7miHlsN58iSKVBb5K7yFAxiwANRw
pj9gRLXgKmc7bMmBriaCcyrz3Nw9pL7kq2TxX3+rOHX0Qx2Y6wcw8WzTEdstC0U8
uwRAv0oa90LBS2MDGXXS71kACBh6p6qOPJ5cFQIGsE/nTAEClMuy9AmguypdhoVr
dT8sJYkvKgOU/Q0SlNj0KKLQg1CUJn/FXuYFwvAyCYwZEiKX8UVqCL9ualYoM9qU
LPjnikrVFUs46xRvrZqo2dhOjg1yGFyGC5kRx7DejXj9OyOFhUkXicZIetwiTrX0
L6MtS9bpCNn5BQLkQ/MM7naIHcuQBg6u60MCgJ/9w+ZHqcfZKz2r4QaHpDEEZN6+
r8+x9xJOZOVUIaqWpNYKwIyP2UCpF09bGjTQgPO0TGzz5B1L4sn9x9mcVARz3HTb
d18F1mmHHK6WWyxgRsnhdhEAijCKu7IXhJtaMaEnSgWyVV2mTmzK/ArRQPZ+SAgK
E0cdmxewVpdz7Q3wHqaxdQGxaIfhkQFykhOwBn769PlW7EgYSQvto6udld66SObu
RpidwO7dEH+ChH2r4mmJRS3F/6y8XAEUcTam0cHNDjotJeMvXYNXcxC+LvLqV+q5
64c8oF89yeT/JxUXKipjcda7bBZmEEd6RpCYZMQuPqHQJYhUsY4wIPzLG7TWcLjW
rLdh7jX9fq5g45TzCXfi8TNAtoCIJeqyHHjVGgASfiRQueMy+ZZvWBJDKVR6T9Kf
tRQmmX6A53Zf8XmqBTxyXpGUDTMn3dItrIJIstzPosyfElMuzilgbMaZOEeI9/Ow
bZjG5yHkQiNaJ4xALxTCE1339gjt8cuMcQ0g54gOQ15KPQhx3kCyIr5HlsOsnYZ5
/0hR+rUD3XYgxiHCJn1JrMEfFTrDdcxSWSjDnZlYPqG0YF1/h2+FwVUdSrTmqinO
5PungcCy2Z2uSoEnQAOd4s3rGD6yIi0qB9IlQxu2vTMnH+pncDMCs3PsHPJIKbol
dwJJj+Bs0z1aqvjE8tGCeuTjdBW+u+V/+USm7NOYos9yhSptiOiOF1IHlP7eDUX/
+we5fTsr9nP7aopLVbzaUHxLqLD0qEJgUFw+HmhOWXsGV8vE2oVM/oYPzRmvpF1N
ZJ/pYFOyrCSzqWqeKggHeFEPvYVoxJ3KukrsQiC9doTXCqrtqmTvOsWY/lIveqNG
f7982LlfDWzOO/ifzg0acEcF4lLS7SNOQa9EDOrxu7eLio9YaxEM42lsJg7qtTVA
Un88/4gfTFEHobCXhnhhWTnOyKAUufyuS03msmbo/m4WO4hvQ85nkaXtZZ+73smw
twwdpDt02qK8hM/6CGjacFWXS4K2dhjXwh+ISBABdpr8X5MdtMvrYJPIZDsp2R5n
O/Clfm7hYa7vJHSh2P3lMV2dIuk8CIiyhe2IGRwzslbvqawV9Kumh3VnU51kbvMd
pBRrGrntqyIJ5E609hQLrx0/8BQvraldb6nZ3W1giINNooJ0joRQ6zra12JubAhp
FbvzDlsuwXsX9IXaaHgJwEXMT6fyyYj7UnbBp4XKv92SlywzbljIqhvvOlsVuEuP
mlrIF+w4FBADCm+o9qf8+hWmcErykVECXO6vfVT5OXOyIHNOZgc6SzQ2tZGGpK3W
vCqPjqyyTK2XZws1c2NBlpOxrXYNr9xD3Z8/3lEPJKifYNjSmPH2tMja1DcVT669
lHEwcoIFVUx4X6lqC47VmSNvYk/DjWeGpELS62Thn5c8/J9gE21cQTmPMAM64QyU
YzFDZHMDqAxeJhQNJsp2PSnJ1T+EH3zxgBF4YN7RMRW5n0pgzPbCYVg5ojXBh08n
T4D8owkuVZ/YNIcVXJ9cDIxawYOl2x+3FSDQ8DkCsPK/ZotWiytBAZ4BN67L6+ZS
qhI2UW0syRnLH5LawdemUM4yEHc21lEwNtHpi44bwxoNBj8GeEevw1zlnXiMXHdW
tXhaVKFAJswS0cf/ftvgHA99LKZe8z9f7Cb25Ty1F+tChhM4sHPk68A5OVJONU1F
LUY57kzzdx1/y6LDoEVsbRdaD+orfHnPgzCtLpOpvqzcj99Yy/UVje0UzDUo3mtL
unThAzM4m90Km1npyUeJo3iEnhe3TMf7QpWImhnuv4uo6NgHjD22EunDDhAIl8cd
tJxQDVz5hCbfWaEfespz28n6ls62+Uow1hV3/C2cZKp9NzP0DWuET9fjs1BglrIn
by6V1NnsmIVQAlBOu1nMFnqykosSzI1cIIaEGKuBFUYypt6QcX8oepmXyFfzIeiJ
9o3Q6cPklcclybo0LEDM4G0Re23SEkwooBkbtDY61XIsWw0FUmVkFzfCp93pLtV0
Re8N2GV2CWhcA3XQ/dM31c2vqcnSywTy1R657Jlwnvmr9lfGW6iZo1Cd45dwOiH5
Dgmn5MqEbnz71ktL5jl1Pj0oNeDkfTgbKujK5+2cRYB47rpgXZIPI+rTo0oRLJ/G
lpmgoHcvAXTvOMchNSDy7qZE92VtoECScFTX/Kg9WltqMmjImJZQK3A+rjpG89Eq
AjWd20sLVtz1S0wySlEhN8qe4nd+vKn5KwUfs9i+mPkxDHRsN1P/qZJl9M5SMHh5
bWOpmpoo/m22JuBeFipkAw5ebly03t+CyYZ1D4yvXsYMqpPIc9yKY52EsBt9S3Mc
RS2RLbhlWbu0COffPPkY7BwPkrCxEq380oRAvjjDMGOf3sVyLZIpl7+06pDhMaEz
mZp35k6zboLpemFRYPoYe33zHssfXlP/28qm30KfpTjtsZ0aKzd3uEyxhFOWntn/
0A1E5+r6YL43jJksrjFQN8WkV18uVfWvYocpkXkaMl3VnfBeZU2oXRZk/LS0Mmlt
3GNtrQuFd0DhhtX7uB+hHKt2cboImT/kFiiJFfNVYrCw69PlkrgD/WN3orRdo4ZB
WLoFH4WMXiVbvreGvmNLya0ventsrDxdQrq4xdw/xxYKOu2DXJWW1EVcPIJuPl2h
sApa4CWwXkC+YEMz4m8ni5E192fCNmd9pJXGCYUnk5UPa8jHtmplkti1xhXRZkta
K2DsvQrw3Xd/AyOfAQ/jVx6GPDaLLDvNDEsomvC/2lYqZiOK+sbD+dGLwn3CHmgJ
r9O17qXCQWpdUmfU5XwFNoad4EKkg9l45ai540wnG8HHecfffxk4aD7tzF7BdFMS
OwR4kpnzbO9Skw4IMZ2lLHBS/T6DqebQ3nXQZbKcnfYMRTOMrrvLJEFKFW919mG/
aNHJmSLXPVyalNx5ZZo9jRQAsK/nCue2CDKRpEo9OaVgpRf7kEnP4SBRKfwt97Xc
zdUjfucoLjFBcfYlmC+QeD5ThqcwOcXw3MYqCT8zFSTHW+umTUSsmUcOPlhc9lj5
VIgjSaqzdpD2HFWBpMg/ed4ZT4ZOL9/l7jZ2Ovbv9v4aIDuahFr8mrBH1Mh+DaBm
Q052bXxw/Wi9WMrhcuL+5qkQK5TXbRzqNqYC3fMxS/QoFbVRN/3ndvUhtpiXUJLH
y0pFaL0AIR2OMr4moTzAYkOvqtLELLZDD87a7BMvJfS/WDQgugyvPH4XWHb572tN
2pAMCw+Qao7v9DoVpJ13F15wQqPjOZZA1MgaATy4lsLtmgIdM3IRCNDvjl081mgn
1VOKZ4OGOj1wahl/aH8MLDZ2D3miojF+mvNyUGrsVzI8HTxhdn2PYYlDfCjgezHr
AHggII4lb4QA8PsjbeeUpCJl568gRXsZnnFtI3b850BSrPrdjYazec7TNVfZ+Ctq
6TLCIW6QzKWdvAeKD0w1TdaRX8B/KPPsrqOyQ4eFn2EZYIYg0t8/I0CuztDxN+k+
j/DJAoX5xRPMZKB9FJKrlLw6Tc98t+VtdjRWZvAtRs79UBjjPOwnr9BvVOZptL9T
gaAtsbEwYgwBnip3tCkT8q/paH92KnFKtVDs2ux9EFzwNWOz0zScFPw8gM6YLi3i
/gAeNqcrU0dQIqE45VQ96sNYQ8hhRGaAuACsXBbcz2ZgLiFjCSSwJ1kwhdGcq6X/
aJLAtXAqGTBfOETh7Cq4Ew56tf22VNplQBeJgv4HlnofaiPWXKIALfFzT/XA/dl+
26GyC+ZKR1KjZWvE70DCv1/z+SSoCKwxR+4gDBk1kfCkedcGe+l1vf5+N6F5nk/8
KGYH012advIj0o4akHj+SdeEQsk+XX2u3PNO1XfKz/HFdJHjxX/wxiC11y6PM4JZ
zDriCII/EIQQsnejDhtDoaWmJNn+qPrmV7CCqauzFnLEJWnUCD6cD0wg8SSQZF80
pmi3wbMrLK9Nfz+i4A44V2iFdc71mebwO7XXjoX6uS744jBFTVWtUtu870WAD3vB
xgLkFg2tahvgg2PW9pX8M8LnaappKjh7iV7MonbDE2FeRxWYh89BgS0qyaAAvTLF
Nv6GS1F92nfdUNoSFfyrHhqcosfqQ+OaLcXyFaLev/OwIBx0lYIJrq4oeWbki9K7
HgL1nI2MxPFWI4ma94dN/96/VIUF98AiAaiG5zyNH5syQhnVH1Z6otWXlH5llxJ3
Df7s7/OtI4pNHOM+u/kGd91E0Yyap0BepGI9Yg9M0Xd10Cg3KvIvt8aYuDpG2pAF
8KeiGLE1NcscTo9/C2VA5xvuX2dEMa4y1+RL50/+yKf7at1U+IlZ7I0C+PmvvSz8
qDebR+lsi2Z0r3QUHwzAaYSvFm9C7xgXVUOveYohiPovuVnGw42EAaVFh1XPRVL/
jek36iO0auV6p5dqlqxpHyuogSxEp3BmlIiHBf4RkePkZUfo2KgyCYmTkta+ktN1
NoienZVBsi+Vu6JrWpvTOkmSGAq5x0EVgIscak1uEnRW5r6EmqHXV9dd7HTKQgAe
3D0arbCW42IAIc0GzP+wm8gIAZms302zmgNaqsStqBSSPBMEQ/N9BqUY6PPSljbz
21qyrXuJbSucv0utiNS8itTsnDdNXmZsxD0B4lJor8YeXoVMcWyOtj+HxM4KVcKY
5WA2G1XBkim9vAGmzdcJDzlhAn4zCHWAyLzIAMXoBx6U3gizUZ7luw6ZsdDlB7j9
xNfNMnkVX+qk+a9unAE/HyW/3dCGpIA3n7sQmq4N8EOTLPiWHaDi+3u0xsqxnVIS
JSALA91NTJDpJ7uT06FGrQpXS/XCVw1Mh+W6pp0SsAuU46Vo9E38EbtY7Q64qugl
dq6qfunbH89ETtkzriWpNdGXpABNRb6o1HceXCPy3KB1sCLGo4jMQvuf126DpFTw
jKkKayJnj88G9lqSNT6xY955RjJ8jnzxWimzzH8K3w9U8K1KVcovTTTJj1oUs1FP
7JQyhd7qHSHYfApvUTUGOZja7p0TCuXS33crvUeTNHPwmc9JIZtcBJQuaKnE2wOh
PlDLAQ6lWp/zOkXgAqvm9FBNfvzIUJYMaHaZEj6sHUNYS3xASfhj3YTUWGck8w9K
xMvrvhWTPNYsALCOjFEggYAp0F+2cn5oN47jvg1+AnE1YURlXQKSqnroP0lIkvZP
Swsv4DUtX80OHkDwuTRn8/Z5QbqOx/YogxQnTZHXIO/hBa3JMeWIWpgxsBf8Cq2m
FqQq7y5QAU0g8Bmy4yXC/uqUJd4VGM+c8AGpK8Po1H/v2bTS2xs/nE+QS4uVQBZL
KxDobdFleI04LS6aTZ+P5r1pXOb9bumNg0Cnw48+ywwjn9M00nWz+GqYIORv9iOd
s7omwkOE8ik5BotS95uojwi2JDf58idPNupKrtt9tAmyyZ+VO/T93Xggt1F7NqZM
FLlXUQWys2MZ6/+0kifnxunMOlqix23X/0+OawB3mPhFJuj0yr/EMnVO7Ro6DUs3
iEkbr92Dz2Wnx8qvgH/EXEm5vwdsqdC5JQZdYfWJ1Kat9irIeZkSMbHKEUKjj4Ot
LqtuewRkOOwkcnNlY7S/prWvGdoek7ie2oUt+5aOviBTf3VtbpuKR7E7iYbap3f9
V2uK0fjPCjQ7o3INEK7BPmbuFJh9sClaqd5qAtWgn2S6ml1035tzLrO7smtfkqBM
p6niEighKh84TBgtP4j7s9lsfinO8GM2PqRX8X+cyFX3CYihofyq+Wub/qT7IGan
uSaygewC6lHee7MGiytlIr0jo230AQBB1wEmKuvTGIPscf2ytzqMN6cStgwx9tMq
xWSruemTy5mcq0RoLHCsrn31ZgEsMf4rD/vIrmsdDorBoqqgvkr0qkh8sCP2spG+
5gPVXUdz4TmMGvFv/fstmygg3YDkorzV3d0uwiy2XHqzKbt6m1IKcKGS4B8Y3ZOY
Rbf3Qm6bF6uYfjB2BO2c4YE0T0yPHoLyzMZFR9hfHOYIIwlRRRry39hTlRkIFS48
0nKM0SHlDKXaxhBesJzwrrUtkEE7fE4V1m9Ql77mlI6hUELRBsTdNdyQI74ivxxw
TGkp2EfIE6c3p/WXBOyikzWarPLxrRc1xiJp1y4sOVWND9SJX62JqYW3BIokl2cV
CdJJZ06FBED60P4H/i8OHavgvDyKoQXz1Znpp947mXLeCB0wC0+znz/GCWKgGAld
5EltE0VmXKzngiTuxhssXaBmL56vhaNAaiKptBrDftOn5UfV6KXOA63VuRNgzL8z
TxdLc/JHW/iuUXmY15VUrmOcFiXcroiD5bcKXzTKEcQOmWpKQkuNC5pF6Jt8DWKc
OoUTbHABsPCw86Kz/yjIpiB1Dpcth8R277RyP/ilFLINqqmwdeXESrnZ/ywXt5f6
pmv9wwBfk80IYAF6IKMUFDvkns+eMHZZ81FJuQmNf6oyFQRiOIRQWrbca4TuxNP4
YFyd+HrLUiNefqW9yA6oCKa5jtHXuYvE9Jt5H5rm/0j7oZ9bZ0PIfaLin1q8ok+m
Q+ZrNi6AfOMnM7wuQ7Qqh9Bj20qNCdt3BkVsjwrFO7X7xdLGPAljc+Fjx+nAe+N3
83jT25FZ5Ed7F8c7tHdUSrgss2yiU38HKss+fmddhgiJ7Do9hsxighUVlu2sthmJ
2PR1hS+sSSa7wDK9LzvrMYVlBW+Ftjpl0CJxHM8fdPsP6lQfBXuAjy/dNtoTKnY9
fwqkGDYw6jkWsain2hMHgJt9rrX5GgIy/Hwreu0y+DY9FGtuZTPcLoT6TL/lvMWa
ovKFuE4owUV3y/gTrZezH1rvxBb9FsMHiw0Xfn6tApJjf7OKIRDG4ncfPWSRKpar
HGUS0d0hkbWbEGf9BBoVuQQSL48Cn8fbFoWm7IxlqqIUVa3p4g0hWjSEZl7APk3q
0F5LfE4wYZ8dzxWgv7JJnx8kPaqzgH5fOOPzXlYubw/I0z/HI7TyGM+EsqKnQ2ee
8id5MiBmblEwCK482LRRRFMFCXVYGJIrr83y7VuCJ2GF4GEpHP59BeL6hYZ1kU20
fOr/r+LbsrctM8UYgjxEMWQQpIvQ5i5iQi4tzNf8Mm8cj4sjFIErc4M4zEbV+SDz
eKrSEPgn5k0Igv6delP/IOeZPwcbWAwsDjLtng5JR1jTw8AGDq1+hjhK6Ne7wnVL
Uh7R+VU1l1KPV/o0ONK4HoRAUly19jG9tnhNV17saP2VVR+T/Gpm8ii4pYPSPIXq
qoJaOcQJEeewG4/ePJQ911jLQ5gdPrUUc34ijBZj4cjWxVRlL4wwFrlT9X+YMR1l
efEn4gTkToKHCffWMESAkepHrkSEV2cM0xc1IjtYRMQu9q8VNNbNlb0PXZ6879Ib
oWUIGiViWtUJcw5t8/q+e81xdJkT1/zt1sydPU/e+n1zTGb1xzLQmkeN/aWYeaa4
702XwyNEpTYbcSjABO7OMhKeiSBZUjn1JOUsrgy2kYmrDWD/gaUtnPbdioxWnLCA
HQbaWOlGfQZX4gM4wu3QVMI1qHYt1C0u/TLSSJ5iyOwoECKytPEi9cjrG4t6LNeO
QCEegNz5CLnR8KVb2Np4EErAnF1P+3Px0SYLZexekuNH2w6uH4J//Lj15BiewbUH
0QFjLhw+q/hEd4sLykQZBGkPbaaIq0xsTlwPHvbyBm+fikXEQ7Vz8Fh1BnPot0LL
JVgNiyB6wMZVl2qMMdNJKFM/JMN8RsSbw6enVCFDhnl5Snh5SoraoE6HapfQRSUK
4wkF5rTUOKcb2h3Xvb25irqSKZIVfmkK684pnIL/yGbYYJIoxiuQlz4ViwloqMrq
OE5Q//iNk5vuLyB+qV7HvKBTaa2TrjAkGDnMdQEMucx1LaAfQx3VaAph7WZJzGVq
sMfzCS5f1uihc3WejoNkisxBBNCQdZv83fRRt8PfoTHbNKLW4or0H+XS3ZDt4Bmp
FvdidbQgwzM/iZKG9mLifjpPUAbVbMbFlEfoMAN3CGHU0FuXMPtwPRP207HhfZZE
3dhSML0jAefkZjqQh8Pvicp1lCS9VwxT46amLaQ9VzkORjVZt6G6W+AO61TBcHuK
W6yoNl1dlAzuz97SDoApd7OdKZl9vIUlM14MMwHx8XuHQfIdBGVb334dpiOy3OIz
j+/YP7dfQc8kerNV1t1/nWav9keN+7uOilmM9oCJ5/UA/xvYSqU8Nrn5DXcrJVZI
Ilkg+7ueFxOoutoZWQRj1jAyeX9UwRh1+Al4MB+UScgw/XfNdkkYc5uXYd5tjkEd
gRhAMK0R6WtVWOihCUXlxfWJ2hksuXASA/9hV4qovz1kFJZYcV5ww22QR97CVhPs
WxMLWNSUIP7UuH0oOQwO4GNDs+uv6TqXumCgWuXX7KiF1LSHVPmVTNylwJxTlWoI
s+6JNJ4bScHcA7zGuFninuTBMt097GsiuYfwngGInoBQ5y6JjieCv08UjzCOHY7O
fPbE5+qmyleEmsvX6r0ADLGA5/B/SrX5BftcWLLtAdD4x5SFQxYvjk62pQcRRdw7
MgIbEHX6s0Yf6spFwnl6aqNERPFjuAENkB4tCVm3bWxuSWixTRr76/B4UJ8rSG4u
FeQe+WmtsJqqHsT5AGBAohDccI2pDUoMP+3lnf/3b9ID22MesAnItrckHvJccmkD
0saCKUuayglCbf9g6EesB69NnZLR6aZc3S//2A2dkim1GQGNVyjCIw7ToaKr7fXH
RMfVNe1vrQ3KlbhOZRAIpbWsbNkYxnv7GV1m6n3enC9pNz6vzFxpbZgGFUFk4f9K
4bKflL4zwzbrtaFP1kFDp4Xa1SN4FE7Yw1REl6R5kSasCXmy2nO1hz1pK+Wd4Muu
RWIvocCbMf60W6uRjNHW2IFnPIpYVAlHdkOsZzKlGIs7X9t3OTCmG84KNSxLa4DE
FzfjdXRCcUrYgWIiOAEQiZIUiWbnf0ysqRNOOzuuEddRH23k1XtDyIxEfGtgNY17
WmPKjZhx3xNoCEercNv/OU0jRuEPuivHH4U8EJ8pbZR771TLAuL5Sg3IZ5jecDHO
/fXBkZKvXhOOQ9A7mVcf9Mx6sl1TGvfbUHQBiFRCaU3sxA16wXeJMJGneuVqntYc
SC1Y7z5087X0UBnW6KDJ7LlYL4vvE1HWxMmMmswksppPlKaei3fni5Mz8AWgLACu
W5F4c1IlehQqrkcYskxJ6+O+iSqfGTtzsAm0uGftHQhHasyYWKdV2X4PlZMNx4Dn
AID5rZs7yH7pkLiQ5r/qMUzLJVsN6DcR95sdOVjAtdA0uz7a7ArBbLANdkjN0O3f
IyRIZRZhWBzGrk6qVk/ecwTwdH0RRIiwGn4cHcLCrnJvPkmwcs11lD2Vx1nZTSfy
vq+5VSTK06PBaVOZjcyyUbBSLwgcAHPCZJ8cDhBs8taO8o7UY1HMn9BkVPPutenh
FTc89CvUOpWbmDVQiuIYGXbrOZx/EhhoNQQZx4tMuWPYqdRVt6XWhxSQU5+sk2RA
TXgcEvqX9rf30XB3cwcCqVKrjLwABs8azu6fQRGHxduDbza79vxWuMQJ+QxAqBBl
nlwyCU/ggf2mn8MXJNgBWd0a4E4qHT3bW2wlWdq9ezosJXF0H/EFkXIzW4DnVgQz
sm767KI6htUFFWsPJ4gJ94c2ZmKLl7Og30l6PDRd3YwOegxz7/ecUcdaoTO0M5Mo
PULEpLFBr61IiHUAh3AMs24084CvyBIX5BqScN04jtNMAbQ5NdMAGm41MblCwWcn
i5/Tcm0g6YVRFFekueGDKBxC8ss8xZ99ooyfnS2IlFysHVqg3lG1qDP+chPl/KVS
1vMNg2kyBsA9VS8bYUeJn78qAPZNjGdqdQo340WnjG5lM1MQikBo2vWiZrS/4tDJ
/bxnghB8/DGhC4S/+pJdDXGKGppW3SLesTm1UzEud4fVHjw9UoCMwTT1YePricIi
vIgrUujzjOWF+wGMiI0cVdARO2UU48gPh4fyvQQV6zMStYl8nP2RUY5YAhiZCXJc
EcrhCbWxYU37UVtQtEInWPHgdsXp159kETe4dYDDzdq7/X0DSf658/rYnVgsvuDR
To3deQkwmIRREGIgCro65C6vuoyiAh8KIsdkCKJT1i48dUBp7pTQLM22JF9TivsZ
N2amKHZjCWNk4XMM0miLLeaKbL7E8Zgumx7ryNKP6PULRDNa+u26iKuE7X88rkC0
zb0SNmZ9/ZA771uCmlncErRgj3EW1Ryq4oAQzFdJpUHJXs1shZJqgMpgnLYSf5DC
RxQ/uLIbUkBOQR6KBZmzY+T4pGiSfH/WD5RqU2+fUHtTALCNcjUT/TjDS2I5Lgk0
W5cSSNYNO/QVk4G9SxC6J5ojUFRWwP8EBHvdMmibG3O19dHvqZG9fKHYj6auAoI+
rHJpYpXL7qPUZN3lPe2bfSz9Ys3dRWK6IaNmBgoNYQO9RBdnESnEeJWt3zAii2zS
5ZuyN/vAxAL8qIrNnxYM80nu9Ew8Aja3esJ9JoQfnvRvY6FDAClsQv1bgxkE+FdF
gZVMGb5ETB8sSMI3ZjpoLaoWUY/cK0s4QndXOKuWrzacFaeLmjgIQSGSBDX1bWzd
+X+qPH/mIM7zZTRw6nPw6spIdi3NFHhMAR95TgWAzeJ143aguuzxB4R/wOnYRgyo
OmwOHf8p8gz5DFWB4kf0PBJegFGmOYWcWPS4hHR/l/wwm8sXUJS0PkbaFyTzD025
Jok5ICvIblB5kKIOJiBiuQocU2utRQX7SLpxXcfSbGncDr/WcQrBOe1uDsEBNKb6
6vOtOWAZlJeadPTDS1Y6mxWgGZtn6kdaI8walrfLAHsuymv+a2pYkr0iYgcH95GS
ugndMutWDyzumgqLbJp06glGQbrgqBUFAt/sk+29VZpEhSdJE0S50yLzpZOvLECT
05OzMSgiWvUdYjTUiAW1nHs/iuFqcVa2h3guaobgCzH5yrlOg5amXpcLpq7XuWok
2wzMs1f5xFP7AjyYBXv8e+gCPCgcsDSVa16F+8uD4m1f0dos57Bn5fT8QY7PWGbl
JZ6d4qxDAdGjbtE1YFpEL2m8zek/Ta4eQRpMJ+V9HyrTCVn6c0uBfjgh9GpQ3GCu
Kib+QQsvqNDRFa+os5GHFIP4dRznhMg9z7Xiej8JOBwn71P5v08fR40yVVcyEpwj
ZIgfmOjKXCfPb7V0IXq4DLt0nzyH43jr0YpXles1UWu4iCVqGIlJFngf1PwQAMSU
hUOHazpQIVUgApu67PvUM5Jepnoih9XjkiuklPJcR/VHrs/PSDr2EhG8P1y21Sbk
klUB27MJlqENket9Pp1yn1Ebr/P/kFXkmTNgrSVnNwcFQUgmPnbEhicMQkHaLsrV
JIc1BakAhkAQa+G60yWeInosVN/D7qEqAHCsw2UHHF0JU63uISQLziDRcteIVvRk
KMJfeyZQzz/U8y+oIApwOxpGKyTD2Kgr2MeuqQNKo9WqbrnW4OiU4LKPwJhtYG/r
/irKjv4IFJwd1to2eCX+EKTIJ6MOrRd1XwxSE9GWlcoqTWVSaXZYvdjFB9z+/sG2
2KKLjvZFrve9G9lPs8Upzq2DAzNH/ONEDIwGp/bRnxiVoiLldBNhxYzbEvUd1Ouq
DIdJV0L+kTyF3XDigqD9tQm+qXQrvSWJxeJANr8ws3mNoFPTvrovHcDlIjTTad6t
B5Vga1qm9HDekqqRQIzyRer202qngrR3PiS9wxa0GjDzlbc9/GPkJ1j/zqHKKadI
KHu2E3aGTT0uepHZZezhv8amFHiEqUvyfnQWnW/CWRUtukCImxS79GHnflGwt0eG
BaZcUeRceDQ7Z7IyXFte9vFk/2RY/4dXvhS/mXtLSqFS/J/ldl6NnnZRywkRBZOa
DnXAJj64b5lsB4oHiHSICv6rm9WdK0uSoVFi+xznx48F/OzBeKOd+y/3TA3GVrWO
ShV8wwsthTDNhAj07jQpIrVb/Hz8mPkwpdjHQ13SwYytw44So6b0+Ulr4fzwd4pE
hdXUK+Vng0d+ynxuIEEOgPIbAqg8Moh9mjdfqlpbWtePiIv9xibW3fRebQ55ge84
090htMZctZsMOxlGTZcvwiQ5DjaavRkoJSIk3wtx8ZDRdRoniWu/PLEO9a5BfOVo
1T4C8P2Lf7LTC4nBwjOR0ZG1jNYa8J2ZWp3gxee+sAP7OLR8IpF/LQqRqw+Fe5cQ
9FUWqU3yWwjizdShbw8S0LTTA7xGRYsmYNN5NdSlXQr9U0YqMDn7VP1gl1WCO8Zc
/v/O3ASaGYHt6GI7qmB/BulQNqKyZA1yKgfYwO3lrqTScc1rDCf5F93TY2AVw0YQ
LdKttSq2W4zwFi58kp/eAom68a2GnUulCjJYeBqigOIdF0TDMkafsbv9YoWEQijw
nBeAaAZtOp6QqCjbcTjLeVnR7NHo1YrvJllcT2WoTg8+u+ctbl5TQtssb4Wa9L/C
XFKtQxPSnXJltz6uqWnGlDfyRhdXPmxOoplf5Ms3tvS6j6DhI6enLCn1nVRfzceC
1T2z/26Sjq1yasOkyy8CwJ3h5czHUuNtzwdVL1cAwV+IlMGJ1JiIHwiX6ADlVm5X
bKxPAAi86aWPCevnKBZhOIFvb4X/CaXj5Uky8F/phR/Kd9+w4zZWzn8Hbodw8En2
T3fNxNacjMLdV7TyNJ/3MA2y/nKQTv4P+s4d0Aoc/DDraJb+RwDevk79fQZYiKg+
wScKAfdS6lKASZxFy5Hlzz8lNlA2tZHq2cQfmBXB8/BBo1qZ/FN1qbeM1P3HSjXa
jJF51mlNii+khhg7MGis92Yxlut7sMuPfneF25aWllEr+lIykZrpZC1FU+RMTBJG
n3Ecf/H4wYJQxwWCPLEp0ye6xJtrwcyJYMXAwOhpc+0pM9piSihmRPov/ALBlESs
DSSrbxKLIzH/4+ZOSI0h5PSLHpZw8Jjv4fD2+1B+PJQtcLyBQj+7UT57W0jHgVLw
coFBQtqINJxBn6rRrshqsJ7s4mTo/6MTw5D3ravpO7uYtusv/YlRc/uVt8Y4wxTF
ojtd0BHqZB0iAjTa7R0to5q6eIMr5MS0/zLjibiVQz/G/VgD7w0zonizOIuXYd6s
pYIaA+liFxPPV21AFArxM2MzQTUuNZ0f1gbQ/7xsyICKVM2nRyRYVH15+rv25Azp
LZk7f/qq4veuFxtUxaLAmPdRAqboWFLW44FrAL65Y0b2dLSTslCMBjFrvPGNbJ7j
kyAqbZKveJTT6dCDFwoYDh9CPhmj71iKMOc0MxaBAxTxBv0ddDeaUVRvtSswgle4
ou+fUzUukc7ut1htazY1si1R6Hi3+x5D6JQooCXSgN6Y175lanJ4Syk6/dn04RWq
AeDrExwlA+2QlCVr3/NZg4yv6Z0ZKJya4dgI6yAd7jWMAMeTioW9KJZ+Gp8IFPgT
97Y3icp9GXQ7vKtbxaosA2I6drlGmUzK+gWkW3DaDerDdomCVafsfA1SbqzPvFx2
iFD5aA3bPPsM+GeJjUAL8COXw27Us6itqpJGUETQPJ8BQ6bbBxF1vCgHiqwwQ/iN
ohOpBTfiAtczPSC2BinAifVRWavdAcHJpmvLOcZXSBaOf0k0And7dhuq06Zatdoe
pFsNKy2OvrRUPe2z8uPLKsavdb8wmxd4lEfJZY5DhifzBchi4TDu4CuL3ti/srnt
WOchJ/ADICDMatlYUx6cpSbkK7QzYVyNdEakqQBP7+XRGGa0eOM3ons/FjDWvmSy
sxqX0q5T+kjd18+ccBIZ7WdwsTZM2WdocSD7A1k0R7SiXJ/3z7mMWsR2M+wZ2Bbu
/nh2MGEl7UELzHkgXSIDNoUza0/yI6+VnJ19SWPx8kcLSuTGUeUbpd7tkWuGrrCD
oWWA+SS6truwYn+X6jRg19tg3fryXKXgQaBb7YNcxTsXM03e5dSg/E2Afr/lUkw7
Va8Uxmt5vwPZetwOTIixRoHmlrLqbfhCNLvI/1b8L1F8490mYeoqsBwSeeOOqSHB
FHZEvh8JrlC88Bna7FBryq9mK4TJXxB+1khRTX44azTmivRRqhNpFdaPM+5OSuZz
j326pwxEeVwQubMzYbCeYlyjZjdaV44JO3lejakZcAvVKhNOtRvkg9elDSpCeUHr
RvJggxLMiNqBDb+t80UGC2Uf+j+oHplr0qg4HNtuAdxqmGHq4TzDlvqK28Tx7f4A
oUX9OOqV79jF6wNHMVKYBjuuGtjqkhX8djJNrUXhusF+c2YfBAdT/NyOPAr2duJ/
cRZQ27Kmv/piky1u4YRy+6yOa5ymLZCXnC4afUngWf8S3rybdug0LyuAx4qmKjop
OGX7SxCoKBVLc+pHw7vGDxkw2bqkos+jLk5WBMUDEMOoTUZrWOFuLiKjLc1EGx/1
2LHtRQl98QOBcHjUdAtRbdLIfH8GuZEmjKjdf6+94dv/rOxIgf5ZSlnrgov4p0d7
njoPY1Ekyj+bvHu7CEdPXKsuRQW15vvxjIwjyjJrOYquumo2nOVXMzK4zQLWlHPo
SRAZvOLAQFyMfYX3geRZQMNwnvjAZZRwpancbXMBBHv0hTkzPF4eOAFvMdgpIWXi
/BxXnkOQa6Msg96Y7azq5sQb+FWO4pYeN+CqeiV+6d2C9lfNRJo9dF914BQhOh+i
dj30dQiH+juxGFe+yn5DfLw4P+YggrUQojuZmF4mKh1MF8OnwOKkqOm3m2zMXTo1
euVTvJXRVcG5yeuvjMXN3QZs1hhS8PNFpXV0ho0MJJhzi+d4/JyzYd3aYFlZvkQ2
a2wXCRuQk0baps/d5oes39TcRhx3q00yGgbEkDKVdfywqFC3qHFhxshhHeIgQ3Ln
3S4smRDsm4pHyK9G0oZq9na+NwdLsw9yEs4AVPdT7KSgzSrq0zAEs3fWzFWA7uqv
9O9pXS4GLBVoZ8q3xWYWFwPzwwWiEDyyx5Dtj8lgbq0VxFrjxdnBYrUGml/irOf5
MQg+K9MKbU5aRepT5UkZ22wnIoPG145ifLkxqUenppJwrEwvLk+KaHbyFTuxbmg2
x8wfPPMltRH+W62bJfF93A8mrD5fJHQFsAf456zaIiqXNCNNuMGDfjKiutHoyWd7
t+e2bJiGMuqBhnn3qy0NA/DMmi4N91mNtdd9SWUKOdYh74np0HIMTov1qw22oCCI
1OePv/7XcNrFwOoYd1e0bvDoHeBdK2+3l/yUZwoz80z3h4W7pZgxg8SBeyyRGE83
uXnJeEusa7hXNdvbAf8ezph/TtpBAuR27eFtx/W8g0igJYJrSCojNi9LpAjfadkD
MLrGVoUntEB8A1v8RlAGTzX9Nly8PsuxOT2pWu+KcjdIfN8Z0uV6zDbkPyeG3BR7
TcBNKn7dV7HVMTVXtyTHKf+V+j8TNC+t6s+4R4iFbfKv4NrKDrvMTYhllaTKId/C
aKZ39+rmXw7ukafa1wS6rWKYyxY9nl+kGF+It8TTGs7gEM5LwChe6J2cXdrmei8t
hf4lmaNWGieuTv9UbYWCodlY1EHu2n4fuj+v4c7cx0IOxHC0i5Os5fKsttBgUxav
wSiYtS8DBuWIgvwmd5PLFxcFpjuklCOLvGkXximmmNLL5kFeetFf7U+ocpJ4o1QW
trFs77cFMfFsRMg1isf6GyDRHv3O1g2pedmSp8KbdewPz+kQbBGMn/Zm2mlt7GQA
8lFnwi1pmzLyR+h6TreMptutSgxlGbuIjRKD6d++7gC8XoXGojG9H7hhCqQNrNdG
NGKKApIaizLJ28B1KlnSy8P3jhktjoRWu8REa0reh6NFXeN6eLgHm+Hms8wyiqkm
4vKRuXTb9XvCWVxyedjL+IurrEx2x/1P99axp+8PabshPaX92F1EV+YH3+Bq1tvZ
ZhwcD+6IwHGFAThTacxkl2YU1HqRbwlTig80LxJkp+17VyWb7CXOTFlgff5mEc/y
0qPcZAA9mmGhfh0HKspCercBPZOrBbRMErIuTdIZeDHGeDIkO3J7c0mpmz8xQXJm
nAm54d99wDszHAtM9IjlyuxYbRucj+n1kMSjthI+vcLzsYbUYLOSRRUNiOAQtg89
F6Kxf5dJ+ynWAuXvBb8jeQZZ+zeQQnUPOAhLGcTNTP8PWE3R1V6+HdziThALz/tf
fESgKsA+yCvFtc+Mf/2FjPJF8l7RarHl+hKz5KoanKFZAqBZ8m514FsiPdCl/3fa
qy3RK6ld30qDT7dsK/NkQ4g3/G5uoRC7mO0OZbTe2L/uJUmdjL1BjWEuZhJZ6evO
FCS/plyVCiBwLa2VBJBlY2YIRT1UZfNI0RdGsWJO6d2ndYRekwsC2PSWNrl5xEJb
+R+XvCyKHYK9A5yo2ebNb2gVzaZhKjmVOV0uR8t9MwIg4na6INJiwy9QzQqKGGnM
doxDtRl2/pgGptTX7wm/tksnCpGpcyBds7golzeLEGun0awwgMmsq2Xs3P7siOoZ
TA49STvk33yko0K3tly7eESLRczafhH7bND447woTkFJFCbKOiukyteMU27imGG6
bgZ2n66DoNe5XvjVaoxcSWy6ClHFhQ+08RG1oE41mN5tic+wKsuRUHf2I8a6XnJh
AHqVGyHOs+AgtcdiSG5TSNadQbk4t35zU7J2aZWpUAMCsw4MFVXvErP3zO4jwrwh
eaMRmwjZFst0FrGnmymBKTlW/bOs/ZZhpNsRmBioykY9Ps7neTekJtAj4iQPjjbW
t6Bb7gWV5DqHD8sA9PhnsVZnnnPWpdHEHpDiQhH1XK1ABH4hsqO/EKuijxCRT+Oe
v/YpuDjQ8JRnbcsCbaIrjmX2jhXvC4qiutN2w5nwjEUvEGB6/uSne+qT0+WrH+nD
ICdmmEk34piObYaiX2YUnp4zcndX6W81Hu04q4iGAlUzYB1zZbnJknpi3TI906N2
Yp9s1CN5opXd1Wh2MJG0NPAJmgzbn/NnUkGFm1d2/XWgdbEd8o99UG1UkZsSQ7MS
zZtc8XqDwTrN+0y9NF7N3mD4q3rIaqY8qoDHkgH95FNTPK0sCJ/GjMp/rhuY4vJ5
SL/ROBw98R1jUNjJ0p3OJIshRZOHDgdgHl9mkV62q2mdgQyTK1l5JqmB8Iu6OCZ4
irtxC38s3V7D8pWtkGlla60SuWFqDzBw+u+h3ZbYTXiOmiS2bL4Sbb5OcaL8ICvB
jtbFInlf4c5ubVeA094gqSmCt0rmXKuwPkk4yQK9taXeAESHAJnFY4kO9LnXuF6z
+T3rkFWyOniSanozY55Fc/J9jm9WELLJlgsgVZgaqpzG2gTR4LSP9biNdDOph9/P
gi0Yepp5Ti1T1M60iauKyWq9nJpMPAcWy5YtuWvAZCLHOHsTNVNVGkhHEk0yO9VK
rcjiC5/eyO1QBz2fSiSf69k5pD4EzNMiJ4WuPLNSvanqP4sjjLUj4UAJf1XZ1uc0
I3WRId1Pgkjkr30p46gpQ0hxTklHtYGJZEy0Ge69FNtvgHlIbRyUXCCR+JJUciZN
d/HSSCB1SiTiwBRjtZcNUnxNRaUr9ic1koiMM2olZlBcOn/c+3dfZ0GiZZLnM7/E
JqUiU867MMk5fyp0XfBeG89YMxe4mD5GUm06y0GqqBG+u8Tkw5nh22gBuG5cyoHO
LQ4BmeJW+9A4iV+8fQ9FJj4LcdRvmK3mgOYI6Nlc4UBsjp5DL43mJRbPLwCfrUDT
AmJAhM93ed7iQW0uD1Ta9wBG3nUW8OgFV7Lhv2DWprkujRmhgwXq2OifvJfXImVI
4bcLrILCYZgnAOuzsu09COvXJepZjwRCMx6jonUeBYU+IebXdPhs9DrM2jtdpCPH
eiWUhmeGKpof4EFFblUTGkFnJ42sfVGKM//uPO9677GGlPVvzoPJ5pB5SaOj6oi9
/hWyqdUgoTDBCq8QX6L+tOvu85XzqCSwKyIWGI4cALH3hJT5jbianJLpuTmb7v1D
FHD6h3zZr7rcXN51+ZUPxxZxu8jb0XQTSr+7fCVp2OgJBUcbMF7soYGN7ezyQOTy
PdwG79HYz1s0OSPhhOns/WtI0W7u0y5eflXbpp1ymIOVi0PPb9uaaxZ6FFCT5aJI
3Bo4/Fzud85MEKGFydLCng2+hjllMmghH3DQ6oLWaMQwKfwQAb4WzFsXYzX4TjxL
l8fZcbtrN2g6tJJePgdMZXpTzuj6fIp1UoKa4j09g/D0h5If41yhPXmk/dbV18ND
eMpBt0OSlX6fRfaM8hz6vL9/tAvHB5AJI07BQG/hBrb59tVvLDPsXBCqsoQTRWzG
vowHKlAbSTSnub71KIS85iXC1kb8vkzYbT9WlGFcUJnWS7++BFghbD8L50lST0hr
+2XR60JyMdV0E8hFGof66v+Nkt+fvATsF5Nn9wdptig3NkfN1LUGKbqOHv1EuiwP
jCLWomJv5CuskBv2dsKX5rr5USVYUgnKugkCfzOGtpB2WIB5d3CV7PIldFJHfgN0
+3qKi+5JsPPLzAZ8RI6RbGvcPS53EgFSXOA3wHhAquyaRTbajVaTG/nq7SAi6ifU
g9jdzmnp+TTLfJktLgp1kapJmF5EPOk0z3oiMm0HdzdKXyiW8NRtkzyWg18PZpLk
9pHpuIii/pFGYNFaKTd9voviMWFRvKeDsRkgX6aIiRBDegSjkArgRG7YI/p88Ejy
N/XHcMRx95CWIa/+NHaC176ZWHHSzOSoGS/BU+kdG/BYeDqD0AwhSelnIUdKijdP
q4Rj0kjr2GP5ui/kFvlLP7uUsGPq9tkOSLSB7r/h/MAfgEWChH2clFC/0NtH8VrT
oBrgReTGenylPVZ1K3ECI/iWST3SyjsPs6O0dVjBSLKrajRKMVowOcpQGHNcbfbr
dR7sLtlmj2mtpZLuQvkKGu+KIdWNNFy9iIfRpkD87K/IQvdG+1+g8CTZnY80sCbJ
j5ej9kTDybcEfNKhpJzpxkm9BM/4MRkFar5aExNed58VOG3Sy96HW36eUDU8eIo6
pdXbFGAgDG/CUc1kXa9J1bB3Tn9YuMG+nUovrrSUIwhVb9dCWKCU9O06+XBHtU/b
vDVFfXbk0roS95o/0JJyFLi3E2iEg3Tvim+oiYVy0U+dq73F62KqJ3OHAa1t1CL6
gsGpDe9pW3LoZiIhtIAunk6bacFFtJTTPCF8nEg6csfBq0MV5PhiWle6WvKsykiO
2zgvLEh5RVW59m19939gVvg8RnzmCeHinp2j75YMNC3/Ojn7i/cj3+I8Nt9e2Viu
kdXWo5tmfttxh3WYwNIU2FDJk3q0OKGUOvlY0RXIG2+7zl+D+w8LraQXVhFYjIoa
0+1bVb8T9aZoeyCHUfzse97MXpz91qB9BC7vrsYSdokiubkfQdQ1MTynyZ12Bal+
DY4KWPvSNEks6AghPdLNHmn1gZRPe2p55ccJsa8RG1KMFyztRWZPRwNRgznmYjb7
Zzsba9dLSPAfINCa0gRmxSIHoX93STIW1coQNVl07pOcrMGekI9qd30aZsADhLa7
DXZXPsW7voH8MdDRC123I7sUKGHIpSOdXhqGRnAHFuYT/69mz0XfTeesdJnPkhav
U7K+vVh4lLqTlz3zZx8ZylLWrYXmCj6wxS6p85wx76J1f9XUCm99XBATC+hOAleI
hFLWvrVzSki97YJdTofX/u0W8YBsz+VvYy35xxNeQexg+zhb8Q2GAftNsGM2WhQa
wbpDWDWA5+26XEJ5S8YnctRoD2bzMpsdPJawOXSO5ZTgWFdW+z34+AXZwApydi6G
m/npHlDYCteJTCrogBAfBCEwAlicPe/DE3esg8HxVIvOlB1bdK8UEs8qfd9JUOPw
V3+M5SPJ5zkOEco4weA5p3fIlPIOx1YvsWW5AgqPjvPmDlR4BPZBjUY7FtWZcaFb
VsRxeEXRmQVtAU/xnDOoki+cDItbTFazqoo88pFoUEFOIpQ2KtMbYMaMB72lZ/VM
VoQecwlmuwvKfL8A0HLHDUIUmVsr5n2joTJtX/6pX5/XlWL7ukIeQRWy6QDakDGu
8nUS0gHXoc27r5/Wahz/eFR14npcB+aQCmvHNrFGpY/8ihhfSmmA5jP6SXNAX3H+
VC079klEEEH7uxBCMSfEj8ODAYdn4z7HKkKVZCCnnA4pysXFyqUNZwf9x6SrtglE
CASC/0uVeMyrDlGUxDi42dM6uKcyamLlZsD9J2Bpfku4He95Hj2f0WmbksnZ7/jB
QvuuWQc/NcOI9m/A6Gm6TwAjlQDj7FTKfd4TU9pdu86nJO3cY6G7zsz/M3YUwW9p
yEvge2myy9i16YJxEWVSIqRKKz9jQpuJQkL9KXnsO3IijyStCiN2Ii27YUa+upm0
I0twhpqk1EtiWAav4yzljZuZozYASQj5MqfX9xjIFB6nLc3vtihtgl6840qHMy39
h9yh2ILH1wIAw4GWB3Zq8noUhjUJKQjd1loUYtsJxMamCaqdsrKVdIxOgzA8Khkh
TfUevH/Mxmxdeln39cmk6E4kKsVX3F7hvWqer9rBX54a1PpCGcyWZEIryXrGlb+0
fSCbT6YxehGMwTYFeXxxrZKXBQ0CEYCli1lCkNR6evGeufhnP2lgCe9sOcXe4z2T
XKJhIT8YhKQHxqkuxTUyZTjA6v3MM/CIKlcGO+dAAHp9NAzrUjDykydz2Nq/LFoQ
f/OojKTCW1MByr0xBK/R1FX3a+f1AV3Zai5D8XUAbiFav9xRSRSdzK7bfLS4nxgl
7fNgVVwbuZikr3xxVYCijNtevdahLrtxB3KmNsgejfQe5TXXN5+sSF/M9GqfJhsr
rnjUaPFVb+K5f8uFzXi60/kzusJwE0Dde6NXM10u4DcklL/RvNDB2oGd5bKY0Yzb
1WB4ygwklxSMHyGQ7g1yhSM2rkg3ktTP57JmMzI4DZhAZDEs6SZQXIAEvruBhDLL
OiA+IOXuowfGZrsmxfdqzzVA4epTcpGj1C8OYGG+xPr2+NRQkigI4WYY0oizrTZe
5krsl30xSmEqyaXBhLPavFcxvuawuCdwmhZ6v7uUoslhn/srYu9h7V3t9nehYbpF
2dYBATeMwqk+ErUmPkYTBdo688LC7vT2km5hso+jZbN7DYjYDmPUGJMiQFUfA0A9
mWh+F2wCucB2wT8vgk0ws7QNYPb8s2diJN3WU1b5Nmwpyohe8aXNFijaGihVPPTj
sPOISCaI3DmQzC3A55Hwd7orbCiZjijihNJnhkx5f8G8/xNp0rREtEQ11GFRNICX
DLtVPAoM6D8+uLkK20Oo6/KgwtMgU2lcEB4k2fSFX7CVQqg9k+DLTDte8Kt56mmu
fV6H5KXAKP+upWatLFftA0fGPg+dkQKN8tZ+inuMxTq2UKwnRvywe2QZCD0oVP9a
DUYSjTlXy7JAA9Qrpg4mHqJyGf3dy5ZeLzw+M/xjxDaCFGJ2oR+Vs8AVVx6l2N+s
Mgyqp2TX87PnjeFP8MHkzZTfIJEUantPV6XpjZNxmaaQpkPqttgrHUKkgis12xBv
TmqXdOYFN/daAXWvE74eyRud3ud80wxHYcaz7cB5a1gQzkfOTRlAxhAUPEZBAsRq
1tY7CujFY0hdiipBgX/Mbb5/BI3xcnWDOTDJEp5YywN6iZYgApBLo3UosKj0yD0V
51mLdaxX/LKjKu5t3Q8kaTzsiMEgE1uM6yOVWOitxW8rHS2l946dP/D+CdZxJRQL
67QXmy/wS+boTQS1LAD8BShL8Vx3I25MCjQUDrd1GzDe5DNkEcBTJ/pouY/YvGmU
5civZuYLCuehTYHfvogdCpLS/tDPDFi9owDgDQLNG1A+s28tnoSn4OSXgFVV5l6E
L4zYThNQC1MFiyWfobB+MX0QJcY+6jC8YwUs3o2Oubvx7XGZxK/G8mG7EwbthIA5
7CQIZ39rxVoSzFSnwd8TBXHlH0CyULSF/P3mwjobBCrat/b82TCQ9jcFRDFyFuLL
AOgogitS/eUk92H6MT6bpkhbbY4XT/HM++cGHEbK/JdVilK6P4XiACvV05B55gDa
r0PAtJP6srOjfypWGv7tJdT9YIfGzEqqS71v1HI96rbgGH86La23W5t3+3mRBhR9
qWWNq4yu2VUNjIlt8y7Kf3nrXvlkPFKXRvOzBBmdkrTu9RnQX8Ma7tUxaWCnP7fG
gl032dBwH5AM3pcVOaXFr1WD6dX64eK+jZ8Nk0yJFK/YWEyCCUMnfL2nYt5/8MGH
kXYOX03KmsfnoAqKRP8f7BrucOxr0IUXa4zEj5gZkMy5i4wHx9ePW5HmqUON+cyt
vnwGL8adE3XM55MVh8YSCxugMST9IqrsL5agId91lcNc1VfSV4JX+pRoa1Vj+bVQ
zbSbuoGOJfFKtQuor1eJFG8tRWHSwJ04RrzQY0JDiHliq0wX0WLjBI348Jyf5B3m
GVlZdpv7GlgohtB/0eeYaGNJDeG6/orh7ovQpQmOfKsZ/yMLk6kBdrUK2/m7okiP
7isvwaeXZkM9AwYTJTONb0DVuqeVPjKd09uHKnlkebjv8RbMqPcURyKO5gLplhvM
oprvAwM3TlIha2IcInHdTOpFhEDebrhZAJyPhLoJWQhCN8BYdkCG2Pdz9bRhyiXO
UsFciSR4RGl3UQCzqJGt9XHZdq+7FTQigRcFiz9vZ2HLClF/F/E0uzYZmShrWwdN
ZC65Zmjq9MAZsivYL9Lm2M3uKhl37T8KsP7rSUP1Y3IyZ1SytmMZDFUdZ4jh8wSJ
j4Ytt3TGh8cTYL+jV/kJIcyCg7g+hp8+/KZbtBNFeROsZ6ahcFqUL2ID5REsAUYj
7rD5yr1Lotr1ZUhFGoeguqwDiTPsDjQ+GXnq3X+uFjwhvnTXJ2iH86LbdH0ph3If
oSeTcTQosHYh/7mTCRUCVH+PY8FsYTuTgED2enw6POe7LkGrwjVIFfT28Y9+nbyV
pdT9VhDZBGYLtcoBxDmy/KAgvkHr7yUkSqaDlN8d8Zgv7kENGLbY5HTq+TKUo1eS
y8hOy5mYSUST2Brj7Mldt0+fckCm1xgui3RGE6c1EzK1ggxLyktJcFT/61CheCk8
rYOIgh1cpgFvJDvcuLVHBqWSqIEOW1hmiL4tSl+jwv56hE8shDm+gPTHJ6TxRqQG
8BjUJrVHqHZM+57DVU2J+H/PuhrvR7vJnTFR2fbC8fxPMiTfTrbx49vVl1g+uCtq
v3+klc1RZrEj/+q0Bnr+3s6+gOXM1gJfbognUKc7MUxrNbSmrLi3snPWe0G++MS4
Q4vRdj71g0IYoh3iXFd7afnR3nLkKrEWzAM/Z/NpfcF4VYtG8FOUeh3KCo3a776K
wVd4wG3OCKT5FrVN1FC+RzFs4yIK9dNegrZ5PbUPJQkYeSaBTXrlBqjEWB+yJRRR
zkVLd7xklZQBgCSC0TGuTwNrbTjWpPszVAAYANEtJJCmD8oIdEjsZTRtKT58RaJ0
tZmCkUK/m12sRucx3e9PHRW/nECf7mDAfofNdcR+y+jSdM0cOpcjpb+SsgAN+D9I
Nqwi5O7UIbEvpkaIyTvdLLfZsXX0kPD66ExtFs2lLY38yfMcyZjdBmKeCl2AZqLn
l4DEXEU1mka1OXYucwQ9OX1y6P7r3uAGLuTRYlKWwUC4qcYaJoMwt7y+7pieaW+r
CxmrieOzx12osmTCkj0UcRqWs75R4qsAZp2fCw/k72RLs/HY+f7Xv8I/24iFBe1W
xWgGj/U7sguL4mXzj9NjsKRt+Ace0zficZ4hFGXCTsqKc4CyT8e8TOSwGhNP+hWa
bqy/znUxDCke+BxXRuodx81oebR9drPX4TnDLiHK9WmFW5P+H6XvNhrnefCo4UIN
uXncf9xjdhbp872RZ+m3RXdWC53sIYHf5BsGcTst752d03teBAjc7M9P0t+Y96Ci
AcY+5+or5qxliPOXhbpvqaQMobnKtdpoInuTAjGXhw17w9UYcwlyHcgKfR/Wq7Jx
N0XV0yhTYQJ8w02St0ElNgIrQyswqkuPkDbxrPaZL08vlQ7+3gnu5GssHKm92AuT
kQafUDV4yEpJqq6Xn9okLtkwpD7qk1nNSKaNHzoGk6opL52Ul/9HQAHr4ass8Sh6
/EySx9ka0mht4i9NVYiicqhYixXwJ9sNB9dPFMdmvrk/TcP6iUGBuTN6SEzdTfRZ
xrYxgQx0/ndqGuZvJxL70UJBwWPgplbID3Jp2eXH8mnEZMVK8eNeqXzOUAB6o2fD
asWdIkeIXs+ftTrhtl0XPWWraTXD/mEsM39N1V1YQyTiPFGMKDUDpwq+rR7xwQXy
hCj5IEK9E4oF9R/bz9s1yQJS5bWp6dKFYAonPMtl2uThkZvwh84668SsImAZdbHG
V6I7ehSm7SStcBmTxk41+C3hclMalB+I5nEgicq2/PwKezn68Hyr/dVvaA0uxyu5
rZtEMnlE2xz+dpu7k+ImvDXhjxc9o01WJf4sTfWPYfsp/f8+K8SAuHVgPp30lDgJ
rVOagMpAVnmWX/+FEQzLaE2CYhCgHV4AfnjJMKXj1J8DKA/PFF/eywR8Mjs7Ha4c
aZNIaZTX6OFUMHN5RQww8PPrQj2G3tkUDb7BQ846LIHBnubKg6KJrh9ft9JGHRYY
TkM/cNWC63ue1hl5aNbt5R+/nkEcp+1Lsl92POfqDz1mLhiGuMgnKKuitkYFFsJJ
aWnEQOGBF0Zpq6OuThDSKDDHumC3W2TWLfBGj0Ah9yXb4yne7yuLnZSJJAUZIt5Y
4Lg3r0J0cVN557gdLKr5FaZzH9IV7wVX2Sdzp7ee/caF8jvGJbrISwbSDAvaM7Hr
VADwS47xhZFPPYcYjFJNLWBZobd1poco5qbbLz9eHTeGc1NrWReg06YwTMKuDHO2
a/Ch90QwzzD1kgggrmasKpm13j9ofbgf+1LR2pFtt09pctwWbzvaTv1DpmYZTNxH
9ncj4+M/iaSF5RxIF/hiMsXPSksKw2r3oi824tTw4Dz8u1OuYdE6AHliYg7+l/6o
fsUvmAaTBlZhmOrHsf6I0dvMcmeB7RfhX7RImLNUqYOFV+PLAbOUWDCpEknuUanR
W6nIf7vYAJA4KBSyV48Q6hZyDenGJNwZb0W0pFiopbDTHjY6J7kV91TGGdNOe9xC
M6dwuNiwJhSpEySLdyclhs3wko5LLYb0Jsl73CAifT+65oL4ySor0meLbBJ/cZoO
1xfYem9Bjxh6JRBLIndnXGfsrWGOlYc3hzl/HdvNYneAsPH5BBunNgmGGRL6X8vA
aO8mMqMlGzNcXyy/A6AqgKfdzxXnz5ISNc0zP4wk/FtwlMnDOJ06b0rfEGXHzog7
NRVTGVsEmQdbBIs1rdR4bLc3m4stFWcHchp5Gcr1cE6DIyOU+YmtoQw3cz0/Ly19
v6NWEHow+DNbe3cM+RlEAA5QKooOlt0bKBXJ0Ndfm7ailcEMbxCv6ad1br44XRet
213pMze6GbaclMO3Ngwdq9USmLJQXRMXSS0efcueP/a4lSYKlvUC+tBQ6W4bDG24
CUQ7HMYQqY+Fit7JJ8Y8C3tT7UUiSqzQnsAf9oKqNfAlSJ8lwH9wB8u25zPzHJ09
33nUi2L25hiI+xfUVUA78kWUYvitydG+Sz0Q75OjPXdKrxU9qmWQqG8lN0PRC8LR
nNcb8XB1XtXxRmFFcQMccv9iuDZzcFRIbGJEqNftTMSzbYuuDidIpA43kZTU6V7e
L6TOsv58s0yeWBDT+M6GKccOJDH49dCr7JZxangpCqhcZGAYFgpQsvknrJ9QdVlC
To+BvRmLJrLRk7ngqtg9VYXQ8dhdxfVq7+iLX0T4HxFX3h3vQBq8+gD9Rom08guY
VNwFIEAYLuzye94KzTnPI5NcgDe0OX80+WTRhK/QesT5DaXVFXWiva66bUiFQsly
ZT4Mz9VEnj5qXgecudnCahflPdNBXQLwzWwChdLMklQu/mHJmhc0vJPOtgBxNcAG
6/XKcEwiXDB6gTjQeuezSwhXk24sTNknLukIR7UBUuZrJ8YkOwLNQ+ugx/dSoeV+
YgUs0HBRy10FAhMTSv1UiHe7OLsOFeqpnHVqHH0CRvQ2JdMCc1fcEOEt3HKpzAGm
bep6MCZzffLM2ShEeehibN33dcf5d6skR8il38HEmrBHzOha1WSfG4DpHhkr9Qv5
QxYMQcLoc5FBQbZXt8eOMaLQ31Qre6KA3cJKj7vvO+qhIsnWMkYCRrDMiJMlaxek
ygH6vW7RVoAjTia5pyoxIfl5msf1iMPV2/7cjMeo9RPH8GxwFqdeW4wZNr8R3Fpa
K7jJ7PRHOe6ODHyg/YMQHYSYMOlthvaamU+p9d8cmTrD6bwSEnohcpj/1p+EHYma
nc2XBmt2OESqKCUfTW1cNaKEHyhNiD7iajWe/ohzzVoG29mLROshmPM6BwqzklMI
u9UgG+AmoqUDO07YuSUIKqY/+HbpKlMcKEQgyv6tVq4b52jEKwJj2XOTtSWUcpfz
aL9rkKG6ebQWzSOEhUtULonzlEWQZOQ3qh7d1++1peIz+5LM6ra8Khio8wIUyH43
J7cRpT4I6B+yXAfipObYi591MlIJMXuJbrEi1U6e6tHZfgCe6+5RZCL1DlhMifXp
lZvoVgabeBCOrG8++Mq20TmAh152c/PAar054+owahK7/e8IFWzxaE5JLob6RhWo
3OCV2ua/UX+KbE1YHbvW74kLS1u9orJmEbQyi1CNcEL20AwIcTp9wK/keOdizm2J
v4aExy3X734cVX+vSde4R2Hk8wHBbpfkJvI1djnydWGDad2CC3Cb2yaC2L9oULSd
t3IP622cqm9kBWMXi0vPyGyhkXzK6Y1kCuVGI+Mwq6mB7qzeIFcr/zIdxoLGhXtr
336jEeSE18dkrMnH2etxcUcs12jMqGISIoRgJ3q1gM6n+agI3ymoQfmo3w7MBRzb
vJHHmEqiva2/MYGmXWWFxOEAv3SiDxfp9hU2T1luX/hHgIBRJz8OGBPXow7qfSs7
upCO5uvPCyBxeNco5ytDkMJC0KFgLYWMEbjBhBL8Zs1gqEI7djKhr6iZ2M447Xvo
KhcE3C4gFcKD+JkpeE9v+6twa+HhWCxLocvGAQDVf++8KFwmS0AF6vsoSJxJivQV
vtXuBSgfYilQHjHTpqAyKazNHIuDV46qu3u39WPKEYETkRquH4BeF5Z4pQM/fsko
wQGnr/Pl/r7kFIe16e0+QLIbo2qtm6GJ6eaf/aet3G/Y+UsSmafg4OJ1BcJPpwpf
ZIR3vsubrqJqS3BE2XbdZE7KpoDiEND30doxjkZYRH0Rp3Y00UxIfY3PxJ7Bzd4A
YFc6U+HT94LDBvlS9b/ODIJ0zNYvTfPVlxyf3rvyX27+lXe7l06YoNgpt5r+SxFK
/vdKV2SfNjFxa1bLXAqxNAlQfxY2rHsPyw2CesV1oql/tvznAoaOSED/oFlgIGfN
UxV9wZhIZTC8lW7q6pPpXAJmta2YeeHpV1SmVKtFPA2wk6smDIkMJs4ZQFK8iE1h
V9d3eR1p7Bp22Cgrz+MLW5tbMuYajH5y0wV0Q/T/Inez75zlAysvavfga+HjUwOx
1tFtZ8V/hfAS5Smk7LSlu3uFRuI37V0tuWqb4ZR0I9hT4i5Wj0POYNKu6eIgCxef
F3k6QugN6F1OuyPn/dxO+A77GiJSIAkT1/vhIVB8XxcOYcj5Mq/0D3Gdyl4jpK5u
K+zKT2bo26xxeEF1xNzWMpOdg7a1WDW0uCJySedlqxBkXMDACfWUIuM5nMIAjbn0
TIZiYZB6JkDTfvIy2zFwI3ujAc+gFXDrZhKSgmot4I9xL/hf45vPahi3bo4MUoUv
cUpWSiFyVOE2jqg0/Nb4spZSGQo0UtabDYiamYVdZHC2chVdwsG+4bSts6SYtjiX
KInC+GYbvIDuCZtWtHlO9+qnqob5bZuMTNIvYJuVl9CMGphZJPLirHAt4eyWzkXv
wOOI4+mMHxJ71OndB54yH07nCm8zCvio9lMKk2Knve57MAbFjWGTV9Gtt6QrgCi7
BwcFL3+c2N5lnXrSRiBsrQopX+PYK0+lOEwVejo9Cot8pmE6mCkwcdcZacjEx4cg
SVUauZtyQ7QHfP6YVCW0BpZm2B30JeRlsSxelOoA5xY3lSGJQUKgjivEAKr0ZrQW
pj0Ic/6Wl5IpbisfGmXQ83yuXJuJe90zpVC253/29+bU3hgFGOsgZj9x5M2UtJtw
03o2DG+xFjyNPjiZeDQUr77MuqFHgajzw4livScnpzud7Guw5WIfA7uSLekiZKQq
aZienJxNMWRxCw1rSE9kqYMuJVNEC2HDiiZ+f9LqAvFf+237Tbr/YZJvHy4KP2r8
ICDmUP5Hh8dGiv+0mUnm5VeVN5pAZPzWDnZ19Ufi6BNFKLz7oC6EoD3ULBqaheLx
+IIyLTmCPmfBG0FS04MgzRc4Iu1UzGIFyq6jyLDFY67Ovy2MJVDBsgU9lYbK2NlY
bcGY6FZvlsp3tOl0MgBV+ycwO919oEJydEeJP/T76uIaF60Tk/X6RjDzW0av9Yvm
wYsgP8eGDKjd3Bu0tgDebs0GSPTLyeL3c4nvDd3yyjPjHeHcxW6FI4V1+PD+vBLS
k42Zn5JK9kzAe6nToCd3coCOw6zxqQfUCx5375XNUjPpR/zMIpHXtcXRWklLa8Ob
zlcuilKgs7dbxFIPD9xfZOjaa+cyHy3QAjBdiVZqJgCEIA4IuvfjJX9yParCasiG
xvN7524YCc7rIgZ/QaUU62ccTHtDg4Ky6XL2dUBeuh2VeR0fm8iLryqTRoNofYSU
BRbWM+D5z70Vo2f0aQpJrC/LFCaRPNk3glv7H+9urzG/QNdp60hVO/1p3lKuIX45
TwOZ4U4u1sMsNN+o3zg/Mwd0+U9aDaSysYGGxjzuWKwMvFa4Yt8SnP6bDtSCMHUK
1EAxjqaW6VeTcZhwTKnik6V8zddyDbpuPWdS6qh0ZIT0/Il9nOFZawHysWAtXaz6
Miild9bHkr+akvKBYFezMQxyOxST32Nvm2HgWZ7gvJJYacWVhWt82ymEkQOMDwz2
6h0aJ3ZOXiPUyZFgBkwdDGxx9jwnPh/4qDwS+8tyT0ftAZUkgbECDsHcaTfBkKMC
D56YGmVoVCGpLhKHsrF9HsescxANwt3Hi0E38Tp0O0QQCh99Xyt8ha+QN8qSbbft
m3+U+mOUahJJF9L5tui2pOPNYcphUDqcLvhcIo/dQ3/HRsCSMBXbb8UoUndPyKXP
85pp2czWaapMgEt5c2UAaRGY3+nHtBb2xbDH9/X7gFjFHNORKB92jUd5JhYrnKDh
i18Nj8uV64AiCD2p8zHbOWtfpeclT6Qe4O5R+LH66o3nxC7hRAoQdPeQlI4B51Uw
uwzKGKGf+54SltuNMmsWvawMAXHBuT+GnMrjGfJgsnM2OAJV822DBiUrW/JPsDLg
AIOL0ZlEW9slThvbcRjDyWilrvVa4N+fJanMwW/YzFUNMpB6RbFelYvYzB778V7j
VwQIE/8FE4HEse7V33x6dDBJcXZl5Q4By/b6etTonidxwEUEulJQbdWqVJdnYK2l
qaMKtoA5UYY71uN6s8IlUMcn8LfnP6Xtms0a3Mk2sfQun3KzO9TACC6F1zy6IZlo
EWQWaw+zpZ+rX6DHfrkfY6q5YYjcrN1MjPEf1Zwjcir+g9D4ydr2m9cPvrXxnCkh
/Uoc3OoirfBjaZg6Kb0TY2dVu/2dfbvAuyjBk6pJaTsQCSjk5Ot3HgeA2lYYGFTe
OFuWf1TasCzIOMkskMYv6qaiDni+WBVUt5YLxbjyFq4/kYZxtnx97H5ltJRJzmUi
l22VtdGpdYcx6owdJmGALXB8ViSMsAZgYqga7JyjmlkhaLmvOR0XAU5MV102JpnQ
FAsPUHK66bBuPqyS5XN6ZZuTrBJJl7ulfF8ZvTEYrB+oBOxiErVB7lhxXUIq1abf
L8ch+nU3H8pWWiYWZPLHJtScqrj8Z0IHk+nuUe2o0+hqSKhJeDMf0oXK620JOS8M
v6hX3uOnWuRijMW82p3w4+jqzO1KJdzXu3JOsOAsq5gIW3eKDMkFEBONQlpML8va
IivFewtcHl0rm1AdiqvFWB0mNwWi1slswYabAuHXkuSR+EYLhnLxbG+Syh79j8nG
QNp8jNtmHnDlVsfRr5G85wsfRCPT3+kNiuW3mZhZJOUtLO37EVkgrYuo4rHMXjaE
Tepzy9WjpAMSxoaPnW5idhAiJHQcEoMDCRjlEeBAViXAlg0yoG/sqKlnagmhKaWE
QR9m468+BahW0vt1I3ia+hVy7iDNKSlE7Bc3uxt4R3NiCih/izRuqjoKjcEfUowV
GlquSnv/SbxfoQ/F/ks1xymI6viF1yyYrBDX9rS/6f2qj482rmUZ06vLaS4ehRL5
L6cywDM5UP93Pah0FQwjtqM4HdDd5KRj89r/yZbBHMvXuKT5qtzt87YWDeyBWEIP
46AxM5M1e3VHjJPFX4LMNBHJhmYCJrM7zmoQr4o72g23Jkzsl1ur3uZzIN+y/mMH
O7J4cSJcf5O37XsvnUAqOvbuRZ2Xjz6ZD1Ni72PDbRY37NAykML4Hrmc3Ybre10o
ATEcd1oJIm65RcDrpB2y0KUXUUAqHrIrqDqbmcHmBOA3Hwr+o3rQyjDI2RXzJBW6
8zHBKrXQeZw+/mk1OYVSvmaZGb2F6PpQ+1zSBRLte3BOmtmUGdBV4u5SJpA1mPeW
pRPlxJ1xBDDatYM8hr5Wyxr45Ymo5k5jzwA3KSqKiioQLfgL20jcAq8wgjark/NO
l47qYZ1V/uQcdXfsX9vXgK+41OM6spl8KuCkzw9B2XJhJCYtgV61zBkGFqwQWGxi
Xj583C6eaaKP2CCsySV6aOJQjDz1vg0RlSwE2cLesYaj/7+i49xy8E5dkOnwsjBI
Z3+pI1rqchVpbXQFU/W8WFOfGbSz+b//eGy10IfHFbjyh48TbjidHmakyOkGBIbL
EoZNCsQRX8dlxQLBrtyZvP4V9vLm4vV7RRIyIfinkrGJZjVN9aUC4RCG4ac3y8Re
OsVFkN86QFA2rcFhe+bWnMS6YvZJfjdtHGfsEgohI/p7A1GRSps9sZYVZAEbeH6H
asCDxJcZpfhl4uXTuUIh2r44fq9GGcXFSWeOokcIo5LHgo/9zJO9uHuKpoe2OlOJ
PLuV1ofjsuyq+XnsShPe8z3vXtbmjCFU+jZcAZDdksUDIskZz9L8nC2R+fHgB2ig
0fZqdAvxaceo/PMJPMaAg6yZut1VEtv8zNur0+Xncwh8dyTbm0pw4w2T26N9DVgP
FIafT2GJPbicHvul+Wq0//8Rwe7YzP/2ILmgvCeP6WXv73hLUVMCH5BRn6XabpbB
Z0GEv9sJN1mIekOVvfSzwEhjvg5REU2Jh4DWqC0XZsMCBHnYzwHhAQAvLMTzHSVG
TvVzi8MaJ24ZXo49zfRH55Xgw3FIkBFXzLKjXzhVd8nVquIYs6jCElTs7jvr34L9
+sGG2bzbT6R74cBksTKr9xHygRC3EL7t1eGCw14DAH72vxfMW3++ETwV2lRPyuNj
S6eTm9DWCJEQJyUh2wXeohXjhLoTfog5SwfolVyz/kIZ6lT/n4Y0vYTV3jiOqM3L
RKyU/Wt3tqYfJJfCXfZmvCMDPhR/XQAFnQ8ct9Pwd7QvEvSSlmjen/Py7is7tGsz
HhYOvqY5HDbbiozIE25UHJ9VZa0CWXN4PuJgpWO/3bEvVjwggbhov2VYm0AwqT1C
rLj5OK/+F4yPL0VnNAPHJRMvj2dan2+n7J2EJ9waefMK389oRUqwKBU4QODD7xgv
XyLnWUW8HwFFhQtNfK1q6doe7V3rSHAca7erpQ1tiLXhwD2KcB12EMnefKeTS26P
bU1J6tG52eNExbE0iku3Xd0SfZ6pW5nfasNEAaktkmgg19yYyZR+AIoplMEbSeHV
fu3TqxzNCgD4nZhCuDNhgYfIJ+VFKw5reXKdwDAmTOAlq6iRK0ID9ogrpnUJrILA
Ya5NxnicpVLWqI8AqxA2LHNx9nw+WBJFhgwqiSynfDM8+15CLDVPZFeDWP52zPIE
T3fNGj5IxvSkotJNSVtQiCLuEpNPyIid8ZURcFS+QMqOmEUv4ipSAZmGjbDygU9j
k2cUWK5YGUaHhiwQnU1QWkytvt6sGu3mvAFrD0nEmNq5DkH7ECN+bkvrViKnfomy
4smAXHZhTbuSS1IJCcRrki3yfjLxT1MCePN4b81yy1WQJ1v8sNRrtNnG+6gc87NY
hr3lhKGCaKhavVu/yeLBM+zEF/kIuLwwEZBfF0WvskLI0mjgcpA0jH0677l4wHLl
7sM6ptTsbH4nIRYhrZ+bhm0eRueBvpYlGgVJnnNgvbdTHwZNZ1iw8901vJ83iyug
GEN3A2EEWtXr1k6K9tMscVHXe4AyCT4F9N/58DCUX/dYmBvZhpRJbSKToYZsb8xZ
+f02/jPCSht49sTL6rXqrAWtyJv5hDPZjju8k+VyhmqHRN6LuUw1cfPFny4OS5FB
MkZtW3tCnI5PPkex09E6wBlCS/Y7r60dE0PTS08Trz0C3D/sQjqXc5sW5u7oBey0
6X63jBPz1lM5Y/51fPFdy1ptrtzPUDycr62ppp/GELgV/9PXXvJdVBYE/vsMw+GP
URXPVMkzHMq2Y3+IgaLVhp2xxJ72TnWOPy2UssRbJLsPiSD8ExJiL4yNRYETHl0P
IYCEryy/ZPJsdKu4QzDDjk8ZFF/2NNFAxaERJiB57qZdAkWkgpRsgCy4MdEPGbw2
ZH5BCr4+thY6w0EFpnnBux3ukGcuISjvfQGEHp5mbVZs474oqBZRJejVd/zGejRz
k+5fIkoXxmkYrt7pYT0C9czFXLjTdcNP1sdG5qonkl8PGEWNJVKgxznjQl6FYgal
QDKCOZXRhz4jlPZNeDeN84IcAK/ZXoVv09vc6rtDEpsA1okQ+AH9zWYMsmWt7ADv
3dUXfTWEf+dHj+SYgchmTsdR/N08O51KDs9UU4x+2aFQHiWc1H8h7AmzRi88ecLb
/Ffj0hmnnoX559XAoZn/In1HvG9D9cvWgPk9rfLAu/OV8akP1NsElxzQAfwSPMt1
QExO+DsKWsqS25tj8RPXHDMQOEAzmh6Gv785Fa0haR2Jr5dD+4P7867Bk/c2a3aH
D5Pa/7AYGRdq3Kmok2xIYXpyDyOlKxRlW3pdkwMc9xCFzRxxCnhV1DRV5Kqu7rpG
kyZrd0aHM2Z9pXjyq0w4dEOU3xwf0RQb5dnmWZOtLDEoYVqPpeCBfHd3am2GCics
kZPOwHOO9qgxQVwvGRJQ4/OPBunuW+sMBWHTnhdTzDNw/sMwPfxj47F2V0UaSyd0
MT/2iTFPfBUgNPOjgVavPZ2baJxRhetw2cgL0u0PC8IETgJ6R1L/A1iU+5FRIO/y
eSQjuVj/BWsYjm+2KQqXY7gVWox82JHLk6mWGsJLY49sTucF0txL7l6CYgmZIeon
BY3bzftH1U4Tzj+1MjXY7ICOiuhNJOIeBrtAHyVrJctxdrFX3m+eX9O3YsLrAXi9
ovpVx6ypZq9/FcuubGaZ9wUxlEuzPvjLXW/Q0RxkztolvKsUXIi1xH1l4aNXmVJI
uaRBue3nF7VVnmXMm1aBxmjKp/NH/gyB7OsDpuJik2to0Y+QxCHo/5hJ0AoJY/SF
CBh/g0recJY+amLV6PIhSx91JzmuGmdX5pp2adnO6ZFiPdSng+c7Xz8PvPgY8ArG
zWnSuDChF/tV/+6+iWcaxsLuGgHQ0DpScN8t3xQoE8mbyPbs8yIKQGSB/zGDsUr1
pjIC77q1nbIsspLxHSHBAm96fM4SXw99d4rFKFB6hHJ1JP8zVs35LuoDRX0HiazV
eNSjKWG1Wujwtlu4Wdd1MofMFml9QF8jG2FlRt/zK6AI5qcDR8zOHypm3ZnW4SMt
EazIF1AcVwU7y3I4lhMRk3YLYRitQBFZ0O0p77SbkN7XeDDlYMq84peKqDL765bo
ck+tHGHXx98eBCAdJFEyunrJET/Dci2+DtPYN6BB7ldFDOyLSSbID4t/BkzTPGUi
+aGd4J74Gw9eXrYTi1/h7tUdv8Pfq7m6iLXGUwroZnVCyLJWXyf7uLko9UrkiznA
IXxqcxuoV/QDEAyO8xDeJJszK+/K6CfOl07KLsFQ0vH8u0/3aCNjEly7l7HqhPD2
U5LskuRL+eTbVWqDzCBi60NMW16RcA0MfOKt8xBSlwy20/ZRJXgKLTNGoQ8J7sYT
O/VWAWdFtGWcmCuM8552oshigl6UFUYLhzC9DMyoEZM5v/nLDbURozwsQ/hmG0rf
FdJt4zdW5tUKI89iHMpnj7boYG6DI7VNWmarjcliuYttb7NT3saSq0pSPSB/+XXS
whGk/Of2m0DnVHfPddP+MR+Ql5aOrqzY4Y0NyORCoTXQri3FgnZhTHvelhQc1JCw
kaKKvFFu5aWD9Iud2QCdyz/hmGnoPjqJumYqHlX1mokwO8c+NHpS8cQutkDNm2CN
n89rCUoFbiOqB7aW9Xt2n8uEp0Z2KoffXNsP2x/E8ZbJq5NQCxLwbMKU3M3QQ36D
W9HhlchkhN/LOKqHjGO93YvZ1ojIvfJuq9cNxegk0dsRAdYfDTiOrOsdU99cUv1W
g2VdC/RGdP0E9V27oohOByQt7Lr/qKjEdWmNNZLDf4aTS/t/8pGtnyD/E0vG3ATb
UFQRPYJlDM0XxdLyf+U2JpzDeFkL+9eBINoO/pEsV2IzBDf8KczBLh1+MiY4Cy2X
jZX5sdFAqKeQ+PGWzsG8Az58T1KE/yKgANYFPR77/eG+CiH+A0Xwwd7a8jUiPoWp
d2EXyTCd4r29MdFt02/v0mruAYzrjMHv7Jdlo2biy8K4pcGUpDU3MyRMdri6S0ls
Xny9GQiObK/vR2FOOVgjZ3BPyod7QsY46BJYAw/o0ZhSESNfRtdEYye4C0hJCak4
lTctuSmncRDJ+yp3dBvdIUlEzAaS6+LIRo5YuFSMReIN6VKTE+MpPFNYnT7LVNPV
fX2vgT6CbEZh/JCMnuIrCeS1NxhWLmkcAqr79mahd1NBQTM47HyJCj3FOcqj7Q4R
PwGN61RkXuTcLSuXn+DBcv2bpDUNhNnTPOwu2Fs3Ihh4gwRsJXMv7gfFZceWI+Al
pTdHj3YnspDLhuYBO+pbSKVHR3dhSsFNkpCKLqSYN21K79liO6uwIhP8ml3uvEgY
jVeVgODahC8QosAW136VdpgCFCxiUGPJwBUoO2MCeUZdI4nT62YWSW6W88RQ3oDd
rL2tnpMDpfawJsIWspLyFO0vRzl8jPiseElvVwAlub/SdRCYvf9bYl9ps43YfkKw
rlc27YQRCigKVlwJXYh/0rmO1cC/lrYnqrMliVgOImb3fagwJCw8t5nhh5HiesSv
StPKqkrmlSDjwYFsvTTqdMN3OsxAgK3Pnsv+88SB2rebmLIC8YpX6AFmcbvgeAv/
5ISm3cWWdjou5oLOikr1qDKm5pDhGE1dB2imhZ9gMyynBd9/tZ/oOZRabyEXRnwc
TSa1UkdOuChF+He7J/PHsHfIBchYxjaIxK1DqvCp2RROoWvT+D4Y0hgdhXmA8GPU
MXUCVNXH2ufRKj8wPe8MMulGIliYSFt/HYUx+/SJds3WO7CGGRCCpSCFwZzJQ35b
PIV/GBfdKUTzz9LkZ51bny613Y+Rv42IlwNWMtj9TOFhExG/J6vBQRv1JLO5HBeT
rNgW7GaHZjHe7itc16DsZ7vL9plYpTJo3PJp4NiGjDNcXL+HdZJdJzSXxF1DEHLa
nQOZ+y/aBs/BPdfW/18keSCWjDgOfzz701Q7w3mU3E4Z+Dbdsk/Gkalv/qqIaSJ2
MSo+enotQs74C3+ru5Go6of/rSxV1gFRJz+ilmHbehsXZkF98KqSP1damQj4TTT4
mOXpILm7p0KHv12E8TPnIg4qOjCLNiEj7K5enKJEjvgiGlHMk+++lOZvAeAM7JkB
d6RccP+yxeQjQaLqVGOhhXQKNP22BmUEKGmoaAVlz98mBW7H/0Gzjah/qqG6p68d
5KlVurWPqz3/+K0YEAuhq7UwjYbOoOtKGmnRccrfN3lFclK6VcC2RqKgO8+r15+b
BwWh4ZxIWxbUMOgeXsYmcZYXBcC2+BcuBzW4wTWkNgQKbifdNoeyTqK9GBMPaLuH
Wx1py0VjpwGlxPzYXQkfOlra1+8RTmFfrSil2uDguVZB1I5i6Pd0RcfI88hb6qaS
2hYxBOyYaTDrbKFFjclCTx7h8v8GkiDYfOxqImzYrX9evGUbzpJZFvL8rwsI8GKc
E0TwTqmNtMj/gYdJcE9dBKagZG4FCadMhLEIshXMKghEUUKza5ID71C12uEXh5To
hx8pR75qkfTfljWt+0iepvNqQThOKDKZOo2/AGzsWIEXsPZbUF4wJQFDRSrijhRw
UTTUwMF+srQeT2qsNZ9ZT5ke926OEfE4tbZ5lKAnnm7rQaE0NObQXAJXT6sg0G2r
FJ8hrJpOGMtrJs46NiwJkiE+3TbZ2BoWe6BysHQIjCMVWugntC94xCH1yOVEVY6b
gCnRkUw63WQX/UBPzZQLCyu8JBCtfGyIK2xhF6WEYD5O4xwmOCU0PnmadZFJ+pTd
dTkA2OY5c5bFXiY1cUfSxQ3zWMaTKRo/2aV83XiCb8pz97StGQKeDvgkngbWNKMo
ONqIBhdxDOof43jR/t1e3wTFOJtstO8B+GVdo4BTPyWmAVvb8BECqOI0KcPQlOK0
PwPeqKRejI8oaffAxse6zk+qU1mM9jr/UFnzJ7PoyeJW98P1STnk0I5AyMlNz7bG
DFb5aCf7GWhornglLkX2al87rCVtqVGQ+qmWq5MBn/EsPkPCd43BNaCucoMc3inB
feMQV4rQS0ND0Ogv+WoiGlLinsBrKUSClQ2GDEoBVmrTpB3m4e+aq7+OhWzZJ/JN
EHPqcsmnVykZnSQi7rUp79iwp6tSSGlK7Q7DmnYVu07PYa27ZT7nKAPbbMD/F2Qj
5MILkqgvaCad82vgmb/6vTkdSjUQcChloq4iP73a/i57yU5mDhzT3pNL2UvBWjeD
UAAbUt+t+GhOJiRnJqBvToeQICY61f7e4hzxrDYi9Lc7rZbi0SiOi7bNF1V0qorA
Va0ZcF/9gstoqNFZ4286SeszHsFhDWQnaCJzSCqkRdsu+XqmOpFOowpjjpQlsDVR
Cw93rTB1eX9KLak+/cELVCg//M+069WwyZ78PH1D2IbrcgobJFvuZN1Q9aqxYQfm
p1bssWl8CWBVha4SJjWzp7yZBJEdlpnsLaGFT5nyRSj2DAld5sSP5BwM2G+nQXtB
xtfMSckX1gXmSD0G8IDODXgC9HxUPB3N6ZQz4YT80DEw5fgX5vDPl64FVNdVbzej
8MfsGvCYpnsHnuLN9gStsuMKpkcPUbnA5It8gFCqdIV0EKZ/2glh5D7zS63yU8EP
+DlRxpS8TbBxo6nHrtFN0i7/hQ+HOIOMPioMfEUamTxIqLtQ7cpeWo079+BVF0qJ
0R25RpL8Mw6982V0I/CGIGZPeFgTLDrcNwa8ivKeSnCVBPT5mWTgQEyTP392p86m
yhVtD3A0rIQxu5B28I7tzt/LuEJ4WSLmIG3EzlgXClHTpLN+i9S6y8z/H95zvy/r
W9F/0zWSTbuwpKXnWB12L+Ce1X54Gogx8Ug3AxDF9gPXcqQqZLmZT60ZXsVZS6RC
oi3ZClacnWnBgEL40/+HgAr/17+2mJ4S/mjwtvX8Wp76DOnInh3A9bvr1q+zvWIu
auFRDavIJQQQ7qAmdTLe2x2fUrE28wvnPU5uiBGM+ZIY3KquvfnIzvwkHW1R83KX
GyQlLY1WpISIFCppOigg/FDWGNuz5bmC/tb0KpdemGiy07FhGyDx58G76SDfMcxq
ZBMO0U4JylIuEqiFjjkkhjUOTKVpgIZpB8V0RO1DtBY25KQMh2Xv3PIVk3oNNCy1
ZJQIdUzik4Y2TMr/yS/SkFTC2XFtorsFqOKAy6MtaPodULbh+as/5PKQ/ibPd8E3
6nqH7fNn4pUlirfKDs1z+iVhGo2aJ8DbygM1qySUjlHYgS1elGQgYOZsXuYuzHIe
iiSZMtxL5k0Y+bwb8O59ncYvuopUksb0LztD/9Y/SnD8lR6yrHDrug2jSHeyK4Of
671kUMaApHYwgE95wn4nVfO7gX2djEq6a2oOJqpT6vcfckUv0HpMq54RXqEZIffZ
F9Q6WdwXs5z9bwMCVly8n7F9dBRy4nMcWvTG5wc2fphFFXZ4fm9aLgcdbsB9cl7T
//P1SYikK7wgYtEH+TqIOUHY3tLsL98dj/67h8N/YzFnjmhY9v/5OVBVBs2K1NK3
jn+0tKgyXXnmVVGS9u8cIYECx6QJ/ZyNkrBwaDg6xLVtPrcR0ImSL3a4eVSP9BHl
DWZVVgZr1B12YpEeMrWkcXw15cXHMO1NGtui2nTNp8mzAHGCGMwMrTLvkMdTUoB8
zqmkD5TszYOchC6oDJXtVzd2Tio8wyQDml0tmgeOP7H0dhcEAGQ57ikqZ5ZdgOAt
MFM+Mx9kgzDNLllPwD2dOaVrfQLJIhwdRGGrq6dUAPExZvOhbqN13orvBubePOL2
+unnwKE0tQHnSoJ6s/yBhy6Ke38bNEG/+rj151PtAvFM41oqKMwBuZOZggmrdf7e
gkfGFiBJuiE1/diMoDDHjemwpWPxY5Khavqe6nwbA5ewIg1DpmRbAxhqPBn059he
3Y4QBGej9FMrBR1oR9NFiF/AySLUiUXA/OnTiK6T77VnROpoh5q6hkUT9dpkUP/p
Ce1p948tb000hmvLmFm7D4vPP4WtHK/9kLl5OHX7L2nQ8dOb8XGmV5aTsIaK9Mea
/NQH16TWdmRngkUOKK+upUVBvuvgksEaOav5NXyz3KnD578RlgYbMmSp5N0qW0iX
wNg9HutKI9UELghncBYg46DdPOZl8vlEN3qYfjha5JGPNFa51sr2zMPlnv/So7a+
HK5IpDirN4Q3sKfggLL2qZaxorE8JCxp9IzaAcFTpg+6Q1utG1Nwe2EyDSxxlC2v
XUWRJecbztd+MUuFylW5R+CnjnJNLlSy+QVdY3PPcfHSaLmzp4FKh9P56Z3Q/v8L
GU3nj9C4Y5J+kpPlLkpXK9TaxAyVkN0tWdvqTRMpdJmCpvE2F/6CUDAiCR5/HZgu
hIkxCD0Wu0HO4bELM7RpvsvYkrrdBV9jU1iOyu457oql+xet5YVgM/txugeRKOI8
ZeevJHPYwF1iQAbGsfrTp2He7ObiIy8Z62yi2DIMzoxElU1+pW4yJ/LVM0QiQOXp
ESNiu5ZcV0c1KJMeIJYN1QZ9P1/N6aOBkBqTJ61oW9xj3xCHrjQRAKOywM9KWMQD
9L24nM0bRJafANYYH5tFrpwJadcatAe4+eTpBB7/lHVnLUpT6x6qmE1zeHUKKkRB
OMDX1vVdutO6irG5PB9j2ipujkdKuWXOTqIQnqFR5g005EF36dy1Y+4KC922Zn7B
UchZAZjGz+Sn51hDz/TAWDjlc/NDK0j6FuOSOz75qwSyOIRO2fpW3z5ZP+v7WWy/
Id3g8yGerbHH7tFLeIKhTKKc+UsCemCFLgW/0zmYIb/1fLsnXqPFiQ+pSdooql0Z
YPgWh+aWuwTH93akBU7KLplJT+c6sEQiMphO8SCY+hnh2q5u3PN/4+8rrzIH95az
WuLMpV/YWyBe2L4d+92pvAFJMHadEKF3bsWWmrqYiZSocMMnx45a8d7QpWzG8Jbz
uDA/O9MwpcW5Yar6uE6wjcOL73pyPYzuTBMJVTzWHfNwbyjdPgGO/0byYZQ06ZAE
JjUPT2iS1h9Bf9YVHZCweupPXuapEgpPUEHQlRsI1oLBL15pQd1hbx5t3Q5VKrBo
A3wR7DzS2YTcGFr3nymBjZ/mEBj/LtbVIZmOHRDfHVQk9LligZ6sJ8x+6eHkzpHh
JBK/SZwQaNke6de9Hi9ui7uFwi1ELC1EwR0Ebs+vDn19vujEeJ2rz/oQuVY1/RaM
wg3xHyTpGii76XpFG+oZdu+MhLA3Fe3n65v8MTAGvGCSyaxCqXm5EB1g8r9BQAzi
IAZRS2MRT1ek8wwc0RAhVIEY0JFWTGwl5V3eH11TT/wfkzIkFD13HA+pA/KqvWQA
iklRrR1bYQbk7bNj0MzLiVLUJ5Mva1/38UxlVNR0MIffa+LHXmiZtpuEAGbsEZbz
udCwueG4eRdEjc7aDq8BUD1AhUdmYL6MVvjm7FcjFuC5Lsvl4gfsLwuJgHGIqqO+
lrqcogajKLGJtxsw8H9+fuEOeuJSnWW/QqIW9Pl1LlKZtkEnsU6i9hZufIqpNkiw
mIm7VlE+MD6RYn2Rie4YRUz9zOp74oi4ycGp9ki981bGf4di03dir/lFrZJSCx/j
Q4ewon54pGnWy94s+Z8V9iO1iF50OJ90WXLFe6k1e0rHE90wCxOj1YzOpyI11A0o
XXXcnnGx7sxW84MWZKDA23ZFzZQO4rQMQII9l9JGJqwls/OowXeptXcrJa0gL2y3
7HdQXKf+ziRkjttE7/9RxxIBw3+/C/O2GB8YYZH98zYWblC5uUtRs98zCu2LqxN+
T7wyS6jAgxQO5E4H90Fg81irdB1ERcj3vAVhSI33L6RHP2fPNoJtyK2cHeuLdGbn
TZZvL9JNdk8/tLk/WtD6sBOdUJFrwz6iP1asCy//kGxbK5XDdyoQviU9tU9AHKct
9U1Z/TO/KETGK5WnFCEuJTMTfkKnMASBtV+KBVcn6edcqmZVmqQlWdsIHoA2ipbV
IArK1duZH7BQSkDaFix8yMNVqTGl+y9mK5jixXIpxAqhXesxnbP1Rgdbtpfk88Se
xwprVHvk9Qaq66U2HGSBbkh+2e5cZmJ81E/8ncvLr+vygwA1oUp746s4SSJz85Tf
itYozEAHk8flfnFQzudWchc2nzSSpst+VvXYgeU8K0MpUUJ1Iwxwl8E2nP2Tv9A2
j+Hq79CLHU+NwPfWva0MGaC+6JHS7TtyY1HS4p2IT/AwdA2e1FVC4aHd1RMBTGYE
qI10y3XxxbdCrvIzE89cGjd+kjkaPYG6tCcvY6CMim0hulNujySo9B9DruQnloST
muypX8B3BokVV8WkvsHt/1zUK9fZjmnf/q22yJxFmXLDbVWE9Zo4UatUcvwU5w5U
D8CWqMtXZjTbEAWXihzKABGMrPyBYVmd1zKUTuLcusvGuOb6kUhh6wgQF1lkPZul
8fiylbrPKqAQdZ7d7G1WV5Wmtk5b0VpGjgEaIRXRjDAZAlQs6MI0ALHjNRZesOCM
KVPqGlc2Tye0Dvec3RmtvD7CEb4fOlYCuY57aa3Qyhs7VbRzzGrbwq0cKSyXLBvy
C2Amyjfdps0+pzYcRMWDMiBtob/8gn3svxQ+s5eJ24WKmkaaUm7wNJS1YiALyhCQ
8bR4HrjrCQEIIiyG0NsgyttCadJCMXYykP9O4jILbBPRXIBZFz32ArOj0P4wxtAL
CezXTpcEODWe1LyglrwYBOaBO6yQkEn7Wn/+ULqymstjpCSkZxVBdnWZ13MJrEnF
6kPlKN7EG0sa5bzNCIi9kFjzBL68Ug3XYQFdRprBdDd2J4hvdWvSfT7xSHdBK6Jv
meASh3N65+Qeh5jN/AK0bLT1BRKfqxsHuN5smr2G4ThPI3gnUquhsOZU+9jlzJG7
pC4yQZRuTNrt9bym8H8CcRctM03cZjBQh54Htf5MOSEYoCueVXJXpLKJiTvEpOld
n8TPsvyaSeeMsMqUGkgxVUo9W8UhQdgDBTT6wqGtE/epIS3fz87OwKKZuSilahVD
mZWATnZYfW8x9ef9uIkL18gueuK7yDsVZkEjRNJSt+qLvYkVZORH9T7FjpUL+HWu
09tJT/XJGoMMCMJf4fkghOKyvs5u4i5IwFUu7uIh2LQIQD25JgKeuIfaTZO8DoNx
9zWQw6sKkbrqEmfCuGu1Q8Zog6nJfnQBoo1lfsNfntdRLhIFhEYPgczO14V83aQv
zv17/DDGZyZxhRWxB5bs5zh20xgSoJzijBL0ckkOkRYHi5rX4Yjp0vRqTJFkfjtf
cb9c4WsE0VLLO5pYLd0RKF1OQSo0vcldt5lqYKrLxO1CUhD8+p1wijDH3Tyk4tAr
qAi8Mm//0jFJ37DffWX9APGE86x8mPaVLdY0xOQawxqJcKoTtsmR9TfdEl9WTOwj
VFqJxJel0znaqjM7aXeMGuyoOQErWwmS+XgojeSdYHprLjkYCPHpEca7hKYAo8CZ
ygIqcNgC4SdoZ8UtQVN5sTv7Tg2rSmCAxyif88ce2nZsesZCz1/m5xlUVPBdU/1W
iWH0wvM+cRIvynASpw+Y1IlLXoFaT/58XV42AFlGhTpY082XAivQguz2QSiS2PBG
PuXmx5WH9hATh8Ism5Ze3Nu9ol0heVuF2U4IRPKGoEehjDPtU0J4mxQk9N/K2LBo
vtpIrzk5o4LT/mUEY8fCFKhsFeEqSikpyyUJVqvTEE/a02/yPfjGRXT0AJYM5hAM
DNtxiNAT/7f3gb2kch0sPyiocA5qIVEiqiFk1uuykZwbjhdDIHMN2UfxQE8EuoiR
cJdkcGWiKvCixxL4m3hBHgKrHCfa2k+QbIG+f0/Usl1PuH9PpnQnBMLSn+L8et/7
TzR1d49PZ+vdRGsw2NuWFzJeO26H4KmhXd9KQix6xtQeRX/4g2mh/Dgx2HzRHHVc
oBSbzSM3JICSnvF4+yhm0GnHPV0EoVFGjk1w19+hxs0J9Cr/qlj4RE/pYYwmaysZ
D/F17SrqGfu621HC9A9KaDKgLJmZXpwvih1t2g6+Vsu4Z1E2yrCp3a4QFwtqXgFc
KvUIZ3CqGVDqLth4Wj10zSSnDd+lai3SURDxsdDbLeUuMg6LkNwAoJhj6FFkg/cH
RxXmEGZ7UZC6k60nOw4q9tgkNgfOAm/YeoaRzPI3ozyj52PlkBpnIVrHCg7/ja43
S6kyYYy8sBM/70klfmxgkIqC7bakSGonSf3RoOFr7xYehsjGg/wcrFt5F9Fw/8ni
8kATj9QvZBhsylfQVyMav7xiCVRSlTYkVcjr2kxNphx+ImUxJm+iPoApybkoL0nE
H9cKM2ZbVEOhcKBJyqtmJRF2ohNDT5t0CHa++/Vv7TqD/irjMvqDIMi2MYy6v+4w
4IMBpG4+gfoKHIEdXH04Zkeg/cabBLTTQZTbdXttswqqEFyvHREUUL5CKZVL26nP
5+ijH445lY5HXezOTpD+yrjj/QpVI/ThdS69J0XmxpZaYV71c0nAiWjRIr9KxBOt
E2TZkzLJeL5ABwUR5Q8DPIukD5Zbr+GrI7/kYH52AnTYoQQvemPulo2ltSK4YMnP
3/fymAY69Aa3YNtQiNGmQjmcgOSIwQ0h3IaDSHcwxGsrHPN+RP2c1P09SuSg+9hY
zTf71e39C+tDaFElh4XprN84X/ykFjRRqC/CSTwuufVUYgEm3xQnEulfKzRlEIot
TTnDmH1q40jmLbV9Qh1ILEbAexzxiK+d2bN3uFVn+HYRQUEskqhkKDORz75TYUCa
ma5Rd53mTeXpZxKGd+uqP3MFdW+IocHoFEaOuhhK98LnhsuEjH4vG6XcaZcRGjgG
BrgX4qpelmYxVMF1AT2WKt/FV27FIr1foCi7h4Gx0dAFdCc5Q9KGQ8Z/lWYUNrrK
R/t51LQd56y68i/5k92NS1s35kpXGPor0yThtd8sjIKGHrHLcwowtikvllF97cFZ
u23V1Ho8bngC7FH3bKqKRvdbp/Zs26uE0+zcRl5HVAghGAvUw11wJnuo+vldOxsw
QzGTCRzjrp6Qyk/a1aVT00oS6MpS8fHD//478QePKDMYhzqsfbaykl4SNgHTdHy/
EX/SNU9bWNR/RD4btjwtclJ9evTN1+XVtHqbLwjsouLwaHjSZlb2tnyQPrEK9slZ
6fp6oRIDwdf6f+l7Qj5tmZ5825ADrMMfPrACkLtA9S5BX94ASZCFC9Bzc3VBp7YF
B2cbQHiXrYrW7b3/hDMVk0BB5mFbEUAxMkfa9wIw1sRbVbXzuYHJMlhaWxuPamJl
us39G7CgUtLdVr2edlHC4x84yF4fM+zhyrrOMeYHiNaM9x5oa7S1O7DeN2B288ta
CxeI7Ses6vzHgyN2umaEXQ4rNvMQyPpkY3Gg09hbh9Dkbm/7zBMM5Rc/y4RtZ+FC
HXae+BXJm0dM/1tRkjhRD9mbtHi7loX3U32CYTcaKZ74Xb9eYIchIHDy0CnMpzs9
y0m7r6IoKlRMy5UfuW7N23C9NwZVDX2WtrD1J7rMQMnLd7UOsdoId6b4e6w/G7I/
zI6ak8wXK0T/Hhn1oMKhgjWJJbU2vwsHw+GKj/KyFeo796JQzF40/lygY/bdeEjv
TYpPA5Ny8xwkxEZYhyGvGFMLj5kUefHHung27VhzTM3ZZgg64t+PE26j82IujoZ1
9WFQl4KCntbWOi5AOlRhhDORxcVcPxSEus1TmXVqFg/FnYAtAZ3k3gNgxfPo3HvA
y0f0c1JOHVYbp45NutNpBFutQU2KLHfr4NAtEqPsXxjTYLsVX9b0/kuOU0qyJtA1
PYItskDwgqmzx9h0CNxL91p6I71cj5wqnipKkPn7LOhlW6NAOpP679QfaVOCI8k5
AqSKlsWgLJtdGSWVRPrxJ1tegZK6MgsFfR9K8jELsHSMS79RTN927UM1dC2lsNJg
xRamTJEyv7ddDdLN0H1sTsP8t+SZ4M2BTzoeNiXOKKwVZFzwXw03Yb+zKSVrLChl
tzYj+sfL3mLEo5g1kbGKzyqPo0wj54rhlE9njDIF773odTrcTOuMBujRtZgHneT2
E+tkILOkm0Qg+LUpMfMgg+1x2vPFTd66VVDz8NcQJvUmAWLvBd+i0M543WNW+wFk
+h5TnNuy82zgUvXefYA6ynXVLT9Qwl0gjGC3xs4cxw3iAxexLuuwSI7Rcbg5tr5J
pZmR9P0xeIFfg2mazsBZgfGxh2h/BA98XIeNeWlCMke3BnGenbStePvF86lgpMBF
XGzHjubYewnjlF06zZka0+WlgLND+ScIVQ6XG7xYXKGmPrMNWCUGAgGb84kHP7pk
CrRHy0g9bLxklC5oNCiE1mCepgTEwj+YDBBgB03Fy1oI98/m2THgyp+LniVavZCW
jMRu/TFAyoeiZhQjZwYSKN4cP3ez2FD46D7v59CO2Z42cyK3mqsjBDdfdYOCqcEt
UbtG88+DC455tTKbq055qmYrmfeIKjV28+S1GBMti/7uAnyifOCIf+XA7kTY5D3U
BJUVRovShJNCuAoowsYuXEixzrCp1XLwtPK2QmhwHvE6DGV7iLYAulI40LK089mK
sLfsuodbEzKJ+EvZR8FsIXVmnd7GFEiFGqv1M1C0WjzEPCAxwGjS9RQE28Tn1bLt
tBBeMMYJj1OpqF6cNrjy3nuYy/FHaf6jVAhF/cOuGWGcDvezpJ/PAkuWOAEhwi08
G75iE7HviE5IcrIpxuPY+aPr7GqL8a/pkkDwixS2Jr3lGUhlvEutYu27qWld0BB6
h6mHIrMAmLZHlsOQotzgrDjmoK5PWEaKcTnyIG1YNA5tiMDpaQBhWIQ7NAFq9kVs
tiBd7+PQ9SkIp3Dj4ptkQ02QinoVMLWJbUdLF8M/avbbBM2v5BJDK0sUCZg/Tr+d
HRGt62SHd981uKT+KzRvr3OYJRl8PttbOdbRNFENho/Q+PXJhwcbO15MCWI7whd+
AyLAuYnYlFcHI7P4voE0Vv6dDySI4p0/nYrQ9I3cu6yP9Ac8G5byKjuHGgfs4h2c
m93EUtLLrjUa6XPUd4eOBO3EzXIENmhpBabjjBq9VqAMv3mAa71GEbqG9EFt1KR0
m4EKja/EMRP3tE07cn2kkqn27g6aH/VkDTqNxB92c+4PegK+e1peseXJyeZ2Sk78
VA3S19cXkS8bO0VUrlHKDrCzhqqJb/ggwotQfLW67wbJzDMajhmug2dAmuSpKrLY
bzdgShEYfkqOG7kr8nJsMNd2Z6z6BwL+W8epOWBXCH19kOOLUibE0gSsj7b7Dx7I
TP/jvOeY0Q6i/0UmK135iwlgYKGXtpPy2881GCPQxPaODRvJj08YpYWS2xbuc8Jv
rB4hkw/T77LpE86JVAwTHxqDJ2XDGgrvmkixV4E24oTPTne7tGVstJTHy01keuXG
facIGXSuMQZcGTMA5aJzpPvpTFAJrO/LWmHpj6E9Hhkxv2FQf2lX7XnA/KK2dhKK
U5IM9CJ6plO+SviPmLILJ4rH+anuPuhgAI2C1bj5AnplIJowhHexPwrWzyqQXyzb
QV5hABAF945fPHKcarc7MoAfaE+CAdfBLaxYVrWpqligHZytKH4CmSgIRptF6fQ2
g53mfYc+5zHt892opREDiDWStTzGV3eYMWERYHDWJ7kqy1CZatOrX5bySDaoAvei
vI3II5RNpGS5UUonPykVFYuhKFOA6bPQc0EBx5NM5daDvs09xImYQYU0wIYVLDqo
NaW4uazzxGpgC0qagwZat5YPlOcgGwo46Hd+65oPMZDvY24uUWUoJuaZXVjHAu76
ZlMC3+jhwddIYl9DaczbDezIwUNegJMRntNK732VU3gvd0KbwBDYWGPiD2PxaxHH
/IAatigZClkI7SF/ALE6OJcERc6bw1QUVsbql8BRsUfYCuDrcr3kmAsgIJiQ8p4s
oFR38FRxp24Fgi4pQ3/vBK71gSlh3CrKewqkVZA3Wpo8MderttfJY8jlQ+ACF3nQ
RAmupyDBI+O8wKC1A4UutAc0WVUYnvUf2ROi8c2nOaG537G3RQA2yqpXH6U0sJba
83CLCy0fQXdyxAQRNnP2Hx0DMClg2tHv3OlkF8OoDThnz98Ro3sI9DAJB+j4I4jP
GpMpr67YvNgFtnEoA2PWyuv1j3qpL7taLUm8TZB3jGEjiBhbQQ6QyFREJf8svI00
blyT9bs2Vi3HZ7cjtCaK1Z7IDhHuztjYw4NSLzZcAr2wdogH2HK16bDx7/t0Ykw7
oorzlsZ76DXCnVZfEMVPiGQWm2sMuOefpMY8D68kJlRfzZKQL9Reb+9+bo8hTj4d
KCtJKcJwzRSlflVVegfRDE1M+4sKT5guUG26SRdDKGEoW1YMPT9WA3OqmHYBihT7
l/kDKjhsKnkrw2Z/MIsW+g4IhICcYAvZJoVVHo7F4fNOCbD0I5fnPdjjQvd+yalS
g8e73LVJdkx5UrkohXB4TH+/Nm4U89OvgJ3ZONmzNNqfoxza8OB6BmoRmJygFmSf
kmXvyepaaIfwZojkSk8wWfJZjov9CJ8IlefrxwAihq5AcQVVoiANtlLwZkavX+pd
pga5ehs3i3EV15zgbr39kz2F8LEV9bXWNZ2nWtENrCbzNZHymblwh4kPeYTzblQs
NyhGRYqmZuHX4mZnQO3Pfa/NuADblzFGU+A5SC5JV45ERlHF+q2F1qRfrrkR5NyX
ADQmMsZAEl/Sj4Q51VK2e9bhSEJR+nxW6slIluZQ6TDGI75D8aOmh0+LZfwdICT4
xauWJXTkU/ov72I+Ay68Vnk+C8fQLBXARrSIoPUpc2nrYBCGGY8oyyauMDr2/0Pj
bgiFdffJVNuKHl85kP0pzypCDdAA1mDig0UsR7SrcwTJwhZn6oXliLM63HRH0Q6J
ije6tmKhwJDKdoN/Y8P0yxMSjVP7nxxyg1y5h6SS4NpQlTLLhTHxc2CCJe5evFOk
8UPQLKOag2gfJi1/9jmHpHyK/Ql/mpQsfvZ+LhTZreURNRilqwohY1/mZ8ISIumP
2ouR0JbAkLpOoYivqUHMQLMgnj4VNizwalFAsmSVz6sppKRxtEoQDceIKHs/4WxI
YgzVzP5c+v9kiQm/v6flyn0BeKIlNsVR20ZAbB1LeC5SGF6XCZRH8GZaj6ihBPzq
N0udrwpXPmabFynhM4TGqr3sUIqBSZRE8jjKUEqXlN29LUinJZqsUOlwzdkX7bev
dwEsQOyUjDNpDHR1NS5r0gMcP6xyVfUH26ZvJRULApAcSjkrFR3Q9ZESX81ATCGm
sBMkGknM2kRQjmabuf0bAbAkpzbZ3doCSpFXB9N3ZuV0dYVtgiRqbqkdxbTCoYHc
lBp6a8dAwmJ2e5yURNvXYKCm/WEQQnofE+hqGS0YzfRvrAIsrYTkZl6C1i32zMEm
TBumuUkowiPomp10odCSL8L9lj774oI1nUV4gPaKLRbRp3uKI0yVZQ4tWTfkN4Mj
ap/8G8DNzy27r1Rhe2dUIOXfFCbRQRYje3zP9tOm1DdOhYKIqViAEk/T/2Nw1Vmz
XDgbfQjXRpUgiFJnEdk94yX42Ozc0ElM0xK85UJ/uS1NOfbNDMlmbp/D9OVDtsB8
EcL0/1r68UMAcjYhzhZTxoW7FzS5HcfEFYYrbkLXfzq0Ll+qHDK0bBFEwQeMKbq1
homgq5SxcmlqwHDYUluvddtIV76cMWLG79zDozsbRpvvzXD/us+baTd6W9uP1cpz
0oad3B2ltwFexCPcAF67rxqcmOZ03bVb1Th9r4GVr1pJ7V7cIsSnvYaBl87PNZai
klckD+0CENpNlVxrzzb4KuhkpVp8kUa0V2bUWUaookYpja6Gb14KrTMjVztdhCOW
xunlPOoOxMLV/ww0f/yJHg1ws4ChnJd+5mTOh/g6EaANkntoHujfjUcYZONwMhIQ
aNaoiZS3IGYDuj+McpVl4gVeXxEog8F/WAsjVRY3rjWo7ciX7MP6bbPhioQBPcZC
NhiTR7OAtiKAy2v8uZrsv+u07rVh7yj5Gb+1rZNXTBrzeoDzDHTDKhf6a+PXXggY
OdXwjvqOR0XT2mkDvYwv7h5cRtDEfTpfxyx8URTpOvnYaFE+TnVRXMXmjrcRdajq
dKVRoSIqoWFMotAbYFpLfT/pM9yPqBsWfdgCQzVFKdO/EVHiAOCdsFR13ftoa3SG
GS0DrsyTHgWKJ3IUvlkD6ZoflLtbvaBXvap/bROVFJKg2seOfKP0wh+4/9gGi7M3
f5Lme6EPmzPOelNKHPfienB7oH/0FNqUYNggYeF7XPNa8x6h0K1HrjnDgBnDnxXw
PuD1Z2hjfF/VU36333wAREhlcWcB4b1Wy4lH8GAQqParI0EKbFhc24YtWmYBHX4Q
oxIp6mJ8oR9VSqNFdVK4MoTboBv0HU3yElCFQvnpKqdtOWYo+bNFMNOVtw3eLh7F
TkTUUYJneLchdzABzwwmQo+DcULFWfcBlvnah8yJgI5mTf8Hws8iJfj6Gz74TpCK
DO05UAmTK2o68Qg/++Wdi4ZBzB1xHDug8IcD6BXuZHjk9gfDE/Ra69X11osWZyru
RBuWHpy1t/Anqg0zqRUw6VMeL8jbj+3uyVIR1ZEDtb6roGHj2OSdDeRjOG9HlSKz
T5SNCxEpYfhbHr75V2+8GuGlFsz+mCD4aQEwVx2hOys9Tjkx1CiiGZh/d3k/L2cf
21XxNnE3q7+giJj9tzYhhyHrKSAhO7egMAov5MFmH0+f4FihaFjcCzhER2gZs4X+
/8NLPOxC5/FsMOfH8UQ+NeB832LKCQ/evL3JRkJ46pj9ld4c/63JrTlDLbfsoV9M
djeq/tfMac/ggHt/MCx+PlD1Rf95Nqp9k9a46Bq6VWzcs5qEprilEXKZ/YD3QTiF
rATzDXnCiAyWqVIi7dVpecBoBljzG9MA/qvt93jQxEx1D4GDxuFST2lDKVccQ3ua
02JsAypmImTU5BG0cgfRXxrEX63v8rMLQedJrCMrhj5peOWbuEzQ9QnbEyHKtzv/
t3hqbPGAoEqPPSyr9qrpGxIAkK482Zd51+QSstlNXDZ1dtn1A25ik4WneXdc3eTS
oBhJeWR3l0dfC/qn0C+8bLay/7Wn+pE0NFl7q+ylt/LMk4Gn/hX1XjtJxfi9KlwW
mT9U+yxG90yP95yDGuAWezEs/DPm6lgDnTSF+tPnSZHYxHf9L4hSvVmePzElycAs
KsMat5RYcsFX1fT3tWdof/BXd0UqPOBnOflf03ZWnCXGwDiT5yArJ+8Rmc/zGuG4
t4mcit+BHtiRtCJJLa94j9nDgLYylojVmGLi80jBErEt67UOHqZT5iX5D1hvNeZt
ptyA2ytu4rKTM92qM8PKKwZMxFtdXVvQrvxabVhI6Mb2ZJZXN9CO/wdGc9qxk+4y
DJ+F6Ze6cDopujRmyGaxo+86hUyWXSwvbbsgUgL5uGGCUyWKWQqYTBasNl3BCe+Y
G5b90HQceRE7/AlFcYYfEx832+hwHd7IQPopKPdQYnoB2TJkHVBCzWnkhLj9VLdu
JTkmwzRQLgeg6bHYaxaruYj0X++/VIciYYJpHvNlzOhggoL0vljI6o3Er67UbGnj
j7t2llWQ/m/hNPebPHvhUQUG2aw83/DUtjx1IAM3pQTy45jr+h20ofCtYlyuMK05
vYznnkWFl2BVKHbf60J+4Nqm1IuVQfzwNx+VFtJTprGVRoyxPwdTWrThIag7G8Br
+DKKkROSO/6FRbS4Fno8YfbRXuQ+ox2K3Ng7lWyqrc7+UulBCI0JzqPwD7AZ4TdJ
t+TzPxFoja5tUi6Xol5uD7CboAtiDwkguwTZ3begnia3nCMWh3BoNLDb8CD5rElL
36DNfIenbJ3N6u/yqljfjAXrUfr0k5EDXQopQMGdk3cqXbgLU9Uh98JZ2nSVvhBx
+eSV0uPwtE2HgQuDW7pJ/IZf4d6vDthFs8R8Tnb9NyaVrWCakc8VW9kSpD//Gx8S
HBwwXJnw0qx+fOzLkNktDVeyxX0WXWTTf54U+OsxPS4Cs4g4dy1498KjlM/cBjEt
7U57ZYEieGB3JXeUqN8Ib/ZyuMpBl7VU8ePqCIB0lZ3GjKfN82zoZmFV1Am2iYme
tAdHLmvMy2XCtj2kwHv/E99m1RdzTH6731B9ShP6hQqUj5rDpF7PwEo1vQG6mP85
G26kpDf/CG/WyplEa0i61J++GbdwyyhQIgNFFee8jOgRl6qooPhVqZgs8YRRR30d
IXGlZq1bBcN82LUyVquAcIDJsNRAB5W5FmeBy+ZUDSuMxEJp4ZOFMj+2AOPYPieA
AyYy0Wt8Y1cbQS9uRk7qSW5RTT4j6eVn4khjeVus9AaFgpyuOvo3ZA9h5Ry+GJAT
z6UUsso52JslpPgs5O6/8ujLt9SyFCdtCgtr7ku8ivVuSF/ffk1dj1JG7tAgcAzm
8dMi1k4AeNvSVkNsQtvKdXXs290814m0lOMkf4Z04GQxtYAmn9E4PunLewBwmSMW
wBFuQi9u92eimJ0hSxxf0SDNNfzeLkXCGKR/AqjaeG0u6DVYtCEbaEbEXgadtDXE
rTJcyge6Bu8V/13aXbQN6VPpxAWiqBAQARNbrLS6KffAWLAgGST7gV2yXELxmRPf
iky4q66B4W0tzu1X7CfdpvEjK/mZMl78UvRvVaWUSLIwv7wN0Aw9BL1YWwINtEBl
jKgA3eXc9/+I+XmpF7I7RTrPcZqlqUQbnRKBjhDrrfImlaxhRmckRcDBCAq+AkzJ
Lpy+LO3DmDXSAyE1nvdg1wL9iQwM60lBVlhB4sxYNi0qK56vRJneuscvheJtGvQX
d0ewmbBgZ1YvHWW6HYdT+fzRopiitE56+7yPLpC2mIkh9VoyCc6GEQTKFW0CL3wt
bNNYVOUMdVr2QwME7AG3cXNzn/CrTbrOgCZwg7dPSbL/NJUb5p7JEnhpTJAM9Ii+
rKE+vCpuSSlUYL4BnCDk5/W4Bq4TL9LTK0yXcb8t19bAmDmE46Y0srcVdoklPfx9
xLP1WtuTBwzqWaP5dlEvQM1KOO7YAN+iFW7yYJI7LAyYm37G1VsGQ1yTCvY0zhu4
oblJul2Z1d4qAnDy3khmobZyiYJchGfPcKnQd0sBOQgXPbc1eOa8Pt4I2uqGUEjC
U8CgWUdCO9jbDeSv+++Mfp4pfjRABZDbiBjJoLjyZ/JFEaPbAJtDeCpqDZYAFlX1
/ZYETZX9ha8vvvkRTXpv8efOldCE/DCvnOLp8j8xMENE78lSpOZJ8iIRf46DiP3T
q1sQ1OEoIf4JNCV5A9RE2EJRs/8GH+yS8cd7KmQsuXhiWQ+WumtBm4NcI5rCrPQl
eEcy/bG8b6k3bgfkZK2Qke3TMI4LzD6mrRtoA1Lhs5x0ao8sEdN39CJH1O5l4DyA
ZXcg+nTmAkp76NvHbi+4S+m6UnBG+UEMYli5Yq/7StD9vPwrfEuViPlik5itHAdC
bOmADY8hn3DcFpbGdQqzZfFpOIPHfY3KlSd0FfqhRg+gNC4K1xlqxx5ZcgstNntz
MXYCi+EbnLyAp/NeuFbCTpAfemVTPyaUhbOokw1Ony/hR+LtSDF+rfEe5eXGSRPq
jhvQxPVCzd7D10OqXRpSFiwUnR8LdY4tQDEgdCVa6SxvEO9YZZYIYilzRWdgDsPA
xRo+YDvkwgTvcZ+Y6VQe2gRYASa4A1fdN1Qk9KaR3y0okWIrYCOGjeXiykdTl/PC
gblWN0liFOAFyh+yYxWJGzr7GWSMsn4/umXSgIknP9mnwP/dzAdWRTiLAx3l329Z
rxamg82rM8jbMt6xx42OcJHdvN906uZIvzaRQxs2o+iRD1cEGCoTgbyQSu5goFY8
h4s0+4+L6khEC2dXaSpPe+vVXg56ggBKjvQygM3wg+/yMbFAr8VGT6CnIKQdqUQA
GuSHoq/SWb8SrUh7LbwFqSMpf7rQDuycXiAayyYWj8bMSXXIw/TXFPak3hFJZpT+
znY32td9YSV+bnAEAZC+o4ySQRfJG/vjosZLXiB76uViX1xUqgS72pj6bWYVdDbd
g3nWnNe2AdHewkOvjqPYvguHMLqnAc6NJmJXENwAOdmsRxpAYZBujRTlk10v9YpD
+TdYQyRSauu5DDBwgfcOCmqETSzvzeFje00LoeA0lhW1G9C7tg7yZbNp49/1voH+
rxK9yQgHoEWWQbE967SvgKyoG9yjntlktOOJmq27QSX6WIl4+s4yA0ZzQGcDwww0
fMEd3D95RSRIcB4ZPnfpFOgjuW/q/hv6s/GkvpuzzwJ9U6Gr0nZS+J0Zb+pb/rcF
cmk9Tn/EfV63kNj38uVpPdE59A7OQYZz4zjqEc7KDTvx1r8vLmXtreL0eSpWgrWt
WzfcpEURnyuEDNLkqhhu3URWoY6qLxBHuyGB8sWB0MeD/ALPTlgvvc//WnzpBRtS
Fa+Ke2Cstn8nstMLcpghXgr0U41LQ4/7/Wfy9l7WgwBMU6t+58ZFTUWnfpwZoCSQ
Guebo0yvi1pAgre6ytyWQ5TArK+tCyODjeTsu9FFGz70pPt0Gqzgg6jLmb7QHVke
I4vrqX97DflO3AL86dlOXbUG+lIYb5N5iuBfaQr+kBSOAPH0R98mzhU0bjDmy7r7
rofLvesdh+JAW2iNdHuWHqfMTMTbReALtwsUoJkIRGicaTbljT4/C+8pLxt6/V2a
0xaZfHDDTDcmTCPz+iwhlyhrNxlQiH+q+5wYA0/LOG5B3Et25XX9MpzRIchLXJBb
NcPflzhSqghn4YowLLXrLgpahywSH/1QxJXZpUXCMU/qvDPmYduxXlKCs3DmWcej
CrE6e/LZshgB8CTRzJHxVKpCmNp+BZQohw6FiBqxnDy2latkTSoNMtQNGfEGZ1Nq
TpWCuOtGLxdC1Qzx9+IlTKgoXg2Xo7uxMPN/HVa7h8mTg9bIsIhyOZNRjO0C17fE
NgIWI9tmsOdgIO1OG8mAAmPDBGya0FhYkSM/CiEi8E1flgLUmxQoH8s9S7Ouv7bW
vKv6f8Dm6SryUZm4Tj1UedH2K+2Q7HlarWnCsagC1I1hO/MAhTmUiqlwyv0tkoHQ
OAU3jenhYHw/i17ouUqanqvRDZG7nwEICsqardB6FyGJJJy3a0S3OdQmyIPiZ0yY
Qiib5d32//HakWsiRfa+R4WQWmwf+WWBfsq1G8NVRL6RflL56UZrNDiXUx6PxZXW
S7F9+w8B9GU4oZnk7q00y0hsidCspxx83fBVT6DsL4TBWxbj0KmM7Y2Z2QBXKSWb
ADplBx2iEKP3teRoI8MYZrC1BBKLfdF05NxTLl7y1uw0TmYGOEnJf5dLxn1JLDSy
VjAJgRVWv9tYGNOk875iosz+L639C2vas/qWP3tdN2QQOdWe3L4vStpFKZGtX2yR
xdNMMkRHxVquv90ckJMERm+L1OyVuPc495ciLz6Fv8q6tCHivLsZjc+WOTJVWrIz
TpJUbxkJCghCEZqPTN5NbK1gAdeVfDAX/K9n9B5nM9uzPqCeUhmUFe7Lo2w+u0x5
BcC37uRbqOFB7c6lWyXgiaY1rWnYh+E9fWb36g3EBFR0YLsQ2vpO7QVOtyXrTF64
0qIGgBsz6oX6hX3EFpTjJqkiW3OmAwCtNnuH6CuhfsemDNAfypLO+6cx13TXdqma
Zmut5ZngUHxlxtW4f9wiBvmJ0Mp4GAv1WSp4qB+9O7h4D/ObIqsui8ocdv2hkKb2
7E8XYlw8BJaZU8XvIl2EcsPg9bBuFvlZ3kM93TyXNrQxJQ7A3lcnFAy6qt7RgIoN
HTWGFE9ICVm1ZOWkaJ9OuD4FDaX11oVXSOP3ku9VwOBiCsNh4pqjJOl0UkiHVUi4
AfcGpLK9S3CfGL+BwtUzSdncraaHa4T75OJbI3NYkHyr1DFORWQ5IvNLUUhB52WC
HHAP+PR9RrzZWcQpo25tYQyJu7eNojybi+NsRXhzJiyBK6BMjEJsOhIE6QuZKXvO
yucQ4xhrJ8V1V0ODk8KW21ZXzWZrNQi6+CAwxM4SA5FThkZ9HJFJFtzdD0NmMjbE
EB98VyqKC76ZtarlqUP2jFJQ7Es+AiiKtTlUaaIVvFbVGxgXHa97Uei3l1bQg8FN
1FpLXndZ5N87KimdrvzXKI9z7Sv7CDpQ2AGoL9f0lKmZFgxhX+XlQ4mGxQnAHpRk
bGsGUI6G9ssFv6tFqjENFwVXz9Mqb1UvjtRFS99jNVDBTU0Y4LBpLnJYvlG2G2yQ
fmrpp2NtBrIVRWTAbL0Fz8UIURoUWSi5STNNNyYJI+1/UNi/SWLi1MEy5KLWImEz
pS7ErcVfYrKBggSL+NhO/RP2F+pQEXCR1iHAnAK6kbmE+N5jMQPbTAAYmcQidVHW
hZNOZwb2zGpCmb3RVxb0Mu0VVScQg2e5J1DqpWi7dAytgD/O8IUcCCz4OH29CXl0
1ojWYOz3/1URFMp2Ig6jZV8LXMnPvlDBJirAoZCvxEZCSBv1eAyHN9o35t67VE5Z
m/BNdU0GjjeB+5ftx1zwmhJTaP6O43LsYp/UEYPX4S1zTsCbGwmHERgWOlvTPdpJ
yNv0tTHEhhW5KjgZ1QD53lYnyhfZzAxbl0TcmiDMfEqqjxvdLk04LM5Xxw7zIlGV
W/r2eRyzr0dHsStWGweTUusRsRHSKvAjYoYTStJ/ec/XGo9ynVfvxQqiuQzDqVof
KmDhCo5WarTxEHz4Gp05TLsSt3Stj4Poc3enzbyaEs1NEptH/46RzFGB99oRMlcI
MszPn5KUuDGxoTLHoZ3IRigbTZLXh1i7gyVwzX/qH2Qj8uNnkc687NrFbnPhwzOY
MUw7WxwtAfxpVZmPoi9RsTqLTwBIblA8nHm9Sse3/0152iFY3qSykGcqWeaWbVyy
yZHEy3I3EAbEBrhkjr/dhpEM3PC08wHbZZHKsryhp5Nl5GDIOaFMEKC9sqWf9BXO
PN+F9Daij1ja+g8if/u0upnxag24JLrM9umeI/tGh1SZRrx+2wjWKg8MJDKIiGaE
I2Co6UFIIROCNMeX6ICm4FM7STyCz7EkicO+lVeLgA5XKVlpxtjkc9TMfkRF7kn2
BFDI+e8tlPaZnNlDsWdq2k+Pv1H+667YRjr4fkJoyWBbI4mNI7Q9FCksbP7K5uDt
sgi0JiWEHWClpQs80bb3kuURnayrjPTXcZG83+8PCel3Fmz1IZ43I9+A7LJMtbkG
hWbOLg+xC8I7jwpbWhPEtVMz4ls/NETxe1m5Ln2P2d0X3wAciBHrDh1B3XM4qku4
aEUEt9TP356AnN42geBY8KGzzWxy1VgNCh7eyCX4pqDAzBruBF/3N9LjDDbepQop
31iIFWooqGzBtFjjqzI60E86oQGTU45apVNgP/rW4WM3EXBbuOo+NpxY5LB4UQCw
LAC40sv6Gh7mYlfxvDx4EeVyjItgotB+uRa+cp2zz9ITzViNNw05rGRZ2hsmY9Yi
s3qkBzzzea4JYwzwbLWc97lZZ+BVqf1ZD2/ktl4N5W+A4h8RpwcZ07uZXZt1d/PN
oQ+1Z0tRw1nWaW9uwWWR2rUzA1gc2gGHz8vKwjzIvbAMs+cjlKztdr49b0cSWai4
IOpbvQZHV++1meUq3rCHipVCAtcdJBfsb0vguLGcY2+rhxCNp+l87X/5PpY+7n4K
v0f1HDrOOeSQCKzjeCEzZ1gychhVhaqvWcUPu4FHU1nI1EZ9T+oX7wmHJqsPJU3u
lYGoqIpwOhA3iBnlXWYlla0WMEU48U17u8wUepCGcHoSyUtsT6DXxYV3DEAQlX18
T1ZUj3AeFVRMMXJXQZtg9/ry3eG6pyHKI64U3q3NtJLScO3QlZtXVIMfgJcQH+nF
h3tpcw5GBz1e6HwzBHyl+uz90ryu8lkpXDKGNiI9V5UTnvaeiZR/XKWPvXmjgVvk
fOQerc0Tev77BmBjtSR1HDVrhJhiR3tQ5BKW6snFBD0kIOuAfLIplPsiec7BhmYZ
CBHA6ZaoSR5opOaorkWqYXWBRtML6251hgWnYdghaXJ1GhUn5RUp1YPOm2BkZPsC
ZNTgWdUrMU9Wk51aAn/m8Tg7PKu65KKtnE616hpj77C9rAjOYCPk+PCC+magrPeO
/xTzR/kn6V2fnt6bI+CDaSS5EohmoX6I6objM6ual9hcPIQWPQCsx+4Lad5meHFn
nV6jfnLylcOB6B73UZCNWuHNJCe1J5+BuA9VpkQoGHgP96FcXQ92xMZTEpd11fDO
Dp8tmwG9Otc4hhCnvd0q6n+2adBbRAQ70eJbHN0qBBVNXIPHDvn32SDPeBw9tZk9
Q9W5ACdbT68jWnXjt4cQ1PkopqMSHh8bt/s3XyZzvbl26fi2FXnn2XB5kvYhIItB
sJtcT283eJzv/LgZtR8Hv9MezGpMbdL4lPsdPhv8SWtLQdweyviAzp5N9siGtIMx
rTzK2HmznGBMYWxXxRTjKhaOoeA2hA4I+1TeQgrrogF7xES3261TzKM8mWUb3YQw
aJvCLOx3cusP0HvvIfmf4IQ41SfBnsr/L4LVX82t8uLuaFRZM3gBBDUA0eiXlKs/
myYcFyy0o8Oeytn2iBuLhTKr4FRtgHCqfs6HvYU0PXfivl9L1LjWetVqWGwaRx8U
nX6yUNodfV7XznvuCVtulZhsL59v6DsmCuDb16W0jeKlc65y1JK62yAfJW4kqYui
qldhQ8Sgm5KVsqF7KH8fugA0EcAPhMoXpbJgBquFdAgbJTG/2Xql1tCOb29PDxyQ
PEAQf8i1Iefef72Z4flnnKmUbfvgVIGqW1tSYATW9ca1dSmAnduln6/VW4PCAeHC
600aIfBUGfxJUrJytYU0n8j3OHi8PMqg6iln2f0itQ+gNp6RMdGJK9Ix/T9g4vDm
Uxx7lHmuIn+5OopCrYyHG92Ea9d1vsSWj3wwIBfb7gZavVtZTLzKwbDSGUemA/n5
5frD7IZxgj8IqdyndwGKkR/DHCJO0zFJU7iWKR4kujb5uRVg13RHgl1hHX98HC1v
OHbMr6zjiGYhoZy+ltDtF+7XVI9Vt6dP4Jn3LlrQ68vvz27cBxLURPRu5AZvgJE5
jcW3VNQfUNw3HBZ/gFSy07JCIebWh0rhuR0T3a/7MRSoQp5rCSqu4VVUoiCfLZJQ
zngJi8u9YIP3fvddTh2WDr9Nq/nOV/5+YoLBPBMaSr/bptl6VO7dreCdYftx11kS
/kc+H/rlWzLuzfSpG9WxUJL8SoQfIZOr0smOnNZbY8YXGRhwM5EZzNUi4Fka+sEA
wtIUjk9k2wGH2pGmuBtmxScGUZTXRlxvmgTSmlylhixIxXNY/kPFjT+eSVP51h/h
H4OHY1p9z7TZ+EEhd9ECahty9Ju4dxj1j4rizSCDN5LPco3Zz51B1woxcSplpZfO
MKi5sRbX5pDY94IcGQyHxoCF+z6UA6qhRfffLogOZTvl5rB7TxnMXXclchHgHT9C
EHEL9ClZaaNk9yGVGoESqNaOYJV9pMxwIbjhiN6wDyF2DhjELIp966UZDudpOOn7
yAl9nFdfxqmTR2hfMSZIdkrmefg1JjscxV5Oi9az1G5HmQn78XFORxBDIh3y1hqV
4Lx/vG38hG0/cAlQIAPoR7r44oAkGn55Vy6iNEskARHPybNgvg6qBx1RE+joAw1n
LEsyLu7iAlESdFdaQFYLjWrXeFkPchp5t8nzPtmJ0E+mcVheFei77vsOOtqjBkls
SjNnuERzl6kUytE4IOAwBkzIBGcFPoGzGbZDeaZ5VfaolG4W/k3ouTWUq9xINvzK
UnTVowp9medkWUBGNtZUR4IkkgMGkZYxopC9S2i5g0gdPHCTJlEfnB4mEXI85LW0
5yESPGtn3zsxiQynUR+lrWpS3lCsYOIWTJJf11zx7SqvXINITsUnDckq+T06Crt2
J9WBkqX/PnRMTfH+5UUt/kRTmzM/36T1h4Z9/sdx3wmpu7BLbxWDbbShxSXOjIKG
HYwGA5ya40AYoZffo3j80ciQyzceXqJRAnPOvwmGHWj2L/oKVuBLkrlF6owc5tZ/
goWv0fgoL8jPt4ZtMydH68dniNXz7goW125tKV0bXQpx8/HZ0jSo3XA1mD4/4GY0
KwopdlcGVWantd0xrXXDyblvmBgVkIFIz4cAUdCTfKPyLyw/KH9m9MxMOZq5f3jV
bUH0IrXmeUz4p9Y7/CHGkBKFSvRB8sddBi1gq3hG11x7A+eKVnVPlrZbWrNbjK7S
MRGvgRtriZmP/PihbxbyIk4bC/G2AhjU1ybCz0nLcS6nnhyTMBlKXYOOR/tFtcHu
Nwy6tK/MpDaDKUxQyAW+/6lmS+WcGl3trg4hL4nhkltts//2OYU1ZKFun5A2krbl
dsje6443UpRAkkbXX8mzMXd/RqFwtiJCJc19zZxrmyegMDQaPAQ+Y4dtWmccS/n0
TFLgkgN8F+bt/VJbvZzb1uJcbRIIjW88aBpuNkhY/0CpQYhtsHONa5Sp0RTi4H6x
GjwADlaZ5lSbp1yYpedzVv5WB41Jf/aYNcZQQQqoiGo9CoHa8b4V0pGuVyaZjkUH
TfNb66GZAkd91Me9wL6Lz9uqMCBnDIQktcXA29Wv/pYMd3KQn0N7RihEovddfkDR
auFUK201xqvgnQHybRuOds/PZHsFmQd1BOJzAx/n0mTZdLgtC7Ukg/g8/FEdDjEe
L6kW54oHyUzNms+LoQUB8vZsSOantLXqfWJbOpsiZoF0RQNWmk1JoamjHPHTn/ZC
R5MhQjl42Oz2JuwADc97+ec1n+KQobEu/7kDlxkwRcULNjRLLpNDpgC+YYdPMO0I
TGF3MCRDzHJxj9shtv36xSKWC53GmnZxyC11rVzslihBqvpcKQMMPx5Uj1YpFN3l
Nb2I1BBjnV5xTMmKpXP1CapZGHWmJYQGkrF9HIj2iBbsYkdHdmHPLuGfXYB0OQpy
rTnjPXhKBF8BwwNd7fmeUCjbG6F61qYC1iHzBnZn80GQMlOfuRQry3f7Ds3WxwBd
JETIZPJNkYm70M5cW7cphTUVLXiinMPTjpAqsmoY3xNLMQ5zm7Yo18XzHUp5TRye
wL4aYsYaKrHY+J9UezXRo/xdNEvsKfVjs7ZnEcw+io9xG6/m+fTwxvZFj1y4jEJ3
pmoe5KAYiws7aDGhIzXw1xMlZfyDm2wd+DX98olWMNZ5iscqY5Q7hzRBfdgEdTPE
vew4xoD6uv4R0TjjBOgMWlhvNtpcmQjj49lUDACl/z1GCEG5wSOo1vBTn4dN5ly7
/J2Sljp9BVBcqmHbikpV+tWo0REmnJgs05V9rgyWKUcKf2cGrc61f+FAqFqzLH2h
rUp7Yx/pdCnM6PUfVk57lxY8cFFx2Tal2eONUvxnmFsNwOkIu6oDwtMAXLpoNXAz
f6enVQlgFiSWo2GXXfmUub0TvDDU0tyoODdluWvLz/p1BPCwPRDp7ZmV/5SgeHaJ
vcIvPVZkuYOhRu37brNISk/CCVnv/cA7TFti7IBwPm6vL8q0dnhPGJxNQDaaPicJ
rSRLmbhbcZiEjHbGYsmnK5IEVuKxdraCb4wNBmURqrdxW37g7AcX5/Dt1S0KWI9G
KNSi5FUa6QeDs4RTVTDxT+OABokgMyJViDkx5RBOKrcT8Xvja7fesBaasAgCj/Wb
h64kiSckmOtgzGWTxhmNRcHvxjXQWXoVk+sbqzmjrZ1SsaOThjZBGNcVHWFbu0vr
nkDSqS3itRcQ6gd1AbFKAA==
`pragma protect end_protected
