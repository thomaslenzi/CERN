// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Cab258v9SSTj8uvGAjG49Pd4pBGs8CxKFFhdK4SlEizcMQYFuNuSrAvLK2k+/XRF
dB3pjpN0aT1IPrboLecsB/Ad98mAaY/o2mrZV5OteHIL2YRmaS9wf8dDXEW+XMKk
z0l4TQzSPJpISTXsNVez2NKLxMe2RaY8z+CGnZnJoe0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34000)
NAo/I+UkKvly5tT1m67upsHuSsO9tP0OJra743D/HZTMR3X52kzN4hTAxjZ+esRF
O8sF6LEZNIxTViJ8mpNSysW4QHvtiKeLE6mfYZeo5bFjBDtxwVffk3lHniGQl7F0
DjLvqhN0NVHMFu7I/uyqtQVRz/yXDmFUrp9LbRv5L/9waqbfeSSJQRKHRdFWhfuQ
g1yiuUJX6foqCz5xnqItjo9z87MLhewJzwr5stsQhspohExA+sBflKe51Qrf1RjE
eBUYzMl1W2iTdI7CTWZS1z+NP8O0hI7A/ZFF1ZZ6uXOS7U3hr9684IikzELltrZh
qV6KZECBAYGoPBKWppa8CObqG001jJV8wQ493WyFSlOl4N1U1g4S+UtEYirvVM+G
4PyalcDYno5JCMYFz1UTNc3DODFuWSx2N438gMr9bNQPKIzFwZ1LazPZDtwFWAX4
JvFTZuR8E3JdpZrpPmsLSnRrT+kG99k9m9u/D9BhIs/KbKcgAcXjSF5UYnevXaOw
Sbc/lTcy6pjWIdF7S4xlHg3SMvJHsIpaYdfqo2iP8vM5rLo8wljeLdy5VfHk0HRE
zAC/SQ72LR5EYfl00A/jThF+q+sFX9S4YIH2u/xF/OGjTxCfYOR4Slx6Bu4ZDhUT
rTnjjyaBSrZV/s9YGGchsSMGIDUOnOffCYDYYK4+QoiFPw1E6Pti+G5p4Qpk6S+S
SZ96cf45ONyYxqJ3WMwEK+DbpviJZoqo/mAf9UMYJGtmHvXh7HlCQCS97wZ3gZQo
jq6iqkxEXGq2ky2g7wp/7SZiVXYX3Ch8rum+GbIHU6pYlIi6fEMmKfmp76LumRnm
qpatFeq/4OgV2AI/yjPrPwfoWquRfH8eLkKEFt8j6+IWqMujF34lc0lSt5IV5CIp
eII/8io7ThfVeWdO1SZqlt4k5pE6HZhpnXLYzREt0akE9rR2W1ARfFdyjj1XKVGg
aoD6fSeB2Pr3r3gXdEEiSt2c07nO5PxDVnK1Kjrw6vKYlrfzlt2mtbv6spZ7kdkB
+Gwv2P8c3oLUq/KvGlJzNl6FMWpLNdUd+Ur1yeSqK4uTGUICMPgc8SIihE3EF2cD
AXoE5gVPT5zuwS+byBwf84KmCh4emwfXowc+j/HBEFpwS6J+Ugs6Ay+sETpMeflO
lZFChdrDSM7r9b6mIXrnxQ+jHC25skO9qL9/7X80qQQZLVEFgjlm5Ksma0AoDoQC
pOU0ftpiDXKHY0oI0+4dRm/RVFc7Azby48KVF6VuV9bze2PbYB5M4nj8fkPZNiiw
XAA3/QrSDUTJsld+lCFNyvZ1XK3Qiu0Dw01KVK5HMGXnczB/OA1wRMJqSnkZeloU
Y+zAcFaWF4bIcWPJSkAIQJTgzorn9COKvNXBNiGOBfTrBsu+ruS6IaOpmWFD60q9
TT2TlrnQi1KYHSssMweNn1x3r1c0KGgxrXKS4Vw41k8q/SiS60w2L9a1rMVoefKM
HMHL7ZJQ4eL3arhRuxB5biotHVUC0sIkXc4OWRPXiiHiJr1x/lupvhyYpoo4Fjw2
H958lXFXbmm5wV3vK8hGJb6SFaCekIRQf402/yrTjwc4tTTkNvt7t+32GAWpiipb
8R080fxXPx6dWMzUEd+VuJygmVN8SAPnaBzFeeXq31fE1YT4R+3lOF9Hqqay6mTy
cyyXNKv1bQnkDp/WNv3WPN4gJiT72pbDAmkaAtPFtvCe7gItWByucgp2SeOLQuZ3
W3fI4qiPF/3aE8WccOlAm5Xx7JpuuKUm8wjce+ijhVYyfnLPzKVXB9SBPLTlAFot
8mwzLlfd6lMdKrNUmbVp5fFd3bg4mKFWDcm6bZXAlIhpybOtIW9Ddptgr9bEcF1M
tK7n2TnxAnVnz0nroAo8rCcGjxQwWMtos2FF7O98qFVfiA1+z2yAESo4oXOUfIvi
vcVySXu9zIIzT6xKhxCoynjlsvCmILJSF59+KN9wlu7c8CfaIvXghUye2LDIAMyj
Y71NiQCmfub22pI98OLX0el6RjIs+iLBLY4KhLKqxnAfrKCb0pD2FZLTrKf2isZJ
CWTA0dnd6NnpWcYQO4uS2j73vTekURZbVrlmyTWEGhdAYdJb1K6mDSDbXBUuncSI
hN4IGTeQbhKuN+weauUBKqfRlCQxjYHcX6ku9g7rvVZc6FG9uRwlLsgZ7NRjOgZK
L1wAMSfExMy2Tugy+Wq5Tne3/xb/4jx+WSDmgMHdPbLDyLRoPz/0o2qiT0F30lAJ
ggUvlSmGm8kREogvRIYCa6ba4kHzFJ/vJ3FbzKtaEQDeCI/71G/zg0bJJoSThzMa
L9XDicbhbl093A+rlZLeApL10zXlrDH+qHSdnOxAIXYpaRPfb7hhnjHw7CWSzH+L
U9zimwSzEkceqPAI8VwgeXOX+8k/HSL7wrHEAg0GeVGzBTjvfwdMFcLD05UnxSaO
rkNyi/lFrs64nvXQKMej9EoHxoLVbO/auRRHC8SFYKN7WngoRDEXwceAHVfh4qRI
x+Y6KMc0kLZcI2lYF2yBgILPvu9Q4EiTGZwq/Hyf/OQTyAarXfFZj7K45g8JBeVU
PoAxNDk6XCRrho/0TW1D84D9ka8y94KB6n2kUo66fMRBmGreuAgi9tYQ8XqBWTDc
H9xsrobIRZvuuIY6W/0otuPNtRQHFqvHS6dHnwrY6Si9lODdQSXsypQNqexPa4/U
KLqGoljk01lKabBMcXtnNflDTVolqZvGeYBST3CDS0UdGppVwkv2JWqOyuW94NCI
MJc6XDgCC3JrwhHqTrFnxoGz52Wo+GmVvsqJd/VsPllA5EDg+RdfIQHrwTAgLL5Y
OJSjrM0SueUfd++8WDeOWRGIKLWWMO5anAPk3auwbD3vpc4yldlHlNbf8qRF6/bW
4bSn6HpwOBahJe+biq91ZRfwdLXLu/1l6vHPoMtg6CsCWrw5FW8PUfxHsNThYKOb
UnrOYF6TbG4KQvCYFdNkgq1pGaalo7FwWKDQYS3/AQ5iV2+q3r9c5wqlOkC3TBAo
Dzl+BPugBoNyfGah2BEJr7FiCqfz5BGFY+z8yxV0LBG2Gk/XTXkb5QIuZW6d82WH
K0+kYU5uwwM85oTrDPS5Fl0shlBssMiKu/2w77jDSdcovagzKkujAqEKgoW4Lngo
2ORg/ODquhOk5l5Z13Tl26Qql+rPAKg8maQPYW9XzCzTgUK8Cfo2Id/1saK9I9YX
1KNUfaKvRwS3ffNLfNqPGefe5IjR85SaeziWQCOPPQIjoa3TpUPDLAMggzpzuuri
T4YSTscXbO8FzcfyRjToIy8t/cO5ECOCTgYDtPfhw87Xuh25skt/qHvmEnskELDh
OzbE65XRfbc0SxtkqqJq9Ndix88eRsndlVhMdOMpPATdwesRmyP+3yuM4aEoBoW6
H0DfVkXGimlExvYNcx3657hXhh9J6orRKm48ZD4rnTu3/cP/zSbPMQNLWz960MrA
XG7yBTKekhVadgCthLCI+29QFzcTM3sdVaD/5UJYNcIKrXo3uQkNg0xoJo99bycJ
8SUKV9nYx0g1HqpxbzRCEK/wqNT6Ga2uXv1DrZL35zs4ek44XBFzYyFU9VQTZv1F
ulmnxtKmLvcyksiP5YRTCF1orM7uznAJh/kMAeD7sqJd/H+92Bn4QwDsE97Wpfz0
0+XVyzCNm/HQ0DHmlDQtSn94pTa9h8VfXxnIMOFefu+2zQApBAiGqLncLGAf4AJx
ckYTWWxqTXqxzqiXwK3BH4e1gGqs5XE0ASdiiSL/cXRutGkYnTiM0eqtTZ4LcKUm
2V/zILcpbDerQMChdCT05uDjwXO58874FqAcY9hESJEKn9gH+r6X0o+F7lBuNUQF
ImA88Z+koT4HaOfSDfX3olGYGyDxOwxLG8KoqDYKG1mQJqx7vRVWyY9UKfBFQMkm
LMMgMslJYlPxXzNU0vFj8SxBhNFg2Btayo6O+Ym6NezzI6vHh1fwJf+VyUnhAEda
CFU5BN97H6HwTu01uIsgGD8pi0m8h//Eh6ofUVDjbqK20S/aC7BXz3LeK00/rvg+
o5hTECVk8UgMmFoM2m1qEStg1R9X1HFJXRF/pSV0fdajKuOWUALSJMN/t0UoZXhQ
XJUnGCEnx2lFIAdXiZ97QfTQR5let5mbHKSvCi0AmbNi9xMI2vaQ97L/5jtvuXu1
6AVJ8C9bxbJx0CbyaqqJzZ8+M46eYxnZplr09xBykoiOgDis10ABvUbij+gH3GB2
BwYeKicReKe+xjKsQi9wIMqSzNmpLP9zYlDZJVWmk6kLQGvDOiAfxBeiVpkaoeUK
z0ip5gu0OQ9B7Ols/XE2irg3IzOBIY92T0uMBObZubrsfFoYeB0EiXoIBCO7yWYI
KVNZYqHoF+WdXcTZODn3p8h/oZnmRkwOFCXNkbkixszF2soQs02/Y14L5ipWBe5Z
fD0Obqdk4V8RfDhdJ1JSbebSniEgaIiQukfwUKSr3W3Sg2XsibtW6E+wYbiNU//U
959AorStdKS6NivXTktRCEzxbgmzf9oO0c/YhMOMqo5Brqtwh5lR62auT5MRru/H
1GOWpqqA1P4Oif6XOEOcIGYCHOQeIux6AA80KqFFsfPQjV5xnAOa32K3UR6uluNb
XwJ+KNLKmbQj+AhbNCR4a5kGweT8fE/6nrb/cBsJJbx8+epZSO1+QVTcWqkFL9Y9
CXKEw4+ADeosteTlnDHevwonkCoy+jNxoMId65fMT0fqLOmI9e6dZsqpmguHc4Vl
Q+XPJovw2rfJ+2bMriDKA+376li/rg2f6/FVlPBafV5dacnKsdr8tlFYcuuVbWw0
MNAqn6yrvkzUBvgJeG+IQzV1aIarr9/We8g96yIOyEso9kyG80tRoeyHIQAHvF1a
Do8beDVFzIVVCjzLLr2lQdgfphaFEPB7Hizu+BdyEh3SdeJvUui1Kh0LO4Su/Lg/
Ri2tcDL0LzmY1GR5xQQ/4ZFokkf7KWAdsYSgm0JJDunk8S/VvGC16mGuFQQ38V7Q
dBowEid9a+gnTKaJRF3p+QbO4HsvJOwTHTNryQb1gkIR9sKdLzFPKblPLBkXfbGN
BKVnuBjn/22u5qSYN0xYa3Ueh5DyCwXwS2clRZ3yQV6Yb7Tg/AbIthy+0cfVGg4G
5DEd8WJPwAaMxsngftz4MaGPr4R7RMHcliA+HUSVTQ9OoYX9kZfB1JFsfNRViQ0W
N8gKbmRct1AMl1KHKT5UWE4qYygHwtEsmknXpnLdeqw5nhnzIb8thhsTPB4np7iU
qyDS6ePUK7RM5FnmATDtwtQCdzPPIhg+4cqIaZRx443yITeQpd9C6MM+KZq06YhW
rCgFZxOlzII2l/v67oD7lV/n3q03hXuQ5H8dxtXF5EQRQiAnTiaY+V3gp9opLq0i
uziQLccybdG/AI3iAmtVCnl0VVmQfgbvSecPGVE/2c9WwmDQ8YWqt7fwKCIppRO2
x394zonxQJY+8K/3pTibAb4wAt54DohdKOXtTjNW08rWXSxU+qAi4P2MeECM1hxP
nBQoffsv9Cp3GkLmoYV+moxMLktClRilnHICpwK9G6RvmJF+VZoyNCev4cPbnbUk
nSoJv/zymQd0uZuw4k+EG4iT84sC+JxNwtCvivfSWjVPGmpNqib4/2/5Rh3TprIu
NtFpy3JiTnlQoersJydnfKqWwtK4VcWgDIqBi0UYfrdrsrXxG/akMz2VfdR0pWD9
VN/muAztQzTBc7rlyjHzanpGhCT9a949gDke4KULVm7OZOBp3/vuEYhQFYsAcjnq
Tih+umYERgeOubbisesjRo4LdmcjS6Ca7NO3wqusU/M4OoE9z4JC5OdDyv+5C39Q
MfROSDFkn3zz3YpHKxasx7JXqeES16RdjoaDBZBvD9IwTzMVaYvYtWFIgozgTzjh
ZXo12mXP1fsPq2+j0QbGPp/FsTXn8urL70tAT5MEbhyAwU5OXQqczEsNpkZQvYsu
CvbdUyiMg008744rnzKOOmXKkhS7/Ox+JnGSZuG4B76+Id42xcjNQUhzoQ1qskV/
2IB+O0Up0TgIpxvQIupq8cdMTD8GYW13zgBcDMGnFdu1lRXJHY0L+skgkg84gIHj
CNDcMeiGdbWODZ+5iEFN42dOdHqAh4i+c44EWXwZcDztebpVAj02KuaJ002aRi52
4+SQ5CkKZpLVC3uTtAsKVU1nJ+4q0trSIIJUEHAjm+P0mXk7Tu7a719CISsSUp5E
QN0f6lneIwQNisuPQz8P1c1L3B4gPcZjBRVstI+xArYEDFjFuPZn/eyuyMqgKL33
cme6u8S+kIS60Sm5Qa4Xsc9WzpdQ4SoxS+ElC7R/yphzUez8FOBVW03TEXiQ9Oa1
S/SeZfkWHc61A0DM9ZcX+qF630Z6t2GENqv4PLo+wYdaBhu1BaThF0tP1tzwquTN
KIcFUlOGZ9YomNa5cV1FLDzNw8BCweigIyCDBz9d5uww35Et046BxVHVzTmeuKQ/
40eU+eC7qWoF5Fn3+oVBsgf0ZhR+dAd6VuRkyDBeljHnFVZ6zjwOvmSWsYVKVe4J
2Hdk2R2pjyoyA0PQrUuy3PFFvCgv8MhJjXnBz7oJu8OO1/Z/SS2YwCVKQoKc+bka
khrWY2IMyzyR/YTutnjmtmcbTNGikN4/dQn9AUXbHwVg0/wRjxoNNm+KOrO5C9se
AjTP8x5tjrkxCSdJFgVBa6obK/lTVnkSOsFyZ5e5+Q7JiSNjA7TF8ap/Nh6s2MJC
yetoorq2e4ynhJ5blH7aQ5vIJxDNJH0bH5e2xRkg3r9bPJo2Gv2jjOqEqh+7L2uy
JHKSRV8ZLo1VnejdhlB4jcEMyyEiiQadklrpSTVbTGuOB9Rwt952yEYNVw7zz1fl
c+FJOqGWJxbpyhfbmjuWCuaQ1h70ROnWHwCzcfKUVUhsJWZoh7LCydoGFgWbBLGm
5FPYQqf7B8HXeqEbtCd89BHWvRnEW/xl6S0d+xLEKi7nPlpT4Poe10ahR5PzOKNq
vMDDTGpNOcxrAOivVv22KQkKI8/SC/3y80cfMPw/oG5bSnL5bN+PU5Rz5LcJNe1Q
1TxjS0Aiv/t2WxI8GO2rVHiQ97HMzk0luuMssudZgW6PO2sm3pTIZ29GsCiredXU
2xGQGlZqK2WdUiT75zGOFukkAwfnHRk4sNd1868BJTw/pKWnNVFz0nzvEs3BHYuF
qobliZa8SzFYNPdKzJwiGt+x3vyI8Ua0KbvHl0mpvxlwCWQ2mDG1kYOTTgjyzrIV
9tkdww8qdAEYYROmPXNVqYQF+Y1pgUGX1FXJfm4FWTU4Ruw3Pzq4x9b6Xi9Q6GVd
qtEdCDxS0S8sNgkuu+7evjvEfUw9iRNpEY/RiFkoQVeV7gg6SxrL3VbS4rNhBFXV
tWwvAU5oOC7SVlXqmKt0zCmAwNzuf4qnjRB5TsTM4XL0pfVgoPgQT20t0xOwWOKp
RKBwo2caVGIuKxkBzIjFe7QX7jH6E4aDS6fYDz4NNjhZDzJWEOWpdWiR3KL4raaB
jGdMJcYlt7P58FxicN9CuzvMN49O9Nrn52g4ah+UFmsj2vHVxfaLKqaEls8oNnBv
QeJeNot7tmABqF1Y/1xH55eRfpqaPo5g+DImu+JhRyI4zs2KpaDl7I7/5mfTBAgD
B/yDqYD5S3E+e8kJXcJlgY72aXkh0jmBFOVylTRIFxsfXAf29zA/WtFSv740UqFI
w4BBz7j1nR2iJ92Q4sZailmefDkOcozny8nSOm5WT4q4oYsGg/QvhwCxxcWs2cJE
AKeM1XPcdyW5tgYIk2G5pmi63DES/dSpVOOI0+rfsH0+k4h5R9iYJVFpAVML3uAy
DEL0ANNugS7mSak1STiWLo0nQ+Y6I0ituHsI2RSWLXLqdnhTaql6NakrVj/VThDb
Gi0hQfDVxnG3yBHh5niHYwkCSKo9De3hh//fnI5x81Wqb7bwqJqxXDFxAmfab6po
o/04v7ZCkEItEa8CQpesQiZ1i3J4LxerygvMbMswLecfsMOADCCXgPivoh3+LeQr
9D7vFVCQo6N5zaC8raTAKtjY2Gt+tvE+/Ps7aSZO3WdUt2MgE25mXlthhrF9PeG1
I5K3GQGcc+lWPh1/20xnJ3yz7WebT/xHrBnzGp9/GAoU7Txg+twuHEkMypRe0F4f
Hngw9M6m2MwIYksgJ5+ZECDr4YMymHiyg4aPYlCUjAcQ8G8JG6sq0B47h216r+xJ
aOPgUfrU9ev7WP0gq8rxmC0ikdZna/qQ4qo4Z62JSOwqNZZ/FGSuKus2ySF+kmnC
u/v8vD9IF2oWDfqPH/SNBToG69uIfcbyr0UL8+tnUSMe8CSQk1k0+4gnBHy8e5HP
s6FxxoTcKOQYk29XAvq/4ltVG2BdKQRgS+VzbFl0894Prde5oeLgIy8BX2uTjUa1
8BxBrrQsUoTajFzftv0Q3kGPzWrFcCTIVoN/kT6mb+Hf57yac9Ggzq0FrimTywJW
93nopiINE1YM6jg4/I3sgFExlrsfVOIpUMpTEPfd/BrIUI+zzmj/p1lmIfCsNBET
qWjqnwDnUuibqjThcTcY/msaUgWpT/vgHppX1jQ6Yh+bXfEUjYZCASlvET1B3w+5
/9xF6mlxLFFeigg77TjdyQi/Pq45IpHm3jhErQ17KWPxU7aRG6EkSr2lFdIzB4Z+
gEbjhVlVPA05qXGStir7ruo9GvAdfRz/vjnNT2SiMvBWhb+xPMzv/SNRDC7N0sOg
x7bqtvv9Yx0HEkBKzUVvdSHBVCUUGmtDM3RP2NZJrbiVgZ3FLo9NWA5LP4kHtINA
s6YYoXZYhbFFWPoIJAxJE7n1SlmIC1iTaM/xM9o0PWICDjyj3tJug+dHgXpeTT2e
l5NoEjPvyOX7i+UNOt+8o0J7QtZhlo/zu8QcvYFgoE1anMMRa8uulGU/93xalNMF
S4Cgk8+tJIWZQI7c9I+WyHDAoV2/g+rwnWkf9JSAyEqD/PnTidgoPQsAK6pmGEV9
7o/fEC+BLzgF37peixcAvDVUOgP23B8pS9FBsBI6MoJsrl59Nkb4vOVrfgYcHIc0
a4/f+FcZnLm79zAUqkNySINfwt5LOf5leATdV5uleHpRKo3C4d/a5R0Ex6R8Wqb9
SyJ7qH1TjdR5n/PssBKwPoLj44vanaBjtr5IXrHrQzyTHnxX8wDLhPe/ckr0lrsP
4EsSzIUlqf2FgEzkc1wOi+XJaI0EvvGFTNprqswoQxL7W79TaciyGBiDBAyLIa5y
Rh1pq0aR9crAO0Gq0auX3V2GVvJWtWb1qF9Q5vsURFcoe+Q1v5YZ0KRsQbx3ayIx
p4Bi5Gu79L97j0W5RnxpH7oTRnXfQtX0qMxaxlqdtnP4yYiawKCZn53r5a+l9X+K
GAqMEVL2T35PLa4QTiKQmlhvycOsqW0z4q0JUMijV7RNLTkAv7RxT66GtMHY9X25
aV8YjxxfXZl3GuzPzX3LQSWWPvZnr2DoMrZo5YwNkZ9I/D4hOVU8PQKs37KcfBIo
V90mDF4Ur13gtZ5/z0kIjf313Dbu3Y3uhofEBEut+GS/epYhJ8qYnNHxtADSUo2Z
Pk9HDP2FpCJkIPqfLGOTfSxepj7YM2Al2HlsngPyGUXX1bn+34HJrdmpcDMaGZp/
A5G43CbA3PkB5Ne11yWjsz1LtFC/1ODRkBtTk75XQ3cQcQA8bzx2sZIu9/DykBby
ErHdORgpBC/lmAceZBa+yKirOCYvrmDst21jK8s6go+gBTSuVZnEcpFMMHyN6n+l
msFqW0GrOrkKBA98cy2x+MxWag2KIIgkixVjJPYFCC9iqM3lp3Kq5IK1IpRkxrGO
qCedxYWDDaMv9jEftYn0CtmL6+LQud0JdZVp7Qy6GHWkXn2kdHb7MjHEvpFpeeaH
YL1D6qjychDdv/OtOn806unX/eQQt2TFkCc5PFpgLxqKjQnkwj28gJUIRY8vTPuy
GtmEbU5RJn/6VDak0ySwaWFAE2/+VszfJ43o/+sQbr0to9BI6XUdrEYs7jEbcoTM
qGsbsCZVkm9qr9J8Qx89HJK34LQ/UT7QfJLQS8JP0LzwtRO0U4JHOX+urdPiAD+T
QqxYOPh7rRkkIDEl44hM4CS7TGBFXdceogiRQ6B6EHAC6LS2uZL316Mi0cMmlwY7
ri8CpY5IA8C3uwGP76rKmzir/0w0VK0WU6Occu+FisuCEibYUXKlv1SC3YqZjkDn
uLryXeRyOluHvz6SEfjOYukU1SHARbAq/XrzZNrqp64DXK82lPeW0b1xUduSpkXt
NHmQJLNNVddeYCcbcYAmmxCN5kojhIS+JA3KuDulDKXVAiG6UkPDL9tl8eqUVdxH
Zcga8T3wNcgTI3EgYhtDAFtxiyjFomsXcQGe6xZByHCTEoB8v/Iupefnves6aLO/
HOvBcmQcGknvSvqO7s/A41xUBDT4clEeB/r+DbGj32NSSztr2IVoC5j+QxWcSSRL
OPMKqaQIhZjvEiVFWMXN16VEuV4pqrF0uM1j5BkzVFHThoQe7/fwlZhtB6GBsWxp
c+F9Cf4iwxNKmX+O0Cfs/sY4JxSGS/qZVZmaq32KQRhv4AGtnG/37zfeQEIiroL0
L3kZS4MPUb2L6U6FHJFU3nW9FlgxTA2y4LQnNtuINYF5C7xz7kO6r+xjq31uj1uH
CKM72Z1ZA+mDS+QoI5j+8UpktGt9NkqZVBlKS1grmmrl9izDfKpf3HtLq7TCzLQd
jvyW36774sptJUBr4rlBH01zAJQjcbqDDNp02BjpRhOS09/VAf+9GUJSxhr7T1H3
MsUiGco/GI0akNHW3hSehXfcXXf91OeISYJPESS+0qFeBaTM0jAKiSbQWPV9Vm9b
YNwZSHw++82Tv6v3pU/2YUVXaAJJAPtofAJFa+vFug9h6tWTOTg7XbWG3fTd4zHa
5kqG+xg8gJ5bQADh8g3URLyuVGUprhJjI1GZF47fgItIZNC6uKlBpjDBzyic8wyE
rT5VwpruAlsxsuwgoBxNrdG4odyvQeIFzwatNuJO+bP7PnZK4vDuvu3aWL34D5hm
jenP2A1V1DxZxNNzM0r8X6WyNVj4k0vvLB38h2jw3vJ9Fa5Wz3bA/sDZwAkJ62iD
cTUiIKWj/bTrq5io6hn1Ld1Oa7JMYTequ9as983wtlLiL+ow2RriGQ2ur1iKI2kX
8i4nfAjrFDuSX5Z0TfoCVPic4Kt4XJai7mXhv7H428C7JMkFAteNVJH39nlbaCBY
CJ2n5jvr1F2Wz/YvdOVeSQ0EmD99nWgUhvgWx5OdEJoGm8eGlux1jJmGVWp0Z67R
KzvsgoRqVamsRqFzEJ9GJeViGTucGOpnj+s6MMCeH9y9uxEgK7B4q1p8vGZRHBOh
357CXrsY/zzktBHWc3u91yJsx8vu+DLY/CF7GABnc2Ck7c/naxa0HXtqw6BpM348
uHeDy2zRaR9owCUTFNtFslNcuekwZ06CIjHjQl73D0Bq8eCgLpRiN2tCExfBXcYx
trabUIe8b+7WPtMF3UpACZJ5yxgrIUZ0e36ztmjolnexrh+vmKtwXdw0rDmk5Fb4
DpCxCB2PlDXqMZYUj/Gk7UhS3F53/9GpgiMEACImBdxTZ02wPHE15ltG8xStIAsO
UodJwsBHlAkRAfSYpkv83zjNJQ6VrLaM2yO0ryUfjcbthrZGbvWTHgXOuL7wXbnb
c9DPO6GwXdTy9W1vH30TQNwI3TQkxPSdRb4fsYlrmGNRCn/i+Vej202s0xrHqa7+
JsHLByBPAdI0w8fQedIicd+PxU9R6ekVU7PsJxWmkHuVqQC3QB9/wxnONYQ+lmgQ
8Kmbd1KnPR8ZtEOOuSAVptJFxUfvPtHsQRXNzNkrj2a5h1djDVQxyRFnZm5ZE3FB
rOqCEgLu7MuLGj24NqzLPT0pP1LrajjY+Bbn85kFX8JsMWqbevjXlFxzG+tzncn/
jyeotHOyEnBL2TtL820rW1kF73GNvWs4UBe5d7E1WUuWtXpQ1+3QEa9TcKp8vseR
DAezgMLqWaK4SdBrPGbOmdKs5jxis/Q8BGzztyZK89KMmJoMU5pNr6Xt2/cotzGI
ttS0PlkpkY63Sho2obsiIvN4zsdyIpGlvv9WoKjHX3t7Bl6OeQvxp0PUcoJjeZi5
vE6Zmk30pgd8oeLq77wIeTHjniJJWHoWJ4WepVqL+p3ZvXfbQUxF1cFerqQMLIcz
IEq0jh5E8iVzNh9br8SFn8YD4k05nGb+/OUnhy7Qo3kXgouI+kvoVEXMP1H68ZG/
HCRnPsY2rQPf5RR1+eHLwh0DQmvofUYNn/fUacx0ZN2gA3nkMNR7lKrFpgxXsoL+
ekcxgjojoVrN86ZjMXD1wQTFfimOw9CBI+q4r/CAg5pPm05TTxbkj/k02pi7niJB
1mkLeG7Vn90IS58Wu2urK+etp+O6QF4GmO8XzFCSR/1hHtkKfnESrRMKl8CUCEZc
1BiZeo57mFkQH7CSkfxTKF5I1rzmfqzp+CLNFp8eWS9v/FzUbY9ipeektiOoA7vJ
3z4uFbhjsvg6dCnfAbxD4+9JXfcwotT+RTCfbMQogmHOsVgQs0ajRzRXB36k3UbC
nN+4dja50O1dFAwWcSnp62qSZ03qOOrMAVHnOt82xNaV+QF821fV/6M25IccEXem
H+MPvLDC1JyW5N2OCAaG6jenjMyBYgOWWk47vzDTeiTElrrukZuup7ZbMlD/KpaY
n53KjrGbY0i/M+sEECrt6vvUubi4Cx4RTlt8FADVLuldFWpHi/jmVxW6zO0yetmP
SZK0NlaGC7DhEoJxO6xrFCFjeR4Yv71OQH1dop2gi/PiIrPFLgDO1uw5EMhmQsmX
MqaU9ktMjMwp+f7IY+HrVbk4CjyAYSFRRZtVZXsNTOsuNaHMFDuaeWEhoy8LqFLV
HMg65ltpcFkbxVzaot5hgaEgqRUD0sHzM9GZCYJ9qVjq2PZNL8qfJGVV0wL1Na4t
gKAKdi+slqxS15VrBFBhCdjMrADBfP5nmWDZ374RBp3zalivrOdqXb+lLdYdzvLG
8kbT1+nvGAbPi9zYSa8BjaNEUIP1OnJBJFSblyK21El/luRvEAqOIFsZOf5A4X1b
kP4U1QiuENMChNfsZp54A7sK5xGBDMNN1VzJQupZ/etKD/yWNaOrz9rT8obljQZV
pVCY2t7X8mX6k7kcfOruCxk7K7ZUosDA3NsKxu8CzXpAVOggMYWnUYAlHnt9XFnG
+a/nMJgzdcFe/CE2x4KBkQ+O9oHh7i6XYsgQA6ljdOktjjLt4sdIMlhni8N8new5
FC2aeYqSvcsvJf+LQ6y/UbqPrS2MieNAuSmrDIg3VeEFLSOT2ENRVEzgulU04X98
wY4lwLo2KVfc9aIR5f6V3xfaxqKRdtK9uFKnCErFnj/wbR4beaO7wT9oHjpqF3tt
2/4lhi8uGQKk/W9T9xJCAE2PSdNzBuA5k8FIex3akgMqbSnHm+58n/Oh9Y8Y4tao
MMvTmhig4usYiOC7A0J6YiO/62ykxDS/ripIlfjUwMJwkq9KPFQD8UiBFKvy0Gvp
caZzSjfn2Z+BcI3u70WI69bwJzQs6bNbtANwfAmaDFC6bluSHp2HO6d6Oh6vedFA
p/G1G9ihFiPsPwDIVVhaL7HPIxF5K1w0qC1xAFd4a9Q3Zj/2nx+JKbjkCcVqm8+i
vmDG3CPGoEsfVGUtWydM4DL+qM5AKB1sZOweAwj9V6yVnXOjkDdTh+rX0Ja9OOJc
JqwQx++ctGHPnRgjJmzKL2KLfNSNrZsmkAwoQavmGG2zcfSmvKAFWC0og9QW82Zw
3J8shrVrk/E5Mx8yqs7FePiwnoC7i2pV0Km2F4oOs49BwKOmEWGqqOH+DpBZldaT
34d+WYJ+39IFxZXTLzv5pXhVxnJVVvXE2h4hT0sxs/udtJNbnhHjcsS3jd3ATEGx
wA7NTfbfh2DAKudWuxwyWMTMpaYToRXigHG3lhyMeCJ5Uaq1hTNRrt9GnG32yNRL
P7QBEy5yobWtwlyrKYePX+UvNw467kfRoH4v7qvbSQ0r5BZROpqqTCMXRm9rXcqF
Z86k/vZ8ddx/xvO2zjpVEg9xPCyvqxgnKZDtdsI8EZZzvD78VQms65pFjr5TujiW
dPJcYXNcH8EicmuhIgyenFtnFwz2DdAcOOKzK3uSZCZje4fCzKoUO/VJAzc1SfcH
Vz9RU62Jr6CWULjZ0fBDRQbTgU5dvAWT04OWTOtIJzurZx9RahPDmic49/mM/Re7
cO/3P+Y73qIBaoTCj7Bnx0JCRUoOldEPMCIsUQXfjAO/7DarDxxaajByTDYy6nFg
4UFw9+uaii9X92Y4NRZBJqPyHQHOHod+d08DJm0vys2/2R9WJtLcrFGfIIkh9Nsl
d9Vf/KH9TjumCyLF3J3nvQ1j1EWBw1te4q66heFFd8Dzp7JDfWNWXclIPZ9Td8TE
Yi4n42ViK8lKMp4RTuUQkr90LZnPVzqxrtRaqQ3tT7nSBtayy8ZcaZGWjie64p67
2MoVyzQUxTAtTSWMEjD+1U+cB4WUH96lV/RBiaQpIu1Re/+noDlN/4wnj4rdl5JY
nQ08zdFib6aBYh+J67OrYbsaM6td1U3Fq+8xpxQqhS0MgvEnPQ80Z35zikbXPhFP
Z/bFVLyNCEbwU6CGElaiibfkDnibdOEQYpmEKoECsNmRQK7qgvwk43MDNI1yBon8
3C0YcN1C/sGxrVrheZYiamfv+suJDAMdANyGjnsC03GGeyFpHh7D+82XqYin4wiV
yym8Vn0708RdCDKxdi/oi0Q1SFHQaF27HG2KF20tn/Th+MxzFzaFIaYjc2+WF6YN
qfpDLCQDPF4vLMi5BJR9qBBRAyQM65EKcSBOkK+MSosL/6FzamiWmLh5qk6S0xs0
j9hrukncAC7XuoQmVnvWrzcE4hr767CkzYOhmn9jnoGfzYDCnb0X7oeR6ml1P3oE
2/d/KqgX6WYRHpiY4yEi7ebTEeinAEpavNd1jG5nhYeZuRg45SpoDuO/qusIyoh7
lsESATPt4hmGewQqQfwPq1hlm3+rHi8otfOLPNee171eOK2KjhxpS9aEI60FGvTE
24rLt5mJK+eU/R7Sk0Je8o/WvqqqTuWASWDfZ/1/t4B+jeX7LTgdpY3LBbVUQHZk
0hH2GMDu1D7CXigHxtAReFWBjUYYqZ2YgUW5qCGU7qPQaMpDMQvh15dZCaRdSj9U
eYf2LHL2biS7dnl4ePNHd8gFJ37tPf9FRX4oMBI+5tWOHVzgbS/zF9kfqtbFl4oA
EYKfFZ4vYP6c96SA/SUadkaAWUum9FhMWhLzbfwI6pmEo9FGvs94KdmNn8StoQLw
R0ekOJANPOqvjKwDCZtgwa/6w3HNKcwx5qOOr9Uw+C0UhIokKiynFg95I1H6nM8s
KeTWCIC7ekwdGzA1qmYvKMGxp9OkC1DsGEpPtcCv3m4PxbzCH2qaZflwyOZFsoZ4
ZMNxQMoWSkBc9Hiu7bSls7D389vN8HIA+8P3VguGfxsoWfX++4s8mBUU3cjs2gSN
vBn3RrWrfmqUOpdU68pQezyl8urnKL56DpOduwqX+D9wJgszDTndj8h8DpTWHKAC
fcofbMR0s6YcRalH8cSKoG2PtwYNOUuyaaYDw5Ebw61rh9LHPnW/lb+AqF2sWtC3
F2OpntrV4nW+YQQA8zuo4xaF/lqMoEGIRb/mBsuNiDlwJF94jjPlJckdURFTcVGJ
uJNUUIbBDxAden9PPncHxermExb63oabhhp9uEuDJJTiUQnA6WNtk0C2yFMRmTyI
BWwOwoFPyFnxg8kH/0ckr6tRfXZN3KXJ4VU1XCJL2vSYjfMFXbmoAFOyrKathht0
asv92Af4UVcmiWWC7jNuT2KorTgSdFRlZ+GnINJsGgDCBzjZN7si4AB8GY3ovQX5
lHoW2h3SU51fA3vvUCIyztucNuYYpyMupLRrj8+L/6QoSt0gnsGifoAXSlkHWkL+
+PEc9QyJw5Lx7P5PJh+upc/wHNhDTxbryl21GRW3uNIDP2+AhvZdiJnvsUFvWyMM
7BhTen+21A/3+scK2nP9uf8t0bQRZUl9iizdKCWlmvYwLs/pF1/ndI/BWYRQazjU
As/Yqa3NzhbZat4zlmfWfR9ZfmZVC1qL/MDnv9tlu9OcMqBdSKn80tzsmXA4yuLn
Alei6T5NLwxPHJM6M0zOrZwVg0pq7U0VYOSuC++dTwXZMrhsN4uVM/5hPfMKoOG9
03qOX527GaxXSQhFCqoz10TSd/P/WhZ16Kjf0rf5iaxgbt1GWBcmJ9+zrQgUt/WI
FEQd+xwb6PLKyZjwVpXHgaD5e98Pd2xozMBiq+HFv1Uy3xTokYVJ/e4QBxBN2jlg
7adF6tJJtnykYu2aMWW0Fz5HFtW9OvJCD9+hlPyUJ0JedA6ecDeSpWO0QK7Nqozt
uMxskdVvpe8Aasf78k4Y8+hGwHjSDhrh+F1iou/msfxnmhlYibl6E4bwX8CmPO5o
BvPxAkbUG1GyZX0ku0UUJjX/L7bI/wQA4cFMnQ81MZgq7On8eT23ABRG6qd/Wq8+
e3C4yrNr5lCYJmwSMwCIC3viuGtQXWwR6NJFG8EIkEg8QDuCdnIeTdweP/6kejtA
5JKK6CgYBb20b0eJMvzp/+IdgogRoWJe2tJWzBnxuyWjNgWXkUuPu5mPrKWm9fiE
F81I8/DU3zEGvGKoVWvSY0wvXUgDVMRnINWyfjSzM7JsipkH2qgdqdCNziTTSEXC
8tgNXCUm4BFc3VJJ9RYbnRBHJPo1PgXHoj7UDcx3Bj8rLriTbGMBJfLnMiscUU/E
vXnf1dvtbRenUXa0k/suzj7th/+2ez7cGJNngYyzOdWx3nMJ+w4JW2NDvuABCosR
l48THd/GQrhSvqygG440M5H2BcqryQ1ZwGiU0ZCS+hMuKMi9qAb/4xjfF4FV5rdj
zeysAqg5SlUKQYF/ndlywE9eh+sjzaNFutFaqk8ekF3BJnI7e8jZqQCgLgBJBVLA
d2pm+qDtt6tO/eEe8wT9Kk4lv/mV8SWLjxOwMXH+3J8rx1Odi2rNfZ1pmaZlh62S
gm+kKwMJ2oafLxLHokW4YQlnS6gGagd3WveS+SgHmep+4XYaAbW6N1LpH7EXfahK
ENPo2kHMrjelSnu5rn7MljyTNrXjL9MdWFLKZEyDKIGwpTpvRtYyy3dXpwR9FgiO
gklayYdL67nUC+OU9P7A50g0GErU/Nj2DCMnZiqFvKxraU1914RakQLp/79awmYn
7n+t9W141NM9TZlMK49bylYIxqpPqM7aquhYLXtxT6nlZs98msgnAphQcdSx3844
YS0wIQtdMSIJlWC7F6prXq1wrpiEuV76lNxo/rKBY0qkQZ/eeHa7r2n9am5yiLnN
52SnI3Ua89k1L6DKrVXJCRxpP9PGVY3NrpMxdCxJyB16zX1PfkA6filZoziTdsJp
skSXsrByLK8pSWQstKfpM+QlFyCZ246dZqCJ/lZ8sOfbIZtZ2j7M2cMsHXV7Cl9J
Nryjjp7H9mYbBz+cCQoN2HBvMmX6tVPgdZdFBRnFw5lN2SK69omB/BFeZO86OZG+
7ravUtvjxXzmZLUvLugX+wd02y47hyNZ7JUVdgYp4hIyJ0G+4SiXkkb05WUi93AW
hZscvXnJtuF2DbNedjJFpv9HhTHBCvPD/UUH4fTCA+Msys+APrFMcqiL+AmizT9H
MyjOwhpZkgp4Bz+xly4ZbsiEkwnW/kxQz/hFiDzJgrTUo56RYiaTYe+f5vIxkmfF
TiWsj1ae1bc25tZtP/mLxQw1O/Dqrl8N9wZ+Lz9xueztZXyuTGp6Mh7ohyq3oMMI
I3q6xpHFf4mdyxklbpH43hCR16D6VUat7ZT/dbqysD3jSTdoj8IZkEvXvIH1D88i
rtP3j6dqsn0gIfCs19LZE3+4d4hSXamdZpz3fAXgry8e+jZkxjebfv+pAOXHCoqI
FDMcv9oCAGh1RQ3RC/vWrdOF+L2EMyPP/Vh++Dg3zrn9EdX7e/ia22ovkk4xZh9M
BCe1ooRep+xmyq2jR1RlDffwfYyMxRP7saLROdSI2H0wC4qjvXTIf/gYVhYveKqf
Po/Ol6rJbSEO6r3AVCHKnlaSMXoVpiK5IJMKCet00qeWEksKz8uEm6blC8ivUeX8
s3WUBEjV8xexHXcvNZ27IkMNtHGHMy2LhxFLncjF7I2tJLau5jZkZGAyn6TjPYjr
BXVRjXuqKaDUGxzrj29qQBnfCjyLUkDxW23kiO/LV7tumP7gVb3sX62BQRoTjYej
AERoCsZLgPy5M2cw57/bHfwZN1EIAAuQqLWcHE3sdoobbncQbO5+f4XCerDqDRvC
fKCzJnJbs80vka4n7qSvWpDbEak+di9XfEA++t/AH6bnT30tErsWuEsnfzKEXMfm
vKkoR91kvUtHIJdXeIqEiT8ph0+7OTEkVmFXyd50FFgIL0A1t0zLgMPZpu3AaVEJ
X4NizUqO5QH0HQqyZoeQzA5216wQz/bbiCBombR+fp53io1/dVNZMt+dKahl76jM
hW0FOH9iyr7rUxKeuyxTtTXrq2vnFkhQcD94aD8swejw1q3dtYQCx4FiayZr9BqI
1B8On7Kx5OBiFYWRnIp4LgiMvCK5rNa7JjR8FLyS34py5tuFfD5kwOSBI99NpcPJ
U01k7mGy27MLst5rWO+h+LBd2S+IR3klB66yyvpPG7hUhEIM6jEx5N9icUtSix8t
wixSaMQfzGZjsNoiUMy9zZv0Ho2u1LP6QoLaBszNAr63smaux1lLLWDcuCRNwDb/
Bj+0Vv6K0dXWnOQT/Kd4OzGJccWylxu1EPxM/RyuZ3smJ4I+rjgPqoukAldW0dbg
6WwPjUO5agxUm1TLCBLRYWcEPSZshvGK56Kapku1vkikF870QCD68iSUAy++1v4J
QiUqKz1RWELKzLNaS0oQSxSrZzY7bwgc5v1hKt7A4hnjgF7wQjZ65xU7lSRo47II
IwOZe5c4YzuI55gRZ4x4p4WLnwaQKmMiJ8LOXq8A88+zQrcTpxM8nc9VeFcHRL7U
vqHX1GlkZUiZKNakTokRy1GfWqnifbMZOga7hofq6tNEnVfgwG07Z/JYpRpLi2TD
FjdNIPtxx9LhivNshzbiZ7WGbBRXOytaS3UykduiRyXD+ctx1OKHyifqtPt3HMRx
rkMqc3V4odkO5LRW9TKFjLtyCSRwn0O6YfdPuJe8QSF43rPOdjR9E/0Zahd5HHWN
2Wi8OXGn0h23TetXZxWwYzkrRC0Q5a34i7KTrlM+ueF/4e8YOtIKJ6z6G1xfuPxx
ZEVdN4OJuzj5D9kNog4OK7I74vnmfjEigoHl9Ebb+iV+Cn6J9Nw5u0sqwoyB68J2
maTFR8BynY9XYxXmgUf8PkgbdTmYA7qzeP41UeLXtMWmWB6foBhqX8TnKMsMDJiS
IyfkJSMXDt512eZAdBhByHKXVY9FM7AU/lW/ZQDqCJll0X8+6bIv5e5xt5iqdu1v
LvnY56Eizs0gXwFGy7No5+f3lhQdnEvELIOsL8Mou+Hs1nesXi9WCAWnNl6VW00h
sI20mlBdTQS7Gg9oIofVjPgLxjK5xk5JpVAbfQ8DPqtVRLq2yR5+yos+KFcUDtTx
Vozlpwf2MRXFCCX4+FMeXqu8XJIaJroUVQd6eP09Px6wU4CcStmIUHksJqum1u8w
UE0JBt6TAv0hTY8Ah1mX14CFBABJHD+xuEbfhx7IOhqf83Wd4K3NIKdapInvrjqD
llPdIVjjzMroiZh8ISy1nkDMCVSuSbK6PhvSqh47V7R2o7x8scMiX8JMIM36Oy1C
LJoJgmKRZotku4cZgU/9Bk0etdSJnRal2ji1fRDmB1wi8f2KA5nr2Nr7KcGPzp38
7rj6vtDHllQ18Z0i+GVgX/ShchFw82CX0OCccAWhAZkXIMQ/9pkb1A0d+EOv7zWR
KrlfV/RDZvQGMZMwEvHnh6HPuLVaIEqHEEpoNfR0ZUG1cwp23zLdDjMHjcTpjsFg
1NWuflY3ZZiSYfrQZ1tp7iN33GQOZqeERb+DjhV185RaFxBH2EqMl6jW+q305NGS
Y+ysupP+UiLSNrcTw+8xCPwqi2D/8GOrrUseNzC4TicBoQfy7GFcSoEREsuhTmxa
b0qVx+6tbhnqqH191xQsF6C/My925xW5XBHWkQ9s6IkKGLqV56/+WeWoSgY+nd/b
lxE7u6SSp68FFmHxw2N7mD1Bz6rIfABSP5UEjsoqVf3YryRgtZNXX4ovlsBvrKuh
6aFsJ7IIZRzz73iQDdbT/GQpbTYNdtpTkXXrOpa454I/h2zQSunkiBmfcPYmMhw9
tXUPFITKhsaJU1I/HvV4eZCRN18hS5sMeeK7KDvSgkYLTef6PWS1l0s5I6boQlWK
U1qyegiqOnHUn2ohj6rlKcFq1ryjXLaFoIN450YnfVr18wQtYJwBDBf080eThBKM
I3SPPrRjxQ1cDtOj25XLeh9mpiXBuEl/ax4/mcpCEdMmpkM77iYY04V9/FOHz7wD
wA2SM5U1bHkmKrdJ3+oi/Aj3xluFy/1WLf3mzHUeHZJd/fZKQgKb3FagurVGMrah
NiIjvQN9culJLj/VFzyi+ely7EjeR/myXv/ADRB3kQM9drwu5tZOEexsfaGCq+zG
DJRaDMc1Pawrbb1ImS0dY4mHz0aWHtf3YVOZQBUwRTA5uVcBW/QhVTm026TG+bdX
NlAekIBPkfjnM44sbJvjhwUMDTir/NZnQOsHetajayjLDaNKWxc+hrvehdJQ9KhE
WPM4LBGUIymheX2+DTAszOTqa9FOsKZo71Ve+Xq8mG4Ar+RgV8tkeMZs4cNH6azk
PZKyKb3xTka/X+buAeorvsVYYKftfK3L5r4pAcucS2E0A9SXdA+Z6CFD3BRGLChr
4D2pKYPfO+UMnp1YmLS0pKmhFCcTAKPPfnqqjKExbjdXMLX154COuY+CBwjh/rXB
G/jaIbPQp72LWkQdK8N1JWY4+uVu5XCEVeE80Ojeb3BX/+cJ6kMFofdQd8uzGoXi
TrBWoOaxxGtynDwwii3tKAOOSlFokzvYW5V24coCmMq0BQezjZxRlGIoH5fEOA9f
KUzIkhkHepLPP8ZKx93UNjIZE2bLyoo0JdTU5ZVZ1YBPz4NhCzJLNY8C+7URv08x
KyCJRKNpCtwJkCdnHBSSP0udp8/MaC7E1sibj8eD7zMbeNXsTvKOpDfKwoveX5nM
31bYoEiGl/Ru7qghxYuLeXKWthoKnmB1wO0/CZ9UR11aJq/5HKbGiEeF82TxEk22
TFF7DSrhlXnfzKhzXn4uvsekpZeqQ8BIh/qLLRKUJPbKPKKy4fSChQ7eCNDRqefQ
wUk+5mAT+9dzpDD3TpfqlTogLwhD6rKdpQRTAqq/aDUEKLuqYv3mLOfh2m8+iS0O
vNWGtFbn3En1wyzLY7LVXo5JiicTlh5GkgdRPv7SE7F2Q5xVHz77zchWw+HDEFjE
I0qilrflYjmZrgOtWzCT3MBBZ5jGy/E/ZRP8Db9gIK1bGf0Z2HtAZ51ZalHjJqss
yaOcPzKCUCjkFetmhJitAbyM67kdAOXyTPrAfFkUDoS4A2OJOPiw6LnoBR9Whogm
w5wUTDRWlec2Q6BB9gvfklXuuKYVq6ITfIerSxAMnGnEr7fJS53YHRKxLSYx4ala
g8E/F3iLTCj3ytOo4rzprqExeag/5nk0c+4QUziehG/PCAuQsC024BWenUQLD9hG
dwuMXmbwBYt/jCv6nJ8psGN/hEglk0e94zwVJ7wg0xEQNl/VdFpnu4uV3qv1Sxih
4Ihe3hKG3hEI7bRBEl7/GZNH95ScVCzhcEorAZgtfj1H9bOFs9lLn4go/vIlbQ55
K+ZirP9l089XgQNMKyvDeSFp5pr7Plpf3/EYt6iurGOGITyObUzDDXbPmL4xRQtM
b02j7RNwYmcxiU5NkByYOgIjSeFXtuXYZ87z1Ayo8ez/Xdu2S8QU6huQhG6rqr+P
QyBWGdKqcayyTRwVdNelTb1lrr36PrUCQ95IAiGNVwkR17R5WkxX6nSRrwMS76dI
DTbn+GPuf4lXHupleR2bEVLIk5VhZ+fcrLVV/rZKyIKl0tdZPgjUf2Vsyq8opNe4
ECnwO76gXp1hx7kl/XmpUf73VYFdLF8OetuyTmcrBWysCCfyMVQAzowir8yNNC8r
rB4C+T7foSZb0LD8LfrkRyv1UISan16yT7EVbWL2bip/opJ7gto40q/JczxUZHsf
fI0xg0Qn9+SWcSfqoYP8hG6MPCA0JcEcT5rKd23OrdjMc0p7fIKuexdw9jFK8lf1
Vfts70qGEE8N4kK1kbMRSqQT+l6agJe/kA6duo5UuBtQzd4T6j+SNjmUdq+hXl01
xCXvoK57lINxRQW7nL1uu1+qeW/GgM8BELtYs9S+UJOXHGaMz8glhjwuVFBtJ49D
FtnbEPAzJrxzTqACTmsqOJaOOIuyGkIke/aFTzujhYi7Ysk92g6ZvMSGxenpJHtd
5bMuLUSpjAPpIelQW3vUZdSWa3HI9+V+GZskwiH3ulIBisJ+/YqHFPxjfml9MesO
kuBFLUvO+IYwiwh+eDvbSzNXVfm6oZZGRif7Iqcdtm94c1VbvXyyX4tVNmWrdnLA
KprB+xxs09uIjk5ej3UJ4Ypxg4Cjjm072zViq3bGQWGMPaLRdroV0zhhrTmK3cU0
/mlMe/Y+lTZ0MKGlSHC4hsxUDPCGr8+LP69BHWCL0Fbn+PoUfs+PngTLSX0GaFZL
Ia7yC0QAc3eX6YHwTj1u8LdS1G+pTFq0hsdPQRo5tccHBkgbQ39iwBxUB83kohTx
BZ7LE1TA2gysfVOwExqfmoVF332tFXRuqI/IJF/3deuztUluY6NLE4zh/jjE6/M9
7j+yIX+QB10OFIuzhV2kE+wcL/6X52Ysx8nU8xTN0V8T86JcsKHB/pKKd+mRW6mN
TAXgZFiYFFbAnl0OA0ZJ2t0ZO6SjUbPC4uaXAhdqYKdsysm09gwN9VV9fxL0xaer
tupVStSy9p6QSZO7VgVjUXNma4mwJ5xpa28s58QQ5U+daaWBme1m9SYsciHlf+C/
2ICkoUNKF4Yiw1O715oFrpPwCXySA8YDQM5MopmsjorZuEZy/sF4bMT8KYYRdKqq
jVjTZvSVWZw58kd6BLVIi4lMZWb+rcKx1q5ZzHMKNvOcykigKkUfBulNRCgYcptp
D811qFqlPJW1/wVgLUAM157faWDr3GqvSue2zQ2i3TZgDfu/W5wjX4AGg5hbnjQP
A1rdfbPG2tBZGnJM6OjP1oOTQHcuIVQ1EysF37utVXtJ3OY1eOpnuSnNzHxenQnL
V4m0K7EY6j10YtcTA3w/gNIEUvS/u0pvMzgf0jR1SaIlqvfiLoehM3/TIwlAO6dS
vOcant6FoFQXZWYUr9JgMvC9LAUdNfqutg4io2+mgR1ICf+UEUW4Q+KugsauEnZD
aRsQ0Dz28Ri5J/Bu9re7z2DmFfxF36k6qHJS4LyYTxRKMu6wsHIH9NbJUs2/JLBL
Z+AUf5arAeAVmoeB9ZkhqsUEH3jC6sXBLrvwsb4nMfm0TaqBIO87dq+rWb9+7Wpk
fCHR/EL/ldU3piHNsSxfCOeG2hKtUmxGdtAUHspCMS2RM0Qdjumyi71rbTJpd/aT
Nqr+ca8ppL7KTpIQt/7SWReGj+wE6DoOpRmShsW/91ZN380YJzOZUf5zOtDJKE7Z
bOrMPBHx17cMBA+yNWZC1B/PNULeAY+jC6J8Ha6DCScPAd4ddEk0NXIwlg/PwiPm
H2gL1l1HddobZTIJ73kBJeiTRt+CYtiIOkPBXqQxHfOzjzjYUSzBX5f8PCtcXsw5
ZimbeZTIISoHn5Tcs+iFz0Hl5F2DAHD7wqTUDthpv4somgkzAcfkERAXWTwZv+wn
rnld+bhVFmaapq0+65yx39nxbws3kPpPzRt9PWf4rD8WppgcBjNVGaDEjUfTxM6C
24PbnGuacKPvg3IjxV0up8qpO3hL7K2gukfnJv81kztmHA7V/1COdvcrh+uzeLOc
iEWDbrVfjUyIcVUsiAG5P5VUxk0N/DnyLCV5wSqalxKZcQtIK2IgbQmKAimumNuM
Eru9g2o1GPvtWr3623CCvNhxvVjbkEAYm8NBJCUNUjL8D1Ykb5ApSss9coN/Bdiz
64b2ZxKaEucEBUBLE6KTgsI5GCxUhWiywEEiMC883O3WO2iCzA4U3Tax0TDvm6am
Zbjl+gYN12XoUM4jFgUwi4TlcaVtfwPEuwAJ1qgdE5qbW/qWtU9NyE/bc2vc39FB
qAmgFsnOUTvEsuMxSjwbroFNk0wemVdksGcpb3bGzrelTWiRyUFIPRyKxDvK3ISk
DLOWbpeKe8BjX1rYKlisU65h/NNsM0XFuGah72qz26bRX7Ltso/46KGzZpdXHh69
8mDgw5c847iblqL2rOPVyqHcHDWHl9NgeyYPugQmHIaHdhKrcZ7WxEEiHrbTDlqT
noRM5guwSuVsHmtum6Od/Xh5dT9yHgpjNXPZAP9FwTadtIR1WpSswWzxJvtNQaDE
vmYrYVXYgVUR4MjUjlqt8xhw3zRshtMb48AVloeiEMyq3dX61EqsMykdmFG8y+PL
DoqIfy4fXmB54UPbZf4lY4DSmM7IqllVa9PCnshKh0u9q+nbED855f//O904VuaK
zjLecA756Ol4qECnlhCzfEI63WNvXlyEpAROYFJ+HDZFnp8Y4jOCQQhLFeKv/HHl
QbZfnJeWYeOR+JKQtfJ/5KI6zoa4y3g9LDxQzOFUtIkcuQiJgWQ90R+WocBWA8WJ
lEU37TYXc+AB4bbdjugwzYyxYbmlV2ZuZT8CauQlBjdA2+lyDGdVMRfgQP5LTz1d
NNPKBzNRtS4VpQrjC/yIP4aj+wysumPBFFnA+ItOiESEvSsgj9wWmdjcrgMMFSqv
fPNJYuRk293DWq73D9dn4wyRK8E1k0wnouFxSRE7fp9rjk6ZWu5gpxi5MWo5NpTG
ubZrq1UYMH5Ll2GNsXwgKVlJaAq89ODulkLPwrG4sImfpggzJ4A32E4ERcioRhYC
qvMgQvl7CUeWdMeq3M7ccs5++Sthcoch9Ocx6XVe+32aIfiD2/i/Vpa8qF5MTILN
HIaaF67UqCF7s6wEdyKSiNPWuhv0WS2+vXUcafZIDfNNQHgnkCosKzr3lAHQOJbd
BocAemTcazvtix/bgBUX9jho5OtlAWfLcPAg5GMSaV9xBq8N7P042W9w007NanWf
LcxyPX0AXA1Q+Gq8S5gnMMhvND2hbr8/mJw+9ZiHBwAqY/vcSLuNrLVldALg/DqC
xGggmroVHGWlYoUauXY5DbbJ684LRdkgqmm55xgDakELj3SaSRsdzbaLDH1H/RjK
WaN8g2P6OMc5JVhYaGyk0rKDG975V9qt55EVkm7SrJhRMC9ZkJXTefFUUd4Yt9sE
9NEad51VcJd8/BBlng7HOoYfKP8O0zvvX9cPM6IdWCBLzggZSoF7gQV+/GAr6VlG
p7n8wMzygPN3eiNZ5m3FllBx6NFwFyiYYB3MzKe3bQoHXpM+nCW27HzO3I21N56f
BUNwc5ZyRZh+0EWMvS5yUGukqKgG/zMvA9SZ3/hIHhHyZie5yQltWNMlc5ZLwcrF
qR0V2zuEZe4Dn2DMls3jIcc8bWvTL+PBExDl6PR2vn9qKBuej+t2JXul3N+L3eoT
eLU8V4iPumLOrqUpebLk7upqsBtxxBPN11iXVBKneLia8D55BipoXm5AaEAWykvR
xiG3yfZjPZzt0aI1yoHcYD6HxKCN4F9rq4ymRrCemPj8xuRgvBD6+u93FwWSpDt9
GfFBb33n5gUMHzirelbHqX+V0NrRMuYfc6YgXq39aDBqhvlktUxaEFKmlHWKt0eq
2Worize7geeEx+GSW3SH0BKK7XnQjSAFFyhUHTNmXywRDEquRnVcIhZle/HfsGxs
nRIUUKDmRr0/3PIV0u6cL7CPyKJ4xWLvgYiEGp8hhFzikXddlrqe6fMwaOnheZ5f
QQqKTO/5hvcsAcnJw+Y07xQnjWJe5PqQT3w4DQ+O6H9+B5tupi0wN4HvacimQgop
Qx0YsnS1h5KTFtZ1PZ5Cwv/qnkOvabbURtQNqpqxOHajK0kfxroCK1bSdcm3gMKa
zUeSdt90W3MvnqtafrK3IwCXENjbZPwPaCLlGNiQC4Zf1H2E1BKQVvePcUaCv86/
bGoqmAUuNIoHjErUvice8g+6XMXgJbIVkgzQXsKfabqTZJmvu6YnrcEHN/55KIRF
s4WHCVeLNBYyOPM+BdyGpJXaAYeoDPFOX898i2+8yEJwG+y60kzzyAAJVIrWXxJ3
d7bf8xmoCIqjl5QwBsxQGrhejGS/3oyLZ+Ll1SuIiwzbOqEJYS26LlorLKC31zMO
0j4A5pBq5zO24+AknZT6ux8eKJxxepCSPPXtBNAQMx2sjUGMlKuWaKErI4+CakMv
FlEpkxurAxr94QFU8VinJtHi7Wg5TwTgYH63ep8TWdX0qA+Awzjd+F2wahwseHn5
rOPSumf7tokP0MbvHofhr+pgG+2L9fO9SnBuDBmdcT1qUQ3AAxhDqIdOKkiKTWzZ
plDu/MFzajBGuruT9rLIdQx6irUs2JZ7FCWCOA7rk0DtibvKKJQ5i+CKz44+ZIRS
Hrd0NnJI2OwdmpnESXKXIOcKNjCceBMSTSDIRj60Oe58NTYyrwzPtwhXP/VjhVM0
4Jt55/n+AfNOlPhf4y2zkSRNmv5TOjjC8nL0kmTdyc69lCT7nZAALtYM8P+ZR4Xq
43rsPkW6g/xxn89Jnm1l2lkB/kt2LcMdLeYu4s2AADn932yPNHu9pC65hZ96mVhZ
uTVc8vzB0MVIqXvUVx5T7pAtDZ6e58jPF1+5MpiDzjlGS9TTcsEn/fvsBQt2HaDY
wg2iCi3yAOnYPP/zPqmcRhXPXS/dhd5+zs5bBR+7u903rz22jTt/irCNpyjYEAhY
SB7U9HisEKGH1HbyaLlD1oFImRvyC6gv/eIMN1GKYFGmaBSTJGDxZ3+3RKsxlNuJ
kO9fTEtfR36hs3z98nAgl5AUhy4G+yjLd04FRH9xVSKqcRwKU/brj3QqxPDR5cSl
CLcAXlapndKpVguQ3YumwjbD/KMldgX1+jY8xrtaALxYLchTjoiTPaWlkREEosN+
3iyKSSteXV1zrjOpUnRvpefikVDLWbitXFD9peXfl59myeX0Tv+YVf5YUqn/hrFm
cgATKKXc4BW8Qtos1J5Ti367Oi8w8YNAIoyuXTpLHkuBtJVGs2O8w2FfCXlxFYh0
gA34ITpzv3eMQKfuhLnwAzHdv27kBoc6uozNIM7izbLRQmeEz+bSBdYN8mfAPBpz
e7VW6DbmWIwz2/+fOf8k4x6QL50FinI5y2jSB+j2Q8RdbYyAj1hvMz7xjwC1q/+Y
w+pEaWty3ztxLhSJZQpjIQA197sfeNxKIrCf8R++brYiHOEfFWJ4RtklbkO/p1Q5
6x54xXUXeUfZi3r5XOUl5J2lSkT82soZdNQMmkQcKaRm15rHXBAFlZMjIR81+RpV
jCtv8eI1im/zyPbXySlgbAiyp092CQmvyemrZVWyaVkhUN8+0Zvv0Cpi8ZxS0ubP
dqUVpzp0nbFyjzSFWzZPva55GX7yY/B+7Wmn5U5nrUETEX7ySQm0u8CUSV1rPack
hGM7MChsvk4UforJwmL59bS2vsW4faLSNaf8ApnhO4j44hwviEVVfh38YdjR08Yz
Jt7+VxDi5AExToH5JtcjdRsQFy3CgyfLljkayfVcPY+2bJEdNbqFb90TxfTzeEya
O37DpnEJWbmHgP+KT4Bv1QLWcSz8+T5oun3o+qmyRuGnES5YXUwNYIgjDjN4SkK6
K5WNn5PWYdlqSg2YBBKWh6Yq3vfyWD2P821RUoaDVj0cAmRzIB+PwvtANWL4MamV
zMZJJHLl997aTSbLMOziG2O5TtQq91Fik/ckJbtZvJUPYUJpUslAppXCS4ZYlgRN
7V13qyBot9lgtQ0d96xbUq3Slv+G60cQkYDz4rhiZalLpkUbv7QFb6o+pyq40DC8
+lYkhIVW9feeEjBRkevx8OjzB1cV8SrvBJiUKEUux7/UOOCymgnGZhazpyzmSVfo
gEvJeK2F2DZxe6gRb/b9w+lIYG1yH1x86Z2jO3ajAVe/1p3zSrk81M3eojyN6h8G
TVGGZQUmu0ymfjxdqubItsi2XGgPrft1/xxRZW4kwjvgeeXYkD1DvuZ0GU06nITq
mh92chtSoLAraQWvU+ivoZdhNta+SDf3KLUNdecsoZgF+kh1XH8JSueng9n8IA0Y
TfljMS/tr25g4bbWq1RpzGuH991CBgjVUWbTGAhZXFnjD9BY2YFl9sHmaWfByxYz
TacMdjHhKil741GNB/sv0xXCXa3xHbGHMB7aIOfNzffS2mRAIvDY/y5bI+Vc3MOL
oLPssDZY8jr440WUO7idhYSbEfJwMJ0SP2wlNdxU6tAEj6sDXg8wxfiBq+/PDZQL
imyvM6IMnY6xwz56RC5HImKdavk76/sN6niIPciqzLNsPeJwXdGLDmEVlmvsEOpt
HFAbINEA4PSGIK/jr7LckPJrMA/9rDu3EJKiyasNdiAekSi6ebICNFHIOGReLg79
/OuIFcKKE1cXJ7X6LZDtWExk5ATRIG+NTOCDUyYwuC1/bGItQNbzCT9qcoIUF3mD
n8ggv74Ag+FvwjJyick08ocxdNi/p3pTMRlSU/SrnFSdJajSjbzbf7Pn7c15CRJd
Y9CJu+Uc6QR46EOpYbd8oXvNhj2WZLVjd7E/7YdNemffCr0CGJvoa/8FWWMv0lAL
9bczpoZYfR8q4V8QPqbM6ecLPJyF2ORrsEdyhp+jt0sNhRT/aNm28WpV2ySYDPxk
bvtQghQqHZ5XtxLO0YivpXI8pCroXk5gB1VjSS+cEkCegyfJDBwiD75eZbFRM808
cGo4U02x8GRNgHHQ3bfIz8GHeKRuuDsNQrpDalLS89WEMeQ7bKEWS9HpaCqEnFxH
1iaQyIdApmaPCM7XGKFgEWLEbOazVh/TvLgZtUsE+E3gJytLMB/fTqTKl8RuIE5x
bNeFQF0zLmExM7eumMcHgb79LMyGXV3haLMEi3L7E3PeBNS8LUEQjxLP+QlpGBwr
cXs5g9Yk5mkY4OVBr2ybN7bVTTw0gTDSvATXLI0Gv7HmxWKWfIy+w8FXs9vqbv9H
s/w1QvDtqPPxLrzdu/Syc557qakrlxXfU8eFKaNsBTmv4utng5XfJPWdX7KE5nhi
kzf7O7BS9bkozpQRZfj6QkoCp8SlBbne3+5ay3vkbpduzZF1Ilsr7XXe5i1/PzLE
SCNWM531evOLO8goe4ZBdNw6JHNi662HQW+cf9rlgVYBpoNGDR35GhMdZFzJKk2Y
X6hVY4J1PjwRzgBacVPmSnNf1WTogLRONo7B1WzTDGyvbmNXyeA4p3EKVOro6Lsm
LJUkQhyDzbujTkpfwm11ZGwblGaK3dvZ9Og+ddQ0EkdsNCXbAa3SrnZ5o5nW+FCq
l5bSjlLcaVUwwBFHmxgqMfMfHTJn3Yxc+PK6/WXwvsTW9t7AdC+zuuloT7U78VcI
saHdHy5FGhNzCwD7hHTC7fxsehBVBH2cvuYrdqLDQTlJgNICq9zx7/Bp6v1AfFXf
B3M6zrQTjMvdtK6WjnU2RqeTpl7H89HJ7PpZsW7kdDE8nmTlcb24eXZTQrkbLdMk
Ks/B8rp3rJAI8dw2bToUPyqe/iBWAVrB6gENcH9yjVDxpp15v1FJVjW1TP6wS0hn
MqqCwXEw87oxvroQLS2UNuWcKHKzIDNMlMf5gXZPZO5Wxj+wtYLa3vW0nYRo9TJD
eFMzBW/0cCx4d9DMueGFNq8nAjeCdt3FjFXdkbTETyBKewE2EJ7X12tMTzCDITjq
NJvKa1blyOre9WJHwCQBEoxZC+2hJLX4bbnslaml1a2CVkOZjdu+JSGpxLiKcme8
NSTINihcZcMVgdmv7meQr/QxNAH5PUUc8Gmp22vi2I8MEUHytL1WbEm6CRsc8WtO
To7+aDUMjye+3aGqjlR3A3CdsWkEyX2yqwVLzTX6uRP5KwogMEGZMFJH4J4bLcbj
qXrAIWtyMyRJ7ka5CzLjdIf+29XTMEZjgpjTojTL5/4sUERbNpsB4lHxP5L1YfQV
3DSPNMJbVnTFO7RppFnDhZUnJXiUnSMzA8Lx1wWkdeEOtx7Cn2Mbwz7/ps1zZqWj
364S676b06Nc8YGjhXfqGr5KzoK52DiijqQSAx7jsYwWWGzFR4pgdYIQ+HOaIIkq
GP+ZDa+j/xYpJF4r+S87k4Udlp1iayw3G1FWGY15e5BWLau+umTxhyQlPWACtEe9
PQm8ro5gx9w/i3c01b6EO6OBLb1oKYAnm8DYuHa64t8gN8uGteYt7NFADS1S7i3C
rc4RvhkwznNocb+BJUhOTkURfzpfaQ+jWdGRJagmjYax2dLRI36SZCwvTlNfklPI
BiiUMhHUQVR2UjYc0f9mQI8Zdb7TkHmuiUw8igFG1B4R0uJqWDrak8kMjKlPVhta
MVPUUMzdE9wPT15YWBaE/DuERBu4z9fcj1a+Hf2FjhYgS0cElmgsoP+Eaz47GKGe
c2Mn94PNPkNam8XVfVCPkZLK6O7Ngor4LTiRPeOgD1FUTVigZHVi12qdet4Z+CZ8
qB6NPyNgtvFFGKOeH4y44kwbZZ1rk6uWCPI3qDGF5UfVgJe9M5ASHdFF9BGwLsQo
BQPhY/rNCmE+9Ns/bg3N84UyFtRt+GhFpS6FmbtzTv6bPEy9sh61B8JeHWAludpr
5ITaHoGUdVPtYmyyE5cXJxmwN/qKu31QR7eHdUON4luMxTOkPKD5fWzQiCQQvFYu
qEQJjaFPll4fsDmb2eddLc4hh6CUFodn55sfMPZQIhBhRN+NYK75iYZJBVOgc4p5
l9Lr74FJ45PzHMb5LWRbowbskfRTxs8JIEOPcvRE9A3dAqeqJqMf4PUSKaQ1x3l+
a9SbNeqiJKY7GS3cXvypzw6EuMz1aWZvtBQ7OUGJnGMyNYr/+BcABx43HpKvljRH
5NFCpboiJ3mra/SLhQbdHrU6n0b4fzD6KVsYh/iBX1Ls72uaiUSWt7fKFh6OPFGC
kQEU4JTibGS4oslc2ZCGbtpoFgNSHlaR0HO6N9D4akZ5KqgctJkNo7hlHDPSRHA9
fkNbsLkkSL8GpkdkYKcpxs+FrXiD7cZFFo9V6yap7qphnzCxeyxja9i95hPon1Q2
MetGbiiTZr8agRNmQeS/Qu62QOILicbPkxmaNu146o6r42xizwr3dNUSMAV1CszT
Hx8yO3rS5usUa2atjbeTtTSy6pR6Gb77uZzCYUlKZi0ePnREDeDX1Xj3mwAqel/R
OO7VmZs9MPI4HVBdxhbMQ7FEjY+vjyMA+rJ9Fjl7CoH/M6AKU4jX4E45JgIXus8j
q/AdkCALpUPO+MMR3SOb/d83OJKks9/+4u6Nk1VtGmiHn6kwtTt0cBmjdNN0/XPY
wBmRE5+QKIfLNbb4jpiD2eGyWqg1hubWrYyu5JCePtCbfCUfTcFuXGAjOvPrvILR
2rXUhC7FzQgZtUD3D4Fbk9JK21DVHeTdZmRgHWwF6/KVEpFtWEJc8qhRouJ03IGG
IyfCDU8YGYdu29FkUAi3mAl58BSkRbJJipFgzUKszJyxYu9GAZdwZ+NwcXSw0h1w
1HXh4dny4SevIxwGSFj1BePW1z4yP5lb1b9XPkOd1y7NI9wJHH+e/TOy/5HAxhp6
dpmuQUDN1r2ORI4K7iLUFlosFKGEkxJGKjnCZU8M+DH8i3SpBd8Pi/y+ypIjWasI
5eP3ovkHt99NH0O4pdhE9muX9joviW1ms4hDnnIpEd04/deEWon+2zlbQVT+wOe7
15UWNdt8FvqIR6G4cXm1jT9sB1DslH3DS4ab3Nrotkkb7k7TN6dELEJVJJYut6zb
qWLk4QgCuhHJB1jJKsLKoxnz+LxMU+z9AH97n/HaqbClatP07FEhXT78bNBb6rMM
i2+2gOkx+4ZZO9Pys6GChnZX1T/KUe5FSivQRSRXWKc0gAgkCwDhPGZme4rG2XrA
9znSZRNjCPjVqUpBJVSKvIA0Y7nUCO5wu0/vzgE6Q+BjIuHbKAS/BH95HHsbt8TH
hzyTM8ss6D8MjfGEPbSS+jJuI+SEJoNQTf5Z4sC3bXIZ3VaugQQhTdkZ5iCL9XoW
JYkLH7UM/QaF/Q5xFc11jGy359Dhn3LohS6v4js3HAaI9hnZIHmlyDblDh1x7DEJ
vp1ns+BYbdtpWQQnhQ1yxYVKkACBuAhGhopi8tAISRv9r7wkEknTUY3qospa5ZqW
/D5PbUmY1lTeU0qy9tkfQddyOxUhod+O90s/ZuasRzfEmHeebXwBL0mzBHyLrrY9
Fi4GedyBiNQUfM/Mt696RYkVSmyh0xaFIn1srJENSlRT20zge/xO0mkfxo3CJNPs
mtgrwkJaYUq2Fixh52+E2kuvZyW0XnVuR8btJ6FrzHxP8sMPniWekq4IILcoFZtZ
H2P2e2uVsbkT5mxXdSLekEtkzQhXN7gx/Nb6SQbYmiTD2GmNZ/m/ihpawb0jSWLD
/kWxcqn/8OsNVREdyuLc9Yzqtn6ju+eh/z7AZJR5/nPgUMxhh1D8XgC8o4+YX/tG
0h3WfuiufhheZUTPVI9MNFc/pCiVzGeQqGsBie070sO3/5p5Zdfi9IrBvhgRJd16
p4aORayN7NCo22CdMmbM3wnMlUf5bAS6CApqaREQ7SGmdErZ3LNhUIOXXrKZAJtZ
PeGBMeJAq5zhXYIDQeq0BW7ZtGto/dMLtTKxxehYcTSUR4+ThNgrYmdCpTynLR5U
4RXqcOqPGLRlMbX6jyy4y4LF46sW/dTVT4QeFpxyufg2inGhr0YppNtHXy2r4mbq
aocp1MmhPhBfR95rwcGNKxPNIVhJc5T/P2k4yBovu/aY3vcrfADbmS2P+EQ0s48o
nVr+hmFyxSpyVzcG6+jAPTBqXjj6ybD+AYYcIodhuFYhTPKCjbD1yLd81K3ooIA6
0QWsnjFSGfWRIfALBKyGGHiDkzlALxZwKb7I8xOSc23Kn6X+b+TloeYsEMG87DCM
Q+jO1jNsikg9GACKpDbxb6yWKFTTyMjLWzy4PII/FKFLIH1cH6jkuIMpLgiI1Twr
iO4KneFacTAD1YYtjhbzLsfCpfhsRdbqxRRzMxw61ZHamdJFWebZbpOfY0enPXsK
Qe1Ju1Qe3YskUdIA85YMAikX0msPa4TRqkbafs5qaoCpota6fq3v2qXxjJxJGqKx
aRJjTKjU4g+hZEx7+OaziopAS+tlCOSeU76XNU3Jev5/nlVKUkfJwOXJ6Xozsldv
JRDGpkagKtc8jMnlRztDDXFLFLj0HDCnFnqkup0mEhuBr+ZeZ/2PGYjgny9y8zmC
/a7QVovHahHUoWwhQ8+zOY8FdRLKpCy1Kh3gWGZngk6xhlnXaMT7VuHjGe0aSFYZ
WxY/dgCVxYJICsPaJ+MdfDtBP+j80chGBoCXIYL58leJx5c1vMiaa6xL5IWLNCZX
tfRIyFvPnIDck8wUMU8ZYsx+CiYlesFKQHNdEIEgNBNSwFg8jvNFpuDVnVXulU5L
I1Rp6fUDI3xZEp1s5Z9A5p/P9mF/YK1iOcmZM4G4yqpC0w3HoGdi5+O5IIhsBM0Q
PjvxKqs3ND4WVHwX/mEkfqYrYR8SMyEscyDSOBN0RFUYJ+gdGy630KIL1cUDPnK+
1BZ6tQ1k67ovUgdU1w/e9TAykrGQQxhnHXjhbFlOOMgTnyQ/qPrqd1zH+hC2b3F/
eBi70+2yZt6kMlnXnSw134Trgj8Y5pwsEXYiYF52ypNRqJFHVS06brXaJGwKVz2A
/lnSVSnh10qOKT+X+b5wdKmu98vNXV0Csslk7k1HGkGFx5yM/d5yIJqbotdl2Hc1
Kh0C6zrNK2ipSGqk0PSolQLw1gDJoCg3Be5l4gf3YakfW/2DmPmyOa2YRNAf7pom
W8ZKVgZw2U1JtGoeqR6jWTpIW8ltA4rg6KdVPaNKZGUGn+0uqrezzg/BCT+YlmT+
VPRQ7mGHShX+SHfy1Q0/l7ylFUB9BqHhyckEjO/d9NdomaLCar5pqsMA4NuPYnVN
VdaTnQ+AC8TcWeg9Po/i9kHrEtvmWbHLt7kTnRR4bGA7wIlZCs10mpNhKTueeUxZ
7LTKOZmIPxTs0FhsmKkp46YnwYG7HUtdsaJy5I2nS6w6BvcHnkNCktShWpGFyyp1
RWdfzzHhjOdJKv4zWqvrRfiG4mRkNmLn8dAC9xZN2/rWiM6q0/RJ42FcLlVDk3iE
Jq5Ry5v+1zUkdhldvwLAYvzrasnsiBhVGT9Q+UAY8FvxZT2DQSipc0ql8lhuTxp0
6UJx/mmAhJef0OZFUMnyXZtq/8w/Puh3UOQAl90U+FsNnDw/Jw8h8EB8EhH/ydSk
5huCwebbBmLAZ9PW/Atdxw8juVMIbb6SZB3XE6RUXmbtG/hcDsfNbYoZhqWjBEQT
Dy/pTpVX1/vQEVHIi+YSancGu6pF0SgqHs2NA3OdiXMA5pqI7tlpMzgE5thCjneY
hR/Ai0TVZD/u/UxIsNSpkdMiiHNi9G/DaKQnBeVwI/jzooPCdMFOF1NKzyQnb8Dg
kIQt1rluY2PzAZ8TtKpuhYeieVQsNdj5bKMXdqbGUAw5PMkCMAxz17dJQRgE2zuk
7rDoI0R40LY2LIPy9rk2jnED8GCOJbmqIgcBFi3azPUd22DzHy3dJigit0soNxqD
cfj9mSrnjSdg13bNb9xfYz3f+BYF9jV0I1+L7bB5TQofY9N6WhNh2NMeDi4msA8C
worTX0cS8nRCF1U+tjxGcYAp2dHKpcP5FwqJwu5oY76AxC9zAB2L9zv/4b7URour
EavbWGFxGGkozFkyHd5lOR+SqXXT9+7HywkGGQa/Ur/pADkoAbAYtWzZ9vxaTael
mLkQpdlCM7/kvCSCb61WFEVjuzvIUWg6SH/RXnG1QcEIA+UJ9St+yyVemCiZu+lI
32s8VZQ4vFlTOSrl1FqWYKR5pgY3YpFR6BoxZxeqQ64vP7fjm5bMeYQWx8BZFr0e
Zr3BKybyyBDxiUpNKtf5eipW3bhUbN/ieNV8jK21YPgyXqVj4quql59h2+4ffeKp
KAbGa7EgOzxBg+2E8GTlH96vf0yJCjQJQapjmZkeduBd6ONkcROjeP3gdE+fFNp3
CRvv3TVU6I0/xdLwQum+fUsUJ5Cmjx8yHln+aCar3/pvCwKKmP7zXhC2B0TnPTcR
S8xkgRy53pQuPT5Uog36c3sQH3qYuQCgfr7h6YhnW0TiAbrlyN4jcwEorChxfVsk
wlhIu/gZGvnO6UQHUTSkK3DkLsRLDl2JeYqd8sP/gdIproBLeFZUw42IMTFk3kGV
ZQ+c2Th0iBBAgiAjwyGSvhGQRaJYbt4i5Nr4ubAqnwHa3uj6ohkFVYhOS2E4CFcV
/8NEolAtfAIIt5fpTBWBLylngmR62NNMxZTGMDx1B+XXIq+0ZKn/fx31ShjWUqL4
JSCwGFF3vUvYYVRPdz82xWZr5XQhJk5tXlNX9I0TFnWaqcZWP04G2JeDuGv4UMZc
pOEfETluRAIyjnGjYMJbPUSmuepggev2nE+idLF0cwNnxi/UbAxKUVxXvBe7xsJN
sczjRX2aXIA/FmHUJMrwYQ1xJdu+6IdLb64BCkxa1bKpPVU9dgXTvITarvZfd4/F
y1Te5DPO2jKIeTceNES3GaPCbBoTQy5NPlRwQ5zLd5VZHXZEyU4fum6tdaXpp00Q
jAObklWti8kGBQKTGKvaWb1W3fQSUFIn0ch+bvOhVTElbPkRwhsNToTc0VhO9yLZ
TxPb0MfnBjY1EP6VwCvG/ff11Ive0v6+jj/KCUeZxVSJgrF/KzgrLvPhuHpaLFR1
nLZMp8ODoa0IVLZYME2BJsrOW7rIPbtVM7LFmRxnRs/GOf0XSIFlecSNTMG2VvPX
xybEyJmRJfqhftb6d1WXvt5uuHUt6ydyMwkz4Pv3+rMOWgvKjJCZD+9T5V/vws9L
hSfNeGZZFYSJeOXTbJd5kDmOn3Mqjg9jqro8+E+t1oG1yYtsikufSILDw9tSBKq3
ccP/DVGxb7Vi27wGI46nGIfFMghifJlyyQePrsNl3GqE+7wXoJr5AhJHdaguqexk
OoaQRr+yTgkCBMC+uUFi4RTafLRYmQdXw1LjhzwP8yqTjplI/AH+QY0wKuJ6/QMD
7X4w9X/mxGfGm+04gG8X7lK93L45MxDz+Z8hhtBj5oa7W98dws8+jEJ9vVLjmiYf
acu5/YG8V+QPXJJhrSrp1+gPnwGcrfO5lv10df8FyoSXiw/3aGlYR+OICU/DUP19
6p6DdPRKAYgO707xZ97/60po7xCA/4q8RaGyXy7+hVsi2qYISS5b0dcdIVxb24Qg
2Z1K5GnaEeShpIxGONKbbZBKEdFXGA/w3U5LguJVZ0MuSQfSA3X/Ug0Jm1yv0Q8M
tAl2kUVgwflyWb/KeJNPY5hBRisU5qDhIOS8D4g3vbIfKQvl2J0GeImBlm2dE5g/
7r+mTzpnHacWKmgzvKo0JKRkd2mPYXGs1VJx8JtprQ3ATCETr4oYrjnpwmSLSn5e
yQ/i+Kcuzp292LCVTgx3dMErKCS/k43Sq/yQdzSnsCSyhqUDJ0v8+9Y6zppLxD6E
3/8cN0GU4Kh76UzfUgWQZ05iDN0sQmf8e6q19kSOQEi50NdTVxH6YaOMMlm9zAwh
HHwkKB6mEgOZPgmF+BGqfZZftArzQJR7X/sA9KhfkvdaqL0GlQbjmL/8Zv9Zj3ST
0UJdeyOSsWs0EOmBep58ZmkQBAJ0yx45DYCr4hCxhRsh2i2IovbK1Q9EzYTfxloD
5QDk6bzn2/v7oFu7llRoZMgculMEqnF7BN+Te5o85xx0NPXqp8peu/sYFYOHoXip
sMhkTYddImJuT9ki+teplPdcDOJGKHlIVaXTgE24QxjZhifayGR3v6Ncx1PnTqU8
ElSqET2EkFx+cuCFcrDetCPr9P2NAVSiykeJyKKi9mRIiuM+hbFoGXs4GckbvBPV
SkJoHQ35sTGqFUCEbaqpmhIa93cNUe2ryi+0/dz6kpAIPqQDm8yaoAqeIoog3Mq6
mdZ0gnFUJZzLWVHZeFdPQBCblJ3AxOwR/aItsmrOa17gm3+OXcxPcPOANWFx4AHj
G9PxMVpttbNkH0DrwWod1bQa4U2aKZIg2hgS9s49PkKra1tdU3Ap4baGpquTeyF+
8+Os2/2sWdXCwvCx9A8iZTqt3UTf1X8abBZT2GF+crkBbUmMl+DHD2wVdwtuCb7I
pZlX2vizRgS5/hO6BlDx6WPjaZXV9j27d3+oh14qgvAqW8jTKo2QA5LtoL7wpqev
GYoFjxm1C5LZw5ax3zB4Q4CjmdDnjZ7pERFsWlFlJGe9G/f+ZZeoiZD7QOQjwhLZ
9czTl6XUbSbAxfEl//18owUpPmZMDaGv/DghECBKuYzLXeWNlPjG7JyYiG2owe4S
E0Go8feeudwkmSmZo2UTqzp7R855SoMsRsnT1Qw3yk3GH3NNEA8FfuO+rOEelCJD
U6vnij0RqxIzRIhSPYm4H/tYuM7bq+diH3+lKnsgdG8la/TJIIr1/d9pgcEPx+eW
2eNJ1i8dxBbR73gSZbnBMKA7GFfqdXcgM1zGyr9cz9HUwUGoJ61dsePqA+/R8Seh
hRglpgIwNSq8BBzZRLmIRrZWwsCf0/YU6hyIu8PyXDySiwZlNbI4/j8FesoOQ+qH
zzZXjd91je1SJbR6DO+tg4dnMWMDDELxDoZDt4hTLSUrR61U2l5ZCGHs0ZBHZGU3
hDhYdN2YMkmo3PezxTSh2n9vmLcJLpf1/w7VW4DsiKrYKrncWlcjg5rJJi/3xy8d
tsCIhvtsAx64dlkPdyuxcUQwhSYIODpke4dOZ/dilAlAtHF07DQmoDvgEPPzHxiF
zoPQb0z2ktm9cH5xynZz+53dhLjXnW7kmtE/HP5+rUDcXG36wGQtVBglZiKdilyr
3wvrpQdhSq4kOA+HuYTA4I34t43pdy1H2KqEbx7me1G33CJe5VR0sOe3ryW31NNT
2pmaDAW+Vxe97WzdL147x/hjqV6FoDnU67f7hLJi5NNE+hP464lzGsptn/uWSaQy
a8S/pTWKo1pkIMcQMUkJiVKjYYeLTesOv71Tx+RmbgF0/DqsSEFuYPWGQAMs66F0
gHNh1xLmL3k+0X1iLLdhz2YABU7E7Kts8rrmdU27Lph9oasKeQcBS1wj0ciI+9Qi
uYIuKS55EmUOOxWDsB2Ajp8F0vB2Lr4mflKE7ewZGNiV/t6MlGIknBX7XUIHz2Cs
o9JB56Bfh4jtf285p9tHO3sCaPNltu7ZKjtkOIe8gyYMzdnHaxw7Q3Fi0SdhrTNR
wYbLBrsxu5k+7gNXMjnJYbVX7OyOMH7zSrysE8+R7Ebj8/pk5crix0v6nGR/4rzT
uY0T9fEffUQU4l8St2ftX8XgYVO+2YwiZjyMBS82CeIJj8pc5Zc4zHIbGqL6zob7
G+wsOjw4xQBn9OChX/3W0+y3fWbgHm3psAe1EfXIFdHDWsNpH3/fQvBdvIqEPDM2
H+WSwQcLWMyU+pfnNOVVt6RCb+bpyQPUuotRKXAGBEegZ4MDYLvsdRYO2Q5u/5kZ
Obo2qsbNtcus4NAYzNh4ZUoSTy6bvhHvE5wsyN+/smW1PE+NvA+PsMfKde2v+z5R
uL2r2vGJ9G7tiI2sso3e3yMNSMTa9TDDDLAMG6dWzqulBfZBLSnTZBdJotMdDz67
lZ23SZ50BIcPpDRF68nU8arnBf1WgvAS+6vx0QtMwxu5OHRBJww4UlG8s6MJqp9n
qB/dE1PULhwNhWwwfDVuqLxFvKKW4d+2ZYTt2cyWYqcg4Qg7hlnUMCTHJffPEL+l
oETfz8aS1PkxTasgLSX4PmZRfBD0BQGJZ7zJvsuhNX+WBhaiUAfPVS++dNRyY9hD
nbgh0Mi3FAPgNH2u5TNGkQ2bnXezJ2N/pNE1CcIYNr6MVEOKi5efnZHbEnzb9VIY
eOKY/k5MpB6w4LqahN/oiel1WI0DZJkma420VgDMNPgayl2DZHFxCsHZy2ffQ3KW
IuXuZRPBwa+Ad/Gd+XAMsXCX8j8E61bo7ljlz2U5LYKIp0t3BeAbVydDjoR8l//7
qHKcDf6OSmybm/4a4ht1+E0uEogvKAMIc4TjxdzzlpA1uSGOAXtuxomLjPD2oZmV
s40arWDdAnTtNklU8JR3498ZP+pGir4FAjCuHuyFk1uqhVivHVhvCD9jcK6SG6wM
VgIVpXSzFLyl5r9AVRwLgW9ybBeqRVm6M9Yl6nVZZEEWiozxFTUfwQKfcivF9Qnx
ZoD0H8NHBb6WOPEegphsZ6VnDmtrmGDTUBeD+m9iV5LMAVWXIdl70FE4W71UqFW4
dV4in/FaNHIBD3MKgqslQvtKVd224fHxioy38xlmt8MIi/eW5z1/tjs2BbRIgZ+b
/KHMf1OWH4wyTHUCe9OovmcavNQykSl24So/Huq/mdSuRMUchX2EMBtoELil9KwO
z45rUeGzraLQaIaNQanUi16/cWtdX1YVg91BpD8dJo8pk3G9yzy/IHQcCwk41EoZ
jibKqATta5r38zdiyWExvGBgoHlE7kI6id3ELnzfRyPP+QFUpDg3Uax2ofrQR1F9
3UpjoOeNyefpeo0Vw3c6JRtlEFuZPYpVsMhJSOtph3pB9gDi4QmBs2WN6wHN1FXw
Sd7RioGQE9GIghPEX/77tOpfG6yIWvnpYyvzjHmzG1m3nGn/hBV9FNX+1l38v+iu
d7Hd1Hu+SjPQLqiUPac5fH4ZmVRB0DgypOuLQDj1mJz6cT+fSR0luu/4RK5ufker
kfxDK2HQTuqzjTAsiVoGPPpdeT0oxKOGsylfCffTWIjvaLLomJ25bFtBWnuVxKVr
Yg/ZZOoqd7j8bE94jZCKhIglMwlKn3GVyAy6eU6y9NpV2fKHjCXRGJ2m9oco9dGU
zSpkmedNeYtEovjoge+arBYtZHuE7qg0J3h9RU9fiNzljNv2j8iFaPXlh4TNHaWL
X6mi9N0DVTsDMT6Bd8Dql0Iq1OsC4U/qLZ1mps/Yjj0rCjSi4iyXJNNSEtw0TBBc
jJKnm4jzGiu6igOCE5XwqiYET12MsRH0BAc7WrDIjkVtVOjUCf6okvklbbEGhgW+
QJHDFoGIC1WQTQbHHYjje0ajBN/5SWrx81pBpoOfLWybQTiE+vvs2jYL+NUfdLUd
Sfll4JOQPiyD3dEe1GWeB2H3uyWxXHY8kDanjlSVfucUOpsH5+4Sl9G2oWRJJBaI
UMG3ZgpSADfe67bh+Ebb7TTr0Zf9zsDfD0GV+oBmeWVuVPStHPeoAipPXGUieuHB
wHarE1JYKG9pIr/eCNoRWHe4bCvCurero/6R6BG2gjd6IGZXEz8irq3RGKUzZIJy
Yy82wB2ypZ5bHZuHnks9NEyJHiq4DfKZd/5k4PTZiNC0AVraULHaiTGFlpxoTgx2
+pqXdHjg89/LR7aCFHqlN9VIF+tnMS4UkTbtOlPfr8jbokZnG6N/2PpYYpHfICrW
4/gT12ChmBOfMVxCsv+x0RyDJN0FbwluEd14hkTLP3PmmwouYciFAFhj2gEIsFN3
odxBKz5axI/eQBYjvz7eBh8LLAclwM3MXPrjUgDi/O+L1wzo27N6le2srPTy0Cjw
LCpRjKwAc4kqJV7790It4mdvvYFlBUnX37yT1ViKM00qHVw2E106RMGIBQBmvu1p
tnKEVlbXo4NBEgBJJ90NSGmVeZS2G6/cqmNYCq5k2W8M9mFPXixHWaKL8Irxw0wd
qwtVaB4p2x9UbozUwaMKM7JunLypHYq9pI8lxdyDueJWiXrOVo/yGDe+h7IOgNgA
efCenOzeZms34S6gl8W5mTBh8iS+wnHAxspKVxWWx/bfxEA4EqufcUOm8Ds+azKD
CkoqsMn4TppW8Dwq7F5yCSpmeWVHCeE8jRzoQ+zs0s/DYCleKetE/AnowKGfMHbl
bsApTaz1RWOe3kmOqlY0vBB9J+UeVkSb35jaFstE3bqG9Mrh9hXK8Om4xFRg5Kz4
KSVCx72twstglHnmYcJoNJYdmhjQkBh6RMUi2hBgLKIjAhUPQBQEicFxfYxeLNxH
uoPpnhAeh1JQDCD31ivHFCh7SDVSnWlQ0pHDvdcea64RYD//HX7KkwChRFkvTWLI
5CKDu6/Z5Si4YMRYKqKT3J9wqLsa86xU1GUhzn7HufB5Ve48tfMBDv4UIed9AclA
XFIJbg57JDjOaB2yb6yuTIWyi3qkvRA0NosUVgyxXUxN7OGVX6zuLerTtJ8FqPQ7
quB3cFItn1RQdXfoXd/ejOMBYbpNewn8FPm0+UybQpUALgv2S/pxRT81FRInsews
JAPJug7P7+BRf0w74FMINXb3ZzwtKWSef1EulkULmeROOas2AuKMKo/lAN01izJ5
clmjvDbzfXagm79+HInLv4BWCNiBxjMDgcWu4ebTwcUaBclc9sbmaiDF63vAl8z8
V3gJSZLJbTeuszVQIDMaW4my+rLx45O2xTA1zhSmwrlsZNrlepsGJqCFhI7uvjq4
v9lazFQ1J2Q+IBJBPt7+tl+8UXfi7qD8WdxDt3znrqhlf3houjGx5W2KZkDshOcY
HorLSdkUH0bbi8qLk3+FZPB6rhOHJHxWwtuya3tDqzBGPh7MPIus+5z2aPK8t0W/
QoPGG5gamKNj4MaWdUlZnU0cNCzTB5cMso30G3W0kjbwdPi0H0zM5MUZaGnGZHLX
BqqnzGCSzGizpfzmvQmOaJOPYnJDSEjNyFJ7Ghv0bdxOUOpgfCb6Ie/Yn7p/msQ5
wS3FC0v2NqhNF2HtvmGOKiSYAaFLrBRIidneJ8Ckv6AE/TzXi6f+Vm2RAxBHgpT4
Pa5UeUx8SocCfjBeL4LKQY9tp0C8PLthNSzfPlH5qVqcwUDTFFDj3zfFnf1sIctF
5eopyZiX/NMlHKWvzfjmEJVq6fgqPO1inPJf1ZYY+/9ycJfQ6nkBovI1U95wGjsW
U7Rx+cSt1nNSCaJ1hyiiGTDo0GlH8ZN8HWEfyZVdhPXeHLSByFW/EhdtI+WBohUb
NWbmUXiJJGgkbuTrRYD3lH04B8teHMMmHHc3o1jxhgO8yZWJlITXa87DffLiBjpd
Mo8sc+bVjG3zNqy4hey55VE2rKAkmmOVWeeN5HMDSZfI7jUdgTIF+2tbGTvf3BG9
07thfoBDkeFBbrmYQkGK2+yzDpFnqk3tgS+7BvWqq57XU4tHo3JX36v+ULuqAmML
+OkSNxK0FAy3xjHwy6yFBZKB7XkH4nXSG7VhlGOXwPJE3zlOVgMZa1NkLfsGzfG9
T4Gs2jnuUB03zc9jL4XnFy8JJmhGLZlB4MOKcf0qENfEU/oZ7ybMi6BWTQmrF+3H
WGLOIQo5UPZ6rXbr3GpatMiBixoiVFBJLrfQBddvBNpb9s7tp6hjCk8sqGqGZBek
v2CmQviKTCtlPJzc5uce4ZMVWhvWV5+0knAYtEC+t+zY68w2NU1hCpIBuZZege1H
ElnDtCjHRQVVOlvlnEUfN16U6L1RBaeKoNZZkd5kcmiMjiujD8/FFyT35QZj+Oti
21YbnXqJvi4xW2OBuBAYzLoGGfKOUxORn+WOvMCUm85N46S+s7xsiZWME9YMCFnN
8h2Xo3T+/RsYq6FYM/rthh/FM/OTCwaLfzHHsBps4fwtJ5QoWFODgJBHopzg9ey2
77C9IvGx7PFNtE7IJqcOFGFyTY8Bq7kPk0t8caMTsHcuqdLKux/P/njZ5Nk+cQej
L7kmZxyxVSFAjjXDIEpaNWTyizDQvRC+zrfvk2U/rAtTBZ8mPzNH86SoQUsuwbhk
h7eUrpMgFFhSAXg2hl5SIiClEZ57QhPlXXoCNByAfovC9F1sRJtxcJ0yeKXhajGY
pHvqZr0KGlx+a2LgwTonx9gBE6HiSrnoSFONdrbCQk4Ck5+LC9UlTx95/WvsclTd
HXA64fFv2ovvJutWl3F375pe2BVIMgIXnKVG9wAmVO3qtH+GpTPcIkdBuspdE5Wq
ZGh48PMR2B2M0Oa9xWv6Jrjvy+NlYYbZDneVKwlqTENP3dY/e04hvv4IIXEcII3H
K7fiZvrl4WB5UOhYO5gE8iKt6cErdyG23AAC+TeZQPh+JsW+N2JW/2UDWpssG1LH
FdA7LYbFC6CMFPvAfkuCuHYrrIL5eIl2uVY2hm4O64aGRAXBSPX06EB167xZPvZA
ME5XgPat+qb6iy69dq8WXsfB//5SYIBzUrdCrbPuzY+UJfLTvW52nZnt+kENckD+
QLWnmBLQxJUgTdRIbZ3wDvU1ajRi0qTjVRVpD+/XnwS5Wh/QWbMadZYkP7oaJEka
zIlem+2C6uEYE0JVX+lfjDukyfz+CcLJytSuKb3AYaMJnF9d1Wt1q1StopyXYg8f
Y4jSW+l3KieppTku6I9jR/AY6Nf8BN+2y92e/yBV6KtkKUSBcCNK6H2VpTePq48N
MceqzZpifRxx6Kmmbi0KqsV7QACqFe/qxcTHdCRk3GluDV9qix0jTJEGy1zfGNAQ
K9fJaSnbp9Ovwxtt5TMud3kBUxY1bhIS2zyXwls5mNqPpD9hZLZZIDCIoR7TEVuL
4VUXm3Am2FP8baNPjXbNRJnrPitVwEUTAI2DnU7SKFQYGhm5EbvacVDK6Czi1Nic
zuJbeV6niMaxv4kQKgu52xKuvlMTYhFLrepoBRPZ90jAXcS+o6eSX32f96v30hSZ
q1s+Gn4pQ3o1pM1tBT3l0b3OceFDaCahAm1eKYAV0WrMjXvCA640c+AbQDMl4WmT
6hRGQDDJ7vBPyYK92C/6VZZY+v8kmgf5ysgT978HUpJuAlSIiMsWJJQOVxfWAnBi
ew0ezqdLDe10NF+B+Xvjwb0/ztjEgVOJla/qmdlOnRC1Bv+iU3xI9DebmvqkwgOI
JDXz42VP+iZQVph9oiYnPtoxuquz3DJiKZ24IPCeb/+pO2/cDqO885AUHsAAVom9
s0VOWmZ8UwOGRQwsNL1TW/+ELLhx6deiHLosqINvyv6k/AvRdRmPaSq9iPdPnSCR
PTANBFifpLirHTY4hoi4zCsDyUWSxHxmBrwlXCo+dKJIg2I05GRxhekl0VPLqSV4
lhVFXyAvT5gzjvezsxG+EXT3JO6AYXdn7FM0P2p9vlUv1CsIR8C5VIE5CefPwi4z
hprKV0WQn6iCFESV6Y59OS9rukcgjaMWXA+NqXfMGCu6zF8ND+Y2d9u1NoCi6ObW
q+1sHEt9wkzsZj2s1iyd+CaPloZjXHalP6AlUZTJDTl0o+hbhXTXfQ/yKnEaazFT
LD9GzMeqCdAapt4yqctVHed3Lid6p534FTnNUie7Yy3j5w88p4N814nj8DdhgXJR
puuQ6v6Ly0j9xq6oU7yDG/naDehcm6BNjXvMU3LmGgqlI7ANv4P1M3xZxaJGQdd7
sgm+wnVJ4VkEgB7GqM+o6lo9gJCVXrbGEZ+cFblBRLUH/9E7tVqRjAXLKk8pqSXT
h7FugeW/BuAALlH0Vx/zeqBVcGXtu5MnD1n8FUDbIE++wpmEkuhY51E85CtC9UZn
F46cikCwn7/V7hZeq7xXHslOah3YcjgPO0RaVFf5eg7Vy3H7XxBIUgwyneylVeHs
t/6ZrGR7sCIxJrVU0ZQju+LN24o1IAJ5vbK5dd/SxkKf0+Lwu9J2uIeETdzHIsVm
8lLrW0/ML3qZe9HlgJ8qSDSL0CdXRX/K6U6R76otFweGgvGj3EqejoWwSk6V0CLC
hlcGJ6c55OfXxc+k0Xw/NNaEgLXTQegQQrpzNUA1Q3qJBv3OiRnAEPVcNNmmUFoW
CyqEfnqLd1NQs+lSlLeQGqNn2+yzX3m1dhH0ZKin6jbVT2K/Aaq8rvGJH8ai0PE8
gzgpNIvNlmrNSCti4dE1qZ7IOi+GKvv64ssC81HSvG3DvJCIdSa+50ForoBrZaYi
FGBJBl1UGUrgNg1gEsXlLa5dLBHgS23f6wL0Hkv+NspADV1r6frhEGSr/7aYt+M1
5EYxPnaU+exl4YxO/Kn8luWXQxDVvCUrA41rCpvt6uVjgGfInjKjkPH1E1cnbTQs
ktRd7cNPwoiJ+XBU3pskkUP/mWrryDTXlg4SKg6YhUiBmFByCIsLec2A/tQhNK5r
I6MEZzjiCiv4v/aVu8cMjuXjo5rg3O4aXyDYLfmJfwFCjp2zS5RvHYAak7LK8GFU
KlQRRXfEv+kAfWPqHmG/QWqRwVvDvpU1OmDBTCeN0U4oYYjPhN7udw/L1ZYij0+c
+kFTIQqUlp9Bb2Fcy41Rng==
`pragma protect end_protected
