// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DQEEhLDAoiw/bN05X3eiSvtrdqSgutXDAm9QXD7LARJz69e8x4ffHcB162zQ4Jgu
jGb0EyZWkPDArwv2ft9miylkqZ68vuKKncr3SycHY4yxe7b3kKAhN8SGWN5kkuLK
20nqsJrJDRlEJT6s9LuXaNLwgt+qjTpTvPQG4JC5RNs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28448)
wfxMnBh3iDaTfvDTemPQCeAMmHC+B7a96DR+d90IE1Q3nCLDJVDNJbgBZey/WrlG
/krWO2GAhktIbkYLgD7wkIuncnJMK5m+B6lWyQZSCYqmLDu8bgzIk3f6DS0sv1TF
zsrUkqscviyGd57CxebAy9lQ1MHMaNPlxfnVNmqkhLgBb/KbA5VtgiP7Y4OberUN
42IzerFvlHS0NNxS8M8Z5aZYhvKi0RvZPpz7vSAKzZxQCX7U9L1z4trE+Pocz8We
kL1sJjS/EQiE2uy6/rriV0h+8Wphhvq4OCgZ7TPc7vBACA1pK5EWSuxv6EheyTJS
TXKwYVtNG13QNRQx1NjrxzRKovnBPu/J/Dx4ileUTUUeTV1lSumOIy5jUh1G/iih
cpHrPffwN/8MugokLDq7dlFwUtYuS6Py8YtaUJZVi5DZSfXOEknsRVGK/rA/RJE7
vZxJyMa/8i1ikpmX+iSYnsCwvhh5siuRhi6y/ZgGgs+BbCM0BsCteYsBhmVHwpyi
BfQUYP1Oe6r7B2yls88rwkt5TPvDtThUsf5xb/PyYnjbId4Ml/vzc5JOQII24Fat
+kQKo4V0SSC0FZxVNy/7JGOZ+AkthL4Mbo18h2otpL6xi+RTp50v8U7Uoe+o5gc5
+ZRc9HuFTsvhUHt9rDMV6qoesSRSa/WBnC2/qFBy2b873uT4Av4Hn2bCbYqm9Vhf
glgjh6F8MctbPilzj5Ee1YKeh9mQIZB5zM6FrM5whi+jOFJ+ba4afO4m73txTl5Y
xcsV6x5K33L50r6ioCB3Zncr7EV8YNgzas9Sbu/ufheHRMLVjZDfd6OdPWHSXO+z
VdByyykqujVxr5fYk5l3wN3ihd0tGf6C2UuuZD/9lp0msQdTvAkMNQ+E7KjWb61j
yV2TyMltRQcuG6UcLhzdSXlBYDlJjfHErVV7vHamfSbqze2tG6ouv/soMuQgTDnt
TCW1XKRKUAcN02gcwH+Wb7Nku2SDu7qP8jkn/umCSHLtCbjmz8AtSZxVKzIdgPJ7
5mOpeZDUScX91RE4olZL3hm6zqn0GA2jN0xWIKNMaojMXe/OFFSs3w6sPMxYWgHk
+BQpwv5eAO3EnkCjhqws8gaCLONYbJn1cxPiLQrukOTbtCB17mUdgdRxCmraCyYH
u1Gt674Nt1Kk0VaZ5SHIORENakyUllN8K9t5eEYSE4lVWnQBdOuaMl8H7i3IlJQh
jsNNW6utKre134di5qzx1Z0u4rHIvnFrMtJNUXNV1Ax++JH5hRzevaCTTLSqQmW7
MIQo0nk0E4Fp08sxUOz8Sd178cwCGkljlCPmyI7u5krboZDurB+R5X7mhUegXh03
QWP38UgAW6T5hRXlMLdKfrulgEwxY2tf4TjRFyteNrmlrLG3Xyov6jChF69A7m6v
zThmHlNIO4nX/1nvw/BUI75St6dq+XtPaw+hG6CDyzJAYqEs9saloyDQfiR4ZE4i
frjqc8iuAXPeMFQHS5V8LfrI1wkNCoohmfr/FVJIWviCttupuha74bfK7Pb9hR6w
p75Orx6Xq9IDktrNyBBmqA3JDXodj5psjMSuDiBCjSlrd60umCtywi+T5aM/yX0a
9gYLWUvPNV9p9we31KSK8XKBR6pXER7o44yKj3VxwBxGQK+vi5I7S7yuG4h6nLX5
OO7jq5eo/Y+98hN9K8JT24ZVWUPRq25Nk2oLvYyXig5bCvWcYtHkBMCk9KuIm5uR
ru4DzCaTxRrr150hPuxz8aEklH6+3T63Z2UuZs3rmm96TshcNqOiGwAE7A8Hs9ex
4aZnIV+NdWxlATfY2wOGWFkjhB2mztU7bf3xNyuZez5N3qeXJh6IaG18JQ+7S8dg
4xhWBcoAPTCJzYQI9LiIIsZzX7ghas1apVJ/ftH9MlaI5k+us7fdFxSFxHk2ya5d
Z5IMykErCNp2njb6UA3m2Xr1AVYVwE/g35ItlalYPzUdbWPqZDJjDYxsbKOj/pjh
8ZbdoI31PoV7BdMdhGVoYAO0BEBhSHwDJD3LVBbP1P9QA2jPbYf6Lx0dKN+W7ttv
nd4sjC3idxJ37YEU17pEV0YHctmNVQzbNLvc5r8hgGhHPN8HwRoZedDkPA9f4Ckt
aPPXGs4NTSOqUXEkSZcIY0PARf5Cmd2fZ/peGyodYQBQ7H/m2jBXZSuaTmAnBv5e
TWioOUHdpRdwerIHlkI+EFLhs4HXEJaQtSba+vg6b/jgVyFQhiv2FX/T6BCiV5ib
vtw/9nplHkEY5CYp6o0rhK9EhyqH3QGrznMaNhEmTNJlU2rv+lKcnQXpKiDmD0cT
0/OL0hfBmX8ZwLv1Rjm0jcU55qovPe7qxq5br85T8ot+hMRYoUfXuRGJH6uFomui
LI2giqRjinW+IPQzhd4NBTb+Pw/nep5NMB+kUgWAVtS8u3n8vck3nQYb7qdd0tdQ
hzSOy8s3e+GaEqtPzrRiK5fkmXpeUC5pAVNZQhh4VnP0NnHaK9SNLOTKTxDPIK6q
eLuvf4kNvw1m348EJCRVFifNLrAz3pZYLYDI6mk9JBwqp02iQfXxfZsn+oGAs0EB
71DJzLR17q6f86smxNWXYNUStLJjy+0VnQzoowB6fOFoy/1dhS0yfz3QA8qt0LEX
65YzVegS67IKnX2JTUKPGRasRnU52qTBMNujBJHnVo4L6J+NDK5t4layxfuGTgUT
EY2PJk85D5IDte8HnEjpYyGFU7R2vgd5teZiurS15BafhSowwagrb24lSBj1tDt5
2KrjXew1fAzdNhMTYM1ZfO6DCLtYMI5lHQNSHRCcfjHWs+Ox6HwWPqL890oR6CpJ
+Vuin6PW0oB0cpEfk/IQuokFCfz5GKqr0c7+XD/ldPqW3NvvBSJR2o8EnguwYvkf
wOXnqiDHTruNnwv5l8y6gZyUkXGYDTPS5DjmU2P6p3FOgjYbajA0qMbrUiOXnHiF
G9aWvU9gS8DnMcbSCmaII5cmduVrnUn8xpTCLGoL1cKQcBb245yKiFuy/U869WU1
RQCOPRU55wAEyndi8zvg7EY6BpeW38Bht6t1hLSsjfXvBkTY+mATukN+mbz0RYbc
VmxS7BsH+QIhDHKvvvwl+fuCCXvnxKGM8uDN+peqdqVDaEEa0g3xzE5Lb/HgRdpb
hdgS0Dftcxj8D/jBCi1ysf7F6n4P3haCqnqex7ic29dsGpXxXDvqkqFZACU8h1Lq
axchAMlNrJ1X1xoxP+l/6SAXZ1+F66mD/+C3cUVxd77StPlTM6LT4HHm1c8Sexev
F6WAmrKixfOzLWD1t6lsBwKp4sjVy+0FwqXvTpKcKkLySlrBolNGrooBdm6JlYZE
DgtT3qX/OCxJbVm9u+x8rcgdz0swEBr31PT8jRgr43WIkB0Zy7f4EJVzzIgxNoMj
jWZyPSXVjMCKlfIK/CvhiWHOfbbTXv/2aZow0fj9T+RuplNpvE8ylyT8BfBtMKaC
cf8vr454rgRZGy7CFx08JXWg9/RlrL+foOg8sT6fuxZ/3ce3FADokkjoSLI1+++5
M8yp9UtZj+pbxLgW4twa7JfL1MOOkPq4JrLFgs9rUkTZuGxbXKCVcKvbbO0QMVF3
nZsfh0kDFuvHRkyJfvROM4BmgUr+yGJ/gaIEUpJ/STblGEhsVT1JdsmveKmiZHfF
ZA/vg+ak8EV07LtDfAl9Hc7bXFYTZUB2NZL5yr9xKncrWJrkT6S/TcJXZpPk/KS3
4tA0E9zKQqq3yn7hPc/UZDD8UOps4hFyRc3wljape8RdO887puals0HT1x3BnJeG
PVJUO35qxos2MVDov7iY4aH2YNA1/3QebmKdw0PNOt5+3vbxQXfwDLAS2T4jf7pG
T5on9mCtnCh++8nwep5EdIJzFZR0Xi7x6vCe7GcwmVjCaJX+saiLANXnHQ96ZMiE
NbJnF+a2WuaPagTUhIOkzJn8wKsxtryjcL6pha+hmw4zDogBxGsDCTIBhIrCR6Kr
lO1oGfLKWia+5pbOYadjUWw5qPV9PWVN0u+NdRir/Z0ePoyJomc5klVZP01C7avy
UrKiYJG3PbpcNcHSIfo1iQvDSjha0aeO0xl+/feXMJTqK9lEGnWc+O6t8ovLe9LX
xhvWc0uzrJ1pnTyyVV7bC8OudTXoki6pJ4EQsB2fHLraDB1s+SwEGp3ZR8aRthbi
XRB6HNAZ0ctyM4ozq2nCdZXcFWDxAA6kV1nuvQVRgIfvGiXikuiLHrEE1NC9MZZx
QB6ym1BPy4dKvxEB3aYG+ByCxs3GO6qPCcQuO3wCQIXoleSSoWkfWYRtYovCueYs
XErrcghi68JoWt21che54cytS2ItA7yIBo/lamZHgbTH7EDOD/Oy1cUFlUN2avjB
4uyEMnudgirFyhMVYW41yIL0Fnh/7NHXokkuqTN87Q3ea3mfXBfg0bs3EE5wMNhg
3FfnC82AEdhy1TjJIbiFMapMcBSbd4+6iM70DjcVQgtTE29xYwKLcJfBqc9wD+q6
0vJ3v+aws5K3s5OKKtubY5Vdoe9MgXeNQM7Csk0b1AB9X2dBCQZNH6ooqCeCu/ai
DbfO25GJeE9bH/R3YMzMsgnCyzZ0c+WlvkYnO0/Lxmr62mqcl2R+sAeQ0p2OPqjv
2kwnabnbjhVQ5JcrvjKTq9ecerLQ49Np+4w5j7aXKN64NB6/KvdQOzBNVrmzAK4F
SFqHo5gy93s/Fwz3g8K/aksdXgGaWtj8Nj8Q2NFxAtsjlu6OC3viY7TAhbBBtM7P
3H52nu26WrlkibuM8Q1arFUJD2cLNfCruLGm1JB/FDTc4u4QlMmIRhKxl3frlMhI
xUFNYZaEt4v7X/tKnfDvVxqzk1G+tf8FJntG32ub4KuzZ+5KAPFMRI9OM3E9a+yz
dx4+nSDqVDU2p7i5b6jBBzMuwHmAjpvA2AiwA93HdthcynUOuX8g083PuVCEdgtq
52ZyY/Dz6ofADIQACogtYqVDOTRSquF1ZQRmhuKO9rlHPOkcoghqDzJlC0SdaLo5
2BYAhBVQZyL8wUJWs+0AUWpfYvLPQG4z55NFlF2/emy2ZTLZ27Td3DtSRQE553cX
GKSwCzRbjqBBoUgvEXV4HSwQXuN4TtaYYkRKd0eLoa6JMkSpo0f3+isoNa1iJxpK
52s0NDvijsopOJuPdsv3m/kq006ZWzYAtjLZf50uQ9CLVDX6mmg/sGRk6pRj7+8P
n4JCJhVxm3uFcWSLl2ZU/u2p9wYMsVwfehYGNP0Q3JnsMhUAowL44rz7fXZIQN2T
ab0G0T9+RsipdnPfQF9o/OOp4O944ekW3KDq7CgBcm2TEQVAzXHS8a1Ww15/Xq9O
iwEDgJqFqfBS34pbPLAivc2uKkRqcUO5fjyy1C0bnuKjLebMEOAnoTVEVBBWhe7w
O158jtDiM3Q9VG7EOKBmAlBGJrSGwMOl15T3KK3tgwJBB01A4X9CV9wO2iefIbnQ
sQ4jDgKSkY5sAtANS310BYLflVPn3qZMZuPj69HGMsNJE3bdvgHzr7lrgbeFqVG/
ChwyiXgVvf1dJLlq3+o44TazDWk9mK+dvADEhsawMSmrQ1la1K/YqTyJ2XGTq1Am
Llx1dupx0rFX6rvbj78S/NlkclkXd7fen+/nuSNaVtT0m0xuYjzXeYRci6m8ZXSb
4muA35MP/lW4dqdUrWftF8HsSlDVyKt0YkhIrweH7nWMh+xFWPKoXMKhEDS0spJQ
ePfELxcsmvonYTJE8dpu0rFpzsaQwQ++TfugO7WwxXPrBlxpypOEYK4iDvpxyxFF
scN3hFxYcGuGndj+OYbZXNfFiu7/+tQdBsCVB7JbakxI8n+eoKnxyvFhIxuzjZ3l
RNd2li+2yvTnkKnBKAGpKRTlIJ5jx6JUJe7T9SKFWjT0YWLR1FkmylrwgwOkYT3s
lchPlefVA6FCwR1n+QFQiQpbk0Y57htp0kSsBmtR3vnDbdGWy4SIH6iXf5KgC0iQ
g8pKFXyd7evDr6upMxwg7jujGOVXtnoRBBOdSC9KX8G5yHeT6zIp7lN1SZbG1lGc
csOihgdS9UQ3sj9dEZnr+I9R4z8yKH44V+iq0BO4lDmkXvk5PNIQ7GaIoGkIVGAr
bP/N0ixM+uwiCzGXp3KX6WDEJF9ZbNZ+VL0aHo2uGB6M3gDaWE88apphDxCaTpS0
itYvLjbyHFFvyf901I+YAap3CGIWFjRrj8+snJ7C79OybqAH2KkAbhWSYJW5ND7n
EESKDhGyxmz0nv9ELy8viTrgiNT85R6HXH6El2cREmaNUEdrFLGjlPg0XT4AFRZw
XmJ3QNQVGJ86uwnYbP+JrSg7iFxtW6Ss8/QomJFRS0x4Uy4d6DNRa+3x1C4XEpsV
eUuBinQt2ZGLEYgLrugv28Vca8dVz7m65s/OZ3P6LJFCkyfmrV8Sh61owbBrBw0E
wpPMmxipRqoavm8jlHZQ2Br6tc8Y4cg7xQOxvbR5+oKPKminGrTRF4zL+vUhWBMO
VOpxuToQlNVmIX06uqJS2oFKz5sDQEPuQCTd44tIY52wuCh+O7gWQIHcLGkM7rRM
/iay1LSu/HejckTNys5O8aFkyl5hsWvuedJkmmVbsrUT2jG4mwuDIKxIOHLy+5Q9
FE3Oggju7AzP1aO3f/p3s2Kx66IHA34XnObynfSCIHxtDskAb4zAENkKeNPmZsSY
oD7bjHNl3IsGsa0ckE2lbrY+1AanUYPaHdG5sRwIfyZv6HRCDcH3XkVC+SyL5UK0
KKRt68IXrRhrrAEVLF0os2Rgitu220C9hEelIy7D2IM7zlOxzkgVk7RT52xkp0h3
hyueUTIv7VTBWHmINPvD/q39yYAYMtl2PHBz9/FxJ5S6Fu953GO7bhNIxvz6jLUP
yN80IlMyMSOdNmODEnLQ5835i/L7n8NfAK2/sjy8Ic7Zhcxx0KSvxpAned4Opj8l
SY8ATII1DLKhzCCySUtTVLC8IfWxD9xUkj7fnZg0WN4pu/xsXQvwadRWdJwaUshI
1GVADmVKc3+xrUlUer/CDE0a99OxyR+dh9f0Cgux064Snj/3cpR70d2DBPRBSirC
bxU5GorQRMQmDNmeq7GAc0b6CGpR7K8ObwceCJVLUlaCOSx8+dONVp4cdldZbum+
AyGyWUS2XQlrQ0esksecXEHp1vG/YBPr1FfAVam40KBcEwNYp40jgKjO2gWkjMim
kNBP2o2P85Km1yVEfXcz0QeW3bK7sC7OOO3CJ8F0N5Nohu8xYruVQG37bLRybXIA
8xQmaxPhxrHQ25pbS95ToV+57Nq1NwFTeBonfM7dCHZeIi1dzLVmuH0X+nh+JkTQ
xxeVS4bULPTNRtWgKLXA5W/VP/lNalUOcsRGJQjFYQMLO+seVbk89LY6ey3nQC5g
v0Gi3+L2oOkHqpKgGSCtB6SGJESlg/5Ja2/qO3q/h5POZ2gcD4Awx5qBhUsANYKY
p//+2xmi5Wdhk7kvHX/CmAy/fA0Vri00iswbE+2M7PlqTvLt0b8xZxpAMJ3k918T
pdo1KDeRCyy0MT1H47Xf6cLsIgA+DirS+Fb3Mk/XTS7Cc2CmWMwFUVaTAtRCUrW2
TmouBA3lfH4mRXWL0ijo7oHLDTKeeCvMv2lq2hl/QOv/fmg/2ol39LQF8p5EFZUR
E0VkMjAI29ky4Um/4UP+uulZMck6cdkfe/ZIcIeRnFwtWFCnZG2M+HOsJFJhpGj+
+ijx+F4qMxuxJxxLm/1rSYTpaAfptm1hmps0a5GGh/4GNX0KIhLNUZOaWIozjrU3
dP+GLaa5/L3QNyWk6VS7rky4qt7e+DAt1U25E/DPn0BxBf9fBiI1t8bqoNeXVHmL
G/4LxJiL3M+I4tSJDorf+5pgww21/B6llyvP5bpbvMzREVDklB+CTbnYqUKkNSV+
/zPdt2sEHhitWjeWbN4U3mZjjQceKR38zk/dGqcdL0bI2rBPkO600dvf9uhX3RLE
AzD8aay68btjahMbreLC2ZIqLkuwAJWF7hzQKRiCOMOfDduB0x6pAtikjzNVzn/4
RdopWPNqndmJ9F9JYtjoJI2K3j4LI/X4kAri2hLxlld220+AFjPalHN5G0PRW/1s
DUMry02wzHy48Kwaz1pYWil8bsOtaMpQfPA3huGz3UDKYe8wNAK7pXpbK21TM+2a
1r2FwmMVmcSSWMg4QVEfANNB4OeV6Pv2VqfyotETP21ArAHSEmyM/nAUgGvdP7sQ
35l8zU88ewccxudqLpp/pq3vpd6d5IfcCVoDfybDxZ6B2c7WDSYRxiKQx9hIyp+f
oqcqfO6z1N7ieJ12aQyEB+l9kt6YU+Nm+rEp2x9p0z93jy4J3fgw3QwNmohvy1oT
rukFmEz9h+UnlEv/9bvuZKMfh02UILRkTrClVP2OQYToWMO+aZ8pjsjJuYR7ompx
JodiTBnuHyZmR10ecgUL2vNOs/GbZ6JpO4CZ5yWddvnTMXm/HyWhjWb5IEzT4PZa
UI+AgVoK2jLmxTYqxwDCX4Jw4ECrxzXYjJA5TATCheYtjdbqxI5iV7L6Svex+i9D
JugJUf63VjRGNLlKEp+ya9OvvPz64lyFceAr0hpBElTGjQoja79VFYUXsH0LJyyj
fuIb8i/N803qsFcLskKl1f8164EHAdYog7GEl6xWCvaEkJ+QxJ2WJMESs8HGYPVi
i/12qHtM1hK7g+JXDK+YXxtmA4RyJGZIhG6H+FbahIfF0phVE3Vq3Br+4RdJHAHd
tvmxfEsaXFk+WnS3KKj06ozIzVG1XbQ4jjopHZFsK7yh0FnEpWv6IgkFgffglsP5
hAsSGX6HQNdb/idtL2zy28FDmK+Bcq/mcPkqx60yO9zQaGUU1iFaxMc7TolwECCn
AOA+B4ltWyFqKFM3PLEEPQS9UPMN9Vc7uIuNMap+9IdY3N92asE5LBeAuQn7HYYj
2n2JpBwCdFTYw24hRJzu8/KX4oKy6g7zKLMvsMBZYdRqmneeN789bFYQpJV9s9sM
eD2S1uqW7sO5OSt0DRs70MrijsyhjywN09+mhaljQIAJ/tKPWVz6SftIhfUW+iG+
6310WlL/zWSWUmX5fgqNgtdOab3Wlo4WXJt91MQaeHezf+s+ZMnUcMyLChhH4TQ4
M/vZiVFEt2NN09yH3C7uYBzjFRx6FB5ELoh+d2ykY5IjK0ZRAxM6vKBTKC0jMIZp
vK/xu/kkJ6g12O9Mxn+7JYyWNbI8CwubOs27TjyA08nobp+toWEfprxVYvHanflq
uRSD8ZXfoW01asRTWQJDyoYlJJh7p0wyUC/ZRVS/QAdnsa0eCK91J17P6R7LYokH
8yaXvwnYFg859+mj5aFyvrztpRek+yx8r8NS6BeL2KBF0vF+l+QjgiloiSI5znG0
BJi6W1SMgME+F/spaHhLPnIZfPDUQGR5PUriGzNKAsTOpyj+TeHtKiCqv0AreCVk
k6XxK/8JZPA6HD5gwUR8EsLr+iIXJB+rS6S5bDsihixLmAlWKqpQLLDE4OWUhMnz
DofSG7URHhFIGt19P/2aDZMhVB/z/3OkLW04lnHmfBP2EgCG0wA3UwraFbqEjOTo
R/SXrmkYXy/27oOkkmrTYY2JwmFVVUwGQxmZj/aToieTCr4mMFkvfkIou1df6jT5
nNmT159oN1T0KeqGwFg8kTfAw6kivw47z/UECLUnzwTNbiGR/UoLfhcBv5kUC6Kp
35fe03iVkk8Ofl5Q9CU7gGRIGD1q+ae9b/kYQ7yein3F8z99LY/iqx/RA647njo0
6tgldDlWfHT8Nbv8rqOWmHKzlNQjc8D8xmL7egmvSHeIHNBXA904H+Bk88YuzL9X
CTc8Cuacz1nHFO7xtv5/2Os1sLSjIMfuKtbbmqEtlmw61BLr2jvsmisfbuuXDqO6
nR5eDdbxaM7MVb+UrfXFqyoVBPUFELsVxbUEuZEJLmeLdCsi7qY4ury+48T5QlSi
In1pP7rjsXOLrI7Ir4K2xUy1166x6aex7xnju+9KFxfsDlbzNbZOWLPPF/5bw8Bb
a4qo5pxJ7NUuPSfgVCRxE6dcL27/eJjvfSfb64uf/wslCHiwWGASc4yaRVYZDKn/
G4wigHEZkBCGBxfo24K7Ss/HwkLVDJa2qhtMPkwdhsg3uZIsbHOHGyez8Lq7NACJ
GBB8D9TCOocMnNEIJyHljqOwlwMc8IO/XYW/c9FNwxDRHGDEsQeD8W32pinJqVMu
tnAduyMOi9BM14U6AyhEh972nmjmcPjhigOdNCORxvVIIT52xIbEe/UpahSJf1jt
QGmLpZvugN6Ur8Wcf7XdfVUvfaxMSrOhKq14c1KqNe2Yvyt/vFjsIP1MQul/R48O
ueD9KgNZx97AkWPkOEXtM3IF7buhvo8XWWP01UQ649w2mCkQ67z8lwpwXoIzLiih
u3SpaqE89fxNk/JrdVsqgdjy2kVSR6E3IhFuOp0kOIeyypxEH9RSiu9hK+z5YjHu
owFcaJeBYgIKnqMq0Mo3Wr8Anxm6jOrFZvPgdIS/CuXxgUu4Z2PE5LmnFoxtiO5J
I1YX1qns+WcYQxS47caKX1BAmvsWSz85YBYiappfrj/ySWdBQ86zNRNqDDXoHuQV
7L1Oljvzb441wHPpUlNSXXi/ydCWprqo+3fFrYgI3ATVYw/SFzkSh6AYXbb2CysK
O3A4izXxbYYXq58McmAacV24b363rzKad7SraGtVoPoUkRVwyX4/z/JfYaIU9YVb
FeVPOApvD99YOq6FOkQdWxyFOi1Js8WmoURhcHNtZjUI6oX1fkAf+4Jzt922gGix
y7Zw5j0QTFJWKH/SrVYWV8RnXRvy8byanFfBO/hryww14g0QDrMuFJB4DSc5s/Tc
LoHDfgvtVEXRJQunlgnQfiLNncQL0zzvZ63HMwkJvwQoHFFydXlYGRcZoWkwTN3T
5jkkjbaxvCQe317rGbwqoN+BytZcTnu5/1bKOT/Sm+66QMpu9UdY/Yx3PA0qT4Yl
nUMgUd8zpxS2254r2knCD4ewxxYPtjj18wW7q8iEIaaabxkMSP9KmcRQhDgMy/DU
21a+ovcLfvuZsYvaKghaIfR2zCN8O4IeyIu/bEP6WFUH0mCvvzyt4p5T2JWpbUsi
bxlkTBVj6VNrzL9Mmvr7ZvWNp6LrM9cx12YjxgIig9BaUhKkQ4pEv3rACLWEw6kE
n1TI8WCyDTTLf7OhYeArQCYPUAZxUinBaDW21/NuA5zVrI3y2JjscHzOYWC0LkSX
XUUj2uUl6VpRnl6PW5KIBWtSTn87FXiR6YPK77h2WvhGN2DYhfiWedpUXsc8oEda
Gt6D2sASqxA20qK17GfLpUJS38JxA7rVQ3TyeQ9yq2AkRWX4l7d05rLH5NL2il6G
cXSUfL40hmO06vUvyG3YhgCedlc0quSdK45TnK2kgeWDuhH/auWjkuCnxLtDyZda
H+yO1QJOl+xi5O+opEEtFedEgm5AcX/qvkiBvRHdPt0QzXLsMwdcQJskWuZZRay2
xOo4ADiAgLfmWDtQrCxzVITf2FaT0WAQBoJFbcXXLCCH10tLpWtuLdjNhCjnxMJU
lSj+zxH63Ckax7oiOss7Oo2uGeEe38mHkvYGhG+u+OYG0bQ7JR00bTYb3aqgnORQ
9W/GOZmtE/9z24XDaPWHD/b4wJ3KMmjszBpmaSoC/euhDwpmUvi1awmcnT1mGb5G
Px9b2oaqHpHHGB8ShdJqsI5xKxppzVYg46RN0bEF1U0c5KjS9GIvbQfyeCrMkWE8
DtaM/1poHLyHzOXKuTWn+FzPquAICtJ5RqkTslymwQmPaIDXIzUdz+8jF0JjQbve
LehPd6DUZfqhIA6bmhVExCJp1QJXcRvTX1jl+B2IOjatVvImzh9Vi2I2pjqpGP+R
lbe+YF3IkehCVYkA5AVGNHp+I7p78rnBI0ifj9ujcIzrPy+LYR5qRmHLheWWjHwc
Q8i59vtBH8/QhWiCaRoSVrgUSohm8h+griotyxL2XVGB5aQdyddbC2JKm6uQrr2A
hSAl68aqCffjjUjj0eDrmYCbaV0kpM4w3GNX+fiJL+NPSqcczxabkCvsikWAylO3
KGJRP5agVg/JjNCSb5u+6yHqiDVOeC+RmT1fgZvng4kZtthiAAsYk3zDmyTwtf0n
ZysHxOvnG8OPmiWUKnJ16Y8qpA35DVrty4N5U8lK++pgimPJTDEqEjJsuEKgEyMo
qsZxlG/Px1Wdgimq0yHtQ9krmk06PXoPwZRogtp5OT38b91icOSaiDZk8CPVh421
k6YQTtEU1hEOkyeT7aVbcMuuJJMg2HHUSfTKuQFMkfl6q55HVI6jdCBWnriuIhss
JidyGQdk9kSkocOGJhUM4P+MRZgusfFM1NcV8wi+0XRIbGIveijHfSuo3e7IvJ3g
fBVCYdF1pfXo6ZPkIECBvJtR4dAZEKXXujNgX0jbwXZjOdEo/9m9FM5CIvoGOhwV
x4G6OqIDBiPP815nANYOri5K6CeDJsfCcg3JH+fdAuXqe5/DsMxQG6xIQJnmccMa
9NzQzD3iRZ/BPtJmdCjzMjVP+r93EaYSsnABUHgBlxgXSY0xmRUSTHbNak/4SR8g
Ndz4VxVoKTgOXKOdfj7Ptn8kkOGct82807q9LcpOtTtsdi8LiY/K6QO/M+rup5FE
/rwHVmOnVcHrvUMOzj9C8wzB7rdiwIEhxGz207YezzoHb01M4mkJ0umFkQzeEzSJ
lrmwKFjSlJCEaJuSK7BbUV8r3fl4gm7rgMIw7lBOPTPj1QZtdlsvF9xxNsi8f/qQ
Z2zKdSt0+CqXVASNqUkTrGToYNSa+Wxg3pP2COevPhqwxW+TZidiSAsskt0sd9g/
fFON8uoN6aDLqAby261WmABVSUxSY2l/WI40JZv2AFuP92En2/Cd0FCKgho9jXyi
Pz4tevAY13AKR+oXoj8BhgoMz3sQi/UCMh4BP9jOdOw3j/KqS9uRFkytndI3Ibak
oqmYoZAfpNca+qtKZ5aqRHEPvewQ/0LnGNQVI455qEp1jhz7yizsctgsXWtEl0RX
ZQF/sfVWTUDKIZM7MaycYg8hi2d2ZWbHDg8sJNrWIu8MVQG9CWL7M+C9Wkb0Op9a
ZFLI0WCTupfY2k9b2UpN/G5PETEMjornDDI6qLR582RpSpXxaIVFNjIE/eCV3la6
uR/ZqlBh2vMbCTtsscdwKowKmzK8lGiPFsyBzm9+RlXSY4UCkGmNtQpIM87eSTnx
MU7Ww60CVIIlakz/UOilRlg9TXqHeu2HZts7bGRevmEO0BdvpePoFcAOr5e0TVZh
XfoawMTR87OqVN/BnmjOGBGegSlVBcAdVsJ+R3/LUlWk2Y5F1XShBrsmP6RehbuT
RAp7vz3uNpd1zVGKblNwfUW2WQjTdzxY+onB1TSMSSBsWnnnL/TEtlpWaRwb3c1N
RVsYQeB3uGyhiEwXrnDkqU1mt1PT41tj+8gUL8IIkB9goARsuquA0sSKqlYke6bW
mNFUOaMpWlP9RQ2axaG3MYUo3lUK2FqJGcn24Ryuz2AunfA2ZB1Be4b0Cx/RrXdz
S88WmZ96khkayIg8KT41XXI7tmZDTo32OVsJstfOpPifn5CmlbnXpfs70ZXIhX/e
eUqqWLMMSwrIK3WdxJh7n7x9RXYWOktgR56nMLtYdARmxHAFduUHqNNTvbKCyiH1
VTi18r02t7jdpduU1BcBQ8KMhlHqh6/AptWQVPv6StnqkRjXXLHhv0zAxkro0S9c
zAuNM6Vs6DIeyNS32CLH1G0/9qckdZR/twIZVDaUEzbRXDz5LLx5PGSYN8Ib2bBN
CTPHj4ZoIatj2DWMIfe8MeHnCCst2w+XlckRx2FxxrnKR0FHaIeuulwA83cMw5/3
K/tzUc5sxFOfQjNFAUhnk522WHNMW4F5ltXaCqJHzdfft/XfSH3n/oG4AHkaaY93
EsiqQGmnDd5gXzBx6Y3EKQ8dVB8W/RflY0CnY1ZocuVyqkB/nqtHT8L7qoA9dcif
1hXg/2IOe7g97OMNFA+9q6EGG9eFVZhzgOPp6c4DCpKUuRGh/vLsUSzxnkjcAyS3
aB9q7Rpvgvf7r6goilNYZaYiTYcmYJQD23DfInAQObbUyMBK+oHhfubZxTvr+uun
N+R+h/ixmNoWKYzx4VGpn0cVAO9oTrs8VXnxttSZyppKgJ/w0GSsSWOGU8Bxvd07
I1lFVGMdmoT4zoQpVkCog96wXSXYsyfC7b+zXNk434k5mPgZJTMY8h/32s0zsPFf
MMf3Sow/P4YjSOB6JjinBRmzw0ELWc0d3FlwLfcROn2QqQPW7MKIxnV1Fo4tvrdY
tK/VrOxiWO7Z1lDPskEZCEOQitXiehnPHl+g+6yXEMftm3sze/am/BEnAN2R1Kp8
Zi+xJ9q9V+qiz1GQ3zu2N5Dc89qMKORjMiLM0U6IAFU/0U66Axkdto+9zmP9Fp11
jrcj9iCmOqO48Y3K3yu7Y2rHCQpc+CuOUsO+gbB5PWfkR66Hxip0LP/nWvO8h1NR
hnj22nV90FS1xVB40goHqx4Q1qSmIiK7UYfUWJITPxTMaZBTeNFyEFuq3C44SQQ1
oJN+uy0MUeFfvim4zlujO/HIyKzhwHIZ1K5/XuQ1f2IDswewSBd7hzaWUQK2JByc
9fjC3re9PjfyN+/PLVvh7qShDk6c4VCRhLQVPVTtXbJcB0W12VYcndUoLCdb8Z4N
uSBgZgIzPNNfVLXIVsglSpCEQI6ht3s1ioumD4Tpp4EWI2XBYIUdgxnkjDa+M+lo
IuAdtaFCMpDaWjxVnIUb6tSqGyyLBZlUihaa2nIg62S0lFeMp0KJmyEB2p0/Rw4H
X6vyBlZVszrrVuAErb+Zk4pe/eOzusIuFizi9Im0PgX286bIbIMjj3KUvFiTRvlq
6gHotIdfEDbDBNM1otXeKJJjKEIFMRrxqrOEEdsXf96Q+ZcUaiH6cVuDSrvjzIcj
uFvvJwkr8lio6ysMhAFcrFGdFglWPeG7lOsdMG+k4hvvyn0NUmvt3Z/o1DkH2wPz
L1RMx9jaVSsJUAp9LgKOGAaIURz5Ae3R+FQoDgHJv+VpU+mQ65KQ3mNUBW09ZU3G
cowTeStGBm8xxPak5LlXBFsdxcLrNL7M5zz+71ALSnDjQ11+uVDEHfYHMbd/7Myt
pVc6r/rIZQ0aw/PmDnfHaPbSkAo8+wnWi8Y2Oo4loyJesKEvToBKA9wJgXHenMhY
SJLZpy1za/tqByR7Qo9Jd0PPtrhXbuC+Ei/raYG8geoe/qLtEYaeqdsJcqFAiEPJ
8JBCEXO/g5SfL9LukAtjIJA08c8CVfU1WfLfttU4Tj6BGfXVWTiUhKIfFClW5yZs
7EY12n0p1N8C2OqO/B/gesAa9zkejoU/lBMLytMFD3tMm+yiyDTl7ZP6DWFx4Z1U
qScQ4HECkg/p/GkC0QGHd80NWTBOWHcnsifePCkZBY1On09dLzrDQdf8TPlWVYcm
AyLXgZNj5ruWF2ninkl+fJs4TzV/XLXACNSEPYToRcrjcVOOqDdTZ+4OTq3caZWK
mj7NGxUNwUI1K4tRC7mK53DYwyaGzfmwqZIylF2+IIOM2a8PmvoAG0VocDqhzgQD
4tEFdmv2sdV2+cfnoLcFN4fyXjzTH6hDiLUIs3qZe4zP3D2JcPEovv6BYcj3YUJR
2Ng2Dwjy58Yt4dFrMU6HFQzvlO3tDfQFBRZTgrxrE1gu326Lf2ynyqBARoWUVUJw
rtD/j30baOBvVCiSWaTGATU4klRb00J1Qu/6WN7aCwzjwB1Z1OEBgldtYk3EGdXL
r74zPtaXLvkBANWnB5Z4CVHArzPR/GVWatSD4+g6QtXwb7OyFYkCaxHQ6YXZgYKH
25fXTLVM/KxR7+DEFh7yZWbcpm8EVet/piWV0V/QcCoTciV1ZuBPh8U8VUjNppdW
ldahETODB6Y5Yc/LANIaTmqE6t3wHmXgBBJuXKrSWStv2yuTcUjybaDLv7SDw/mW
tWPy/Hlbw463QhxbYUrVHJVfeo2+IAOCWDpy0zSO1+uGG3APYxkp59n1m2P3GOVH
cTg/QhFcuc1Bi18INk5NdRKGG7APnXqpvhVjinNNWlpNrK9W/DX0JujifAU2I1yu
HcPgoIijHiV0f3tKfts2gnItqPVmJcIeGZT5vTcCgjlTB+BpKm3+FjdWTTI81odG
prm5ux0iBFxyWB8tx2YHMKl8Yj6QtMNiYkNMoNg5MXPAtBga0D5bihcAs8K2fTx8
tsRHRTXEKIJ/4b9iKmC7d3dX8g0k4UNtXjbAF+NA2QIs9w8b6sziGU1BTEqumTz1
0dwdFNSs50yup1N11D+V2WGH60YtOgW2qkE88P0ovg1X5ZfWZn1YOtIF8zEjeDd+
z9u8m5tk2qwWHT1SzcMNDjTVeR/T/kVcXYA7jYf3TLjFxXgM/7YASwPFjSp+O46E
6N0SHQGhgC4H7ABsLJQlZ7xjMKEmlh0B34zL+X47uVCqY8epwBy1yZblPxt8pnna
WBouv473bHOQ0xYw8nxiwgYA4nna8hfvLXAlGROYxGV2TtrMzycG2V59er4lCg8J
hctvq9V5js4LCgw8mX0izCN6JLKSXtAPM+VmVxypAQeD7+Bs1Rr79fsMQVD7FCGs
mP7JsU1Uh+n/PkjGRboDKtMfcSc4nSANNepqw3K/wvzIXrjPVZHvq13KKeY58vQt
VRVFtNXQzjm+bj2yIPe8IzFV/cvBLlI1nmQzWpJSzME1o3ZRm/Xg5/D6BGiXqxWi
d/pUX+2P06Q2NC4C8jY8fLsAgFxbCWtBzyXko+k+6N95wDGw9bbyzJgD7OG2Rvz/
TXYz2N7yowj53tnNU1K8ppxOlq4bRnqjVYPGuVVTwTt2GtRRqnk/3QzvWt8PRrxf
hSSHoH+okjYOHRJsD/0LBXVXIbxAvAAFsmBgURmSvde7IgaFD5EJkCnrvsl1fz1l
Ur5HR3Yf5Ku6WLXpAX22rDpSVTZ9YnZ0B6R/rePFwMJfVV5TUG25jC4hhL4MTMTy
zqVfD2iWypaK1LnF8cwGZzv4cWXcmt7u3hqllSJit8Dq7b+ee/49UTQ5rle+qvoZ
p3bQkp3009SUJJ53/brmzs1fqjK0KVLJvH/dNHwc4oz78zkPQzDfMutlacACbmGX
ACYpRz7L2EwDOt2NvSWAJgdIoJh79DM13H3g6nCWd3oRokRN3oYJKXP/VNjt0mVg
+bAR+IKtG1+poZQBab+8PRJ2CPTs8KhEW/I2hR9T2bsY0nQ99iUr5vcdogBOMQ4Q
iwyNeWos/h5OL1VWiRayi068eS6Bw6EfIXK3PGutUVkZf43mS4CFU0U393fXbIFN
AzKqJsIT2g0qopqBpUf2pcboijP0yH88zdVDth+k8l2uQEeXyFVeC2kr29fOePbS
Fs8a+Zm/pp6sdp6+ZCjtxk2ZJntqo04PF5Wr5QUo1MtWrcOEMo1/4wBqdgLNjxaL
NoyY81HE8QC6VmC1qD3alppUvWuN3w5vUwkY8lWI01kPivLagaijx4OteI5hjS2A
t1cLgUO3QHXNWTbjRg2TJHJksG0G+njtk6Vz7Qv21zeLkVDKTecsccmP8oddgKAr
i9RVTzWDP/rhrHDBnlyGKf7cQ3h60HNor5Wo8F3V2FrnoIwMMLAGd6QSnMuWmfmO
k2dQvuP0M0YYKWagZ4hRA9jHUCbXiguGzgNrEKSMV88r3O37fnwfEQJ6fIlDf08I
50ZDoQoqjS4L6EpEAX9HITnsoNDfkOy8eB4m9X5Hc4c1lDcl+dUwLnr70mts1vPB
E2K8Feza+U0cQeE8Oe1cU5TnQxiFLG8uDOTJ5BjmLaOooHeDW/xwZXs05BLyiJWi
WbwUK9xFvoljg1WQ5aiJO6qyNsgbkDp+89Pl5tiGUpyrylRbPnlE3j+ENmNZY9Nv
x/5ivrkGw/PQKKSQL8KMAjf94Dmu1tPIMZIA9pcdCIjs4M+SICeOxtlhTXLbIrBG
lkNk15RglzQF4Qu628v/Vm7Xt1DJPQBeEfFynRDK6uq4s4mYbmWWFCHE3DFheoA1
em65B1G+e5Mbu3n0AnOvmL4EhdFJoqIyKWpZylNxGog+BCWNyh8eFlmpqqbR+snA
ANJTCQ09EFxzziZVMWb34bz4+hROHBECzjymgw/gxaPzgVa/Tn7QVtSo5E0oGZxB
u1VPr8OeemN2autURh3Tp3VEiRuL/ep07uh7UjFxhg3N2lJO1+S9FUb9jKhQh4tW
RadbbH9pHV7413FJhezt8QYXMqkKkIKNa9xgvz9W95AOmRYi9rWTXCaqzRExpEMw
YSwHA77huwAacygpMflFMeB+g9ZvghXDrzdRZAqUuA02KDKS6oLzsFdl9x6QFjek
PVlNPsKqGtJf5lvZ2q1Ed6PNC4cHcApVOBCpIeJV/dhFH3GSjLQABPO61CiA6JAm
zN1V4R7lA5LUhYulh0exM5KmXGskpIyZA9+ERHycGYagGzPNa4a9pfM8omkElUzA
wq72Jy/ZqmZQv/Tnd6vWgAJwDyZBxm3gD4fVZoMRdTgDBcgjHFCHEoDPu029a0bU
w3/FDzyv5hRhDH/fH+Vz+neO1mnnAlLZa10keZMn6i/Dn63qSJ5CXnXWuwpcFdgm
bU++79rHQcxlzCOhIdt0X9KG1F8YAiP9T1IEUy9HkRs4knXoyMvo58NjALOFQ1Bg
k7cVubcVJXS7LP6KGw79eVH/X/nwAbH3ft4UeyDbCWgNO3YR7C58mcl0uure59LA
Cn/XDYRNiM3FxjSrHZ/4T0d/3WctvM3kTop1EBUSrL0I+43PD3fIj8d+GZNE7wKO
dSyzcvEG9nA8ReEJlNht0+kDc+R1+m1cEL/okjfjlwbdzFqkX9CB+R2KR9CJ71vi
vQGq10lR5ZWAR6kQuAvBxr1zgBQzORnf9+FMgyIeSdgbTN3p1gnVbsGmsctLAvu5
DEwLXxVCMPH8u+4JwQH0iK7ExmZXzwgKtt8K3WDU95ibXA0XGqP2PxhgADhH3J6z
qjamSgEcaIKzZIxElCZUVu2NPVsvYBBUGs/GJEjo1Qn9jGOKBgjFHltHsOemXlQV
4A1JJLtv2mbHy6gTva5k7sh30h8+7RPHD3sv4BNZE6RLSi0JmoAG0jSD9SkLBaAK
AcaYJcNd2kayA/yJtqVPUYM1W9TGoWOY1lf43cYOTpxxLVieyRhw8tez05hyzggc
Y0ZHihrOA18k0Un6pEU3CPYoQt0A/kIOYrIs00nD2JaNjr/9jiVPfbOmN4+9aUUL
jjPIJWCMreG6mE997BMbdhOWRfPwhaVISh0cM901C/hNPo9r2JWUsZW6iMokfzE4
+Uz08KZ2sxOu2zyePMBSuUHuo/5NGufsL0xYg6MxtnXsa+wXiFbc56DdXIZxPuth
59Yomk54dOFMGw8Vbk23Mi3kU8mf6cvKcJa7UghaEqS0dYLuRqFR7QPDNlvbfdgx
4Lu58dFfsQB2s4Wm1by222LUvDxTHb4yDe8AywxD6PiPzTD3TY7PjOz+2oJof9cy
VVlQa4nDYW0v0BcT+/+oWR3PBxnnFIuiRfH1hHe0Eosv+oksaYITmu5WjXqJETbE
t4ZTkBthhvhZo4YmFmhddAVt8jRGytiX8gVjAK/VQDUmB/eLDnPenhnVD/XurdeT
5SCa5t68STREILq4//1yreQX4Ef3gmAf3o4d8UYMHnSyU2nHloaBYYrKqDR7cYrS
HxkQB7x2kqLCwrrHkw47LEIFlq/zZt+b1l5wkkn2n44TLggay8g66pB0/oP0YEcy
7W/nusKm9d9h/kELMVw2loURt5wEznZ/eav9mzueFKys7NU20M1Z8mSDgLfz5G8G
JQmbjbmAZwgbIY3fCCUMG/jlUBpK+GuojqNR3G5yCTMywdoXeQ0ai5V6d+UOlcbx
cDjmzmvwUhKoHsNCejI+zf3zzFM5Mcn5nOm1IiEBBHE9HpzvXZveZZDJsOIOWtUv
fiyl2dpNCCxXdy59cMZFwrRwI/2mOaU8US+GJdOyyOkrbGoREZA2Cmm203faZnP/
X49PV3nc7jBkDP5Fe/U58aKlH76www4t7SnivstoUCu58kDGRYVNvhvHVLdro41X
vyNFVYe4t058GHOFeApki3JzladYp90rEbwOUgCua/zIUIMxfLq/ZzDXv7b6uIaE
UG0m+GmD5l6iCPelfw0j3tohgse0XPI8wzCFJY8lQzkvSP2UIWZ7PoyoDDS5WIyU
Vdh3EFKRpt+ZN0w0r3r0RrWiD1W3bArQr2LDNsvK89Qn2Vtzh4ga+OwRVW/N+Kio
fuQs4wICB5Z6AStA4bvy0WIZX53lcnxIb4h1rRi/YpuPWZZhMCuXHC8MB08HINLR
aH8z7X8DZrqpqli4uL7VolYtxYHP3hnHG6L9dF3gdbUgRKUa15kBW5u5hOJSIPoc
dr6aKXNH7wItUYEB7Otr0a6rTCnQJTfkAMTGI/3rZQfkZddJSi3eJROokaKB9QGv
Pp2kHDjbnod9m0aXO3qmocnHI8eo3hujrVnqPiwRl5/c2/uuxCm/W5t9of7KfrcD
BzOa4BchHVsPi1P1Otv7Ao8J/OKh/TdbVjyDLhgT707SggAfOCFQ5tgAenIpDtfE
8aC/v9REtsyw+Kh8cY5BnzxW0Hf9BgZvY/YM3ktYVWcWyrV3ApMFQ4EKwhyuVKdX
ZZt5vh1pMOASlpi9FEuVuq5FI+Y75tqln/hNk+ylLEgnwDXN/EtPU2lgSboGd3wC
+iv5e/WS3aD1GeIy2dYIZAESiBh7gR1kXEgAojM3bKCvJAJ02Ts//yw6gkPhAvhT
6mibvwbAeJ3BM+58AnlBrl2ZL5nr6l4hJMoKdts8Bovl/YqnxGBJ83/RWb4tyE9u
LHytqaYRQXy8axbwtdM1UR7tjIM/mkjx3h/tMzHK3nIwjikb45XP2G8a1lPBIWKY
x/0VxN4Fz1v3MeTq2Y33k0x9LsGCT2tQP2zAJ76Mb74JGX5TVqYwEnstR/u9GGS/
+DWW9d3woNZMAa0HVZI36jpqK2VJfWC0uCweCHrImWqilLxuj4QL7sp58UhBnGff
uj4dexgi4Pv1bMcH7/TBewrPUshYrc3Fst26XasJdrKJ6s8xdUwc1YXPOX+jpH6I
s4uS3Gm084msBVClXyXUgwGhoC63prwNnUsyjK6rqFcQY9k15FdgVoGsoicUvmGe
rmrQ2VAg3zCjA4BJqOoN9tnubrwW1twy11djC/X7dyyBfPAX62yGge1oTwHy177E
ub2gOaB/HhYFgqW90ZAJExdBwZeUjrEtu/P4J9Yix9VyiDDuutwg9OtniKi5kcDm
c/iNzUU2KblQiURNHDryw4O4eZFX8ATvxqqkliUedKr6EgJqODwrj0IwnKq3wzLF
+l4ZLX8Bn3ZfqnLBl4r8nRIgKmcHqLZbKC82pZDUCTTbGAgGgsSpSYItDglOGHdb
cbIebZ7Iqbt4hro5LikiFvwzvpVbY4SQkPWncaxY5TrgdMqiXwmlbzRKcAMobPS9
LzbMpLRuTtperTwmIEC3kFuEDw6o0g7pfD/J646/UFeTcpgTM70rgpjmiGbUYJem
T5vrXw38dk8olyId3sz93VT8ZfdYsSq9reuUXZMET5e3ugtho5CMmWaoRHPkhhyZ
OH60iXmWIng/VwSCNXIfKTiZtpaiRYiQKIGBGF2uK4a1TTZZrLb3fvdEg28WISXY
tgOxMWWnC/xWvOGxGLSX7dzk5HjTnD4cWykznUhnKYxUwGhr3RuUv3D3OWs17/J5
gWy72WuozUpMTUit6nGLzU5XWptWvFcNDT5K8zRxSPw0KSjeHkGb65edyX1FN1TK
ebzsSK1SOkWYTJJRoC0tJo6wVsZBpD+aBQMNK+GUHIU6SJhRVu1e12dsf5Nw17b+
EX2f9x8n+nDmvZtW1aAyHVO46bLHD98eeUU1OHCVM8AfPIsjx9GYisaiQHg1C7VC
N+i2FdJyxb0kwDESl2VxPGWbFKTPzF1crYlr8SmRx0R+lkrJbH+siTaUegJHr1Ph
ki4ZBGRmSl/awxvkAXQgqJ4sqgx4R+vcEepwUMmoXxkC6Bmg8JHjFzL1MkX5H94o
5+tfznOM9/AUNQPaAGin8C3PooM/SWUSy/xfItQwik0QL+5jd/MJL8IG8BureZFk
hmdbtWfm+8rwIBC2YRLfYjrqBr4viO9mCqpJ97gExhOrLyKhrsja0hncPJU5pu2H
cYR7ZAzXhwAJTwGFK6KewoqlBn0FZDVnSUOdHzm9z8g9tKEOVedDJ1X3UymqH+4y
Z1yiBCmEa7Fas0+7DyGoyqswPRo6lrYNB7ntce3MWl+jhyEdHhaeMi9sziWG/XfV
mc4nHzc1wV0ZzGtM2uXXzYFvxgRNMkxL9gm/9EddNrGJCPboH/RvZeyRi0x0GKFH
NglaJAyOAv73jCCI0csqEcdKNqLZCha5DhrcjDvQXXouiBHO6Mw6EUFdjq6Ll8Iq
yzDpjTAMeMxEg6oVP9Fm50znc1f08IMWWapXClZneZG74wVZNLUpqZfZ047wB/FY
mdPmvpxEZOxRtkMOafbGPk57scdRhyFIiO0jlDdr8ljAvlDM7ZBJNbG0YL4JE/1t
28FTt82+QDJrFJVfMPBPBHBtGCOwwd7J+IH4aAWVBVqI4g5ijKkO6P4T/DedoOxE
I2fqDbM4Cf+QQ2CdsZcx0BPA61M0LuHThDISZmnHfjgSmaxNfN1xMAJn90SLDAx8
KJ803vsRoDyRgo6zC0O+qRtVQW+lbAR/IZbkVegOtUQE0qNtpfOrO/c6hjV5SPAZ
4A4jq/lhN5yxy9Tb8f4Bsk42cdmykN5vZunZDB4HtXSEBk71jE+jAv9CyCZODUfh
HfNA0lOOR75jmWTzYxCDqIRI8UMaGh2Kcwjdin921IfiS34SbfiN7qdmOemMfkpw
Pw7/XChzEidbnizKnAAwATqDQOvF9HsBOwaXFZrbotltDp/tJHIwcR+yek1wiKvB
0YzYe8fRjaMohl5VfQXAZuV/yS99yLPtqImue1jEL2yTrNPXnkd4G/MlGXChqql2
qb6Gm3+ITVXs7aFwYzEElVm0HalbOC8cSErjMEs5a2vk6O7UgPT2bUAcG1H3bFbg
Hobf+9XRzkEd/vOwdHGHKDbB7bs48lXxhZm829tew6R3DvD6SGgWbMg3ZOGNaK5k
9SRknKHMzxRKfRm6FkaYUGUSPTD9RlYNOkFFCtixFWCF992R5QMkpLNTJ6vJeH+N
OlCnHbNoqP2Mi3epr/e/ro59VLyUpcTuciT9b9KPkjsmjejxW28Gv/gidUdsZT5F
/CsdfnOsOrUG8OdM4xPAdwTReWnJCY3AvDVEgmSqzCXAcQ8JvpSGxnlQ4dF/qv6n
DuDnWnb0a+D+pEpZk9VH/CurglvMfxu4puG9ZH7rGVkki8rUJZLvzscN1/Ry8xHJ
kD3x1fJCJGmgSk6aQOyrM+jXYpa0aDzdRaZd4B7Jhwl9mZY+wofkwdlN9OcC0qZl
BfmpckPuXuUZFTAbej0Zp9l355PSgnhA48GO764s27Ekqj7+5fiVrDOWtcsqLmNc
zK/x0hRHsnh5iIIIkZOYPH7PFKpF3iuIGTphAFwC6eO/FZv75tG/FUvgq39r2+vJ
zxXy87GiI1sBd6gmf/gWysUKvKXMRskbjOhF9CiQdGfmOoaEMR93Nbq0s8kzoBEr
wpvFULMIgnStltwTvNaWQMVbO/svy6+AwoYLGQDHY1yIGd8uAZIfEbG4ki+sU+wo
WJFN8fDF4blt2RUYTDWwdQZBDb2glvQcj6Nt6A3+5hoThX/ImATF6BXcN/Z78c7d
st2y5EoJ9G0vb/AxCCpIIPnzipKir+6gXpY76uSjqqkG6cfN0VaC0QNa1L2HPffH
pGrvwYrG6z491UJdntHWyjJhkP+DyfLMqdPyNDrSTD4NG9tSVvJfL+7eB3Ka/phw
dYLvHesWXMV2OUVAcwc5J/8+0/5Gujo5KDQ0uCJ+J6ORLwgJ77JOWbe3x83VfQT2
vGfnAjwVdjucUS1Qz2cDTGqllYZc8/0It18nJVHApRNV2IcDI2Tzo9W6qlsrzwks
cdfwMQ+JYhCBBJrkOvEH+q+OHKl3svlJAWiIq7KB05hqP08ppMiTkt4FS0A7FUBa
FzmApmWeXsySJZk9LlUyJDIu64w/81DsL/dPhhR6vs0lDrSj9hNhwZwvumgWNu7N
VtlsTW3sCJuShAqaEPLCfmrMKlmVxdtWEu54cGzC0sawZveJMJNxVxEJiVjCjQYK
H6hyY3KqvbC6MvBb9x1lNEmExroZDlEA0Va4hMzE+FLDfO3RMo+dTaXZg06+ofDH
ACwPLm32MEe3WuxK9IlOD4TTxPXv05sz11wtHWRByZ8XEI9hsw2psAEcsvLV5AUu
4ATLeW+6jCSQVgV3pdBJ9vWDcbXt37gtkGJTVV1YiOyGsSXvn9MRrHGcdMkVYwLL
uIaFO+0+//fpzI+TuHtD/XHDpet/FuptQlWFZQpBDCqxrM9Fwo+DrMVQRYA54aC6
uOEMj7uGUeGW1gvIMYkK4DjcfdJ4Drgb0BuUD4/oaNMMv0DKbXSs1E+CHDIsYn0o
Tql9DZUwPRrqq3m993ke9o/+HHtwpGcAUUA9yXeoVzWvUUmBZgjFW6/uGA+zLYuM
TrYviR+xGNvN52pZdKUQfG4R+MrO7II2svL9WQDXbCx8ljNVf8OVZGFyaRi1yIDv
DGkvln4Scya2ZpnyuxHK8HSYSlrzFU99r6M0g7c8S2QlFLOj87yfMzDuQHAKBUX2
awHrwxazcgsjfHtAlH4AubqTI6fyfiJPxLzu6rGaHJuCBNXHrehLfUMIvgNj55UC
/FuvUDRqzU3yzKOMuKdwiRJIvKAyDaq1bqGQZOcpT485HYSO0QqSqLuwh7HMJQOW
zoGCnpAQFXidY67cocKClh/cz+gFe9CWdIz4Qb+0iSmDqvrm3fCxkgw2iE9Vfv96
bLUOFLlUfyLYmhN4rw/e6P/U4KSHefWbtStAMEzMFZGiQ+12RePNHLclgE+OTl13
42DIchTB/B5FQqm+3S64J7SxzSW7Hq78n8lPDMalKK43x7bZCbLlQMVfSWKuggGZ
m+IDZm6g787g3eTPXg98LoiEy1bNcduTNhuDRNbYGef/JLfioOtG4fRDyb/m/gs/
wrPHFblp+JTQbjE7b8njnvNxzCBg7bFi6DY6Vi9mb67YYajsn9UdZYxk5IccUG8Z
3UHMR/iz0HbFOu10fp7u0v2zpJwYtCXLAi/3OB3bqZfgyK/kOiQgqjaMF3wcaRht
WCsgQn6z2WFhMM4Hr/8CM8T51uCDW+qn+lYiWaHolGWgK5z1/oPOZG8Qs1MgNwAc
5jghI6FRxPWdIec3WLWzTUzAwf6ZzXDMv0ZVCnup3yDP095kv6BQla3txinM9Eq1
oPBPMjQftJ4DEi3de5B6CODtrWDFLVUgN7wIgR1ldqyF4yt2v8IAizPnaYO22dAj
282Gzd6S9MX0hvIlNmv0bY1mdAVLwnP3zRgWk7Nx5GyCQxLnVpwDl91YxvsOyqwu
RhHoAEb1obZrXu7lr80l+XfrdO6Xt+TF8HNuwfxTlS/ssgdkujvZ0Y+XxGXyibB9
29ZbwDVHa6tBRvRO2Y6cSA1zE1LSdloys0J2GpEm79IjdKG/gmV7uaa70ogQdLId
GdLwy1rK+zyQgW8PUaUKd0KrXXKYuM+S1oxEb1GR0hkIS5YvxHjkJxDiZKap4Qgv
9QvewDX7iOE5/aM4ZELk+PcyeR4JkYQPIr9ODxSeSS0DfebiYXNhBCeK7YLUwCbc
9AqYdSDAdPzK88kGZyIdvRxk8qraBkFd6QS5uZ4Ykus5dDrv2ZI0UuMeaQKzIGP+
lF+GHTSPu+Dw5mWljYzqFV6cettI31ILFKkq472gNetjVKEc8mMjFXbImnPfvE73
HqZvEfcTajYXxYIhb2pwsC+bZvb3d+4oB7wHt2FXUiX9OMHI1uFpXzFPycRb+H6S
ta8cXdlNxE+huJw0DmqzNfq6Jqvx+x7yTZU4ivHtL0pvlArPg77IF52+i6Nu9PW7
mylJMuNsBwd1koqCn0hcKzL4sGMFmY8wab9sJAGA4H0ZvfupiF75donRbok2ykcN
oDD8ISbYKVhJFydP1T5nF+VWg654tpZWukfJvuuM9Oz7hXXjnycSnGyIty5TAVDl
kg8jfY5RjzbYJ/dKcMdRfMKxNoH0Y8DmtmpeW0zUCip1/xdIMM3symCXUH8wjrP1
eNX4j3x57mfQhEdls7NPCpNFhuDViHzwGYLA2pbDeTWYK0DG6OvAMWFOZXt606ge
XxP7bLPXiGepbA0PDwJggsCv4ptB7aE/PeC9Fd0l9SjCU3bLWQNwpW43eOFH6IE8
8QuV+jWKpg6H7ZPHWBr+obVveeadtZm6rPmHAHVjnTG8pV6Lk86JAU0gLCsl79TY
pSvemUCDTSys4B5ZKVs5dpJDtbI/TDSxJGJBl48e8IrIQQ2ejohugCOpgyhMIgzA
KKfpYzyW+Ssp/662AkTyaV6xjPY2qEWLpvrxGRdtrwu0qnF3H6HErQZajf0u0ZY5
8weRk4Lw4wHv9y306X6h98ZUcUCybX3+J4DO0PVN09iqcgF50YqlSqc1vF6NQXJ4
C+DpAMkQQHoos+BSrkJ5y24ozuPOvBQ+v68yvP55yVJxjAtyc+/ptBlFlQoj/SBC
hMmv4Z/TLJapVBv+A1/Evk505PW5Mgv7cuXs1R+917+PQT/CHmBihUKWkC9K7Cju
0VClfrHaJQ/1etByLuqqYALrC7DzZe2Yta8QfuHlsNM4C0Yzn8J+OKAxcrXS1a9k
SzaOV5ct9oWUYQiLdZMSiFR+gWLFB82FBVeVgTczjm8vVjmmWeq918/5R/Vw/jTo
OAiqwzhC2tVuDEtklx/LawfpCzO4Vuz288qOB/o4geJOPbP6Vl2EikBo7yt7WYE/
+5VBnlac7ewnAzcqHHnkrJmwkN+zR7Dw3tsQg5u460kDx9HJPLwkKVrJGztJUXFU
uXNm86bhkDNh6PdybVqow/dy6Ju52XpUaJhs4c68jY+2p7H3CgeOrQg8PpTK4S4N
b20cFeEBwQZfbG0hjW3zZ5vWM/7zNNTBziGTHyfgGl1DmgpTJSfq9Kol7nhIDaPD
O0YbcIeq3p6zTgiATjDKWMA9MrXG3R0xVdhUodMLbELpYAIGiMWVMbvsxk//jytt
G7AoEhIv4cJbHC0ZkgRn17ScJdnNgDd8AYdMBl1UXdKW/tcFzf+e5nG4648SBIsu
xI+cWQtmu8SFa3czd+M16QzLGk9cEcWrUvT5OutRpXLeRVrEdU/RKly4pQU4FsGg
G+1IN2Wq4yIh8yhgxbpwTAFfbcPm925CCfejCEs0UULZThpH/vTuyqpykKUi2yrC
NXRXDw6fG9HmTeGedlWC3TeL/0VbmF+e9vAOAz9HpgXmcrhL1U+dp8GwFlLtKU84
cL5eH2EcrqnmIO99OHtrvgzZ1CRE/fXRvSUV2Hfh4NZA5CAR6rXaCnGcWFbMcNXW
rBxginbC8aIBCtlPmx4FBz5XvkG/lrMnpPsGsY/36zAdJddkP2Jifw9Wo+pfPGTW
UHpJ6wgnYUKh2vRt/vByd7aKEf9RCDfPXsH83rrTIlBPustbzIG2h1pMsys2CbXk
zmwc5Jb7STCrjIQIPADgdgl6YQRzt26LbPRj8LYZG0q9v/cSe/PUjsxWusGqnzxj
q+CIzWeAFsQPJ1+ZQkT/y194RZhQIZzwblMPCiXZ5D1WLzTJLREHJessyuzYSb3o
VttY3FA6gPb2fl9OtCdjk2RTF2mgNebT2Id5v/3zfGBfuGdzHBA4s8i32axGrb7Z
wtvIfwEanhVTWZen2M3Ul82fhwo5x3SfhzgRzZFg2HOYubMSF4BqXySP9822EuDQ
uXPDH0jKgJStKcBWtySf6Rzm56BztDIGyyUtwpQ24z2h6at/YSUlpRr+eOWft5an
KDGey7KLqio95oX74DlWrLwUp7/bQDM4v2hOx6idh2G+EQlIsClyOdvMa2eqwMQK
iWsg9drKZTNIoQJ4kvOiYB4k1c+kI3VDQ8ajBJOWPcVXXQVSX/iNNRHdL96bAaSs
6eqBbm274jUyMQAvLcW2CYyv73nMp8sBwY5md+d4F2c2E48DQ0ML3mPof5hNi3mq
UkiL81iPdOaBcPnSPVpnU0yxQZJDMtzR95vFBnRVzmEHq/mPREvjSMRhGvtKcYm0
TkRhWx2xu1yVXxcP3tvEa4WKy04j1j8FQ/Unz/hwKO7VbMk0OFa0Sh2sd5m+sp5a
w8uJ8yNh8Y51Q1A6GBMPepnjiKOgabLORCs69zoQXDSr5JxEbI9XaiwtYclplJMK
7lThFmR3hCUUH609+pl07twlg8Mis0sVS85A7rtTG9S/e/vjUBzV0S+3s3knOm6+
jeee3q5/BSyoGjBfJjc0K5ffDeB1uIIAqKh1XhivnmVXY/ayR4P9/QF/2PLsFoBC
PZeqcdEzr29wKo3mwypzxTn+DOnHX4CrhUK/2N3VBuQkWweqRCzRWqVtR+QvclUd
N5G5TuBv48wWhejnzRsIE4saxz6SXkDf4rXY4f/Ailp+jT8VGgRmTXSYggfDJibA
qxQT6G8qxWX+S3eg7BJbxggHfjQluvb0Fp53HuSX0Jd8Ug2IpC/6K/7IrDz8NVnJ
6S9ExE3xrkKfb7xoQOiIOZJWO/BgPh4sLSZ5Z0W+GnB3vK3LfVsmw8Yq6Qn1W9IC
oiWEjkzZiJyS0GB6mMv4Gz9K/9nMmb+GvWBPrjJF7GCZchkMCC304s6G6kX/gX7s
QpqwDYRvvx9v8aXSFrtcdWoZBelR9p4rONHtF+dp1z/Kk1swZcrCS2I16/mRkl8a
YfiGgK+N+mHoUCD7iSA61EREOk9TPaS75ZDyvGCP7FQUZ9wG7WpjiH/qwALO8Ccj
dK0N+ravNGHc7ejaOFhQkyHXRXyPcLfl+asiOac13Uenpgli3NB5CvythGJWc35P
iiomHOErxBT9lqO4LR354fsF4a/0EL77YFIkVgZbQvOLHmIF59SEgID9BX7aMdBl
aAf5yF9zTCT9657zB43vs4HBrAoZwJAcg5+a6ECXnH4c2oOcyCQt1+dHYKfAcGZQ
fMex9VoPPE2I3hVxwggPWPFd2xpDnssdrfVX8edR69sRTjuGYsutpFhRrY7CgAfl
826wrBGmQGkm22Dk+VK7f/UVrjySNjndkvHymG54sP0ARGCb04+0YdowBWa6eR5v
sogS/ixklb+uuBEWFBnm0T359xeOmqITo3+4dh287co2Zw8C6cSkPGD26Wyg5ROA
xBmnpIqjKNGQ3zH6/IVxitv0IiLyLec4iCpQZMXtI7wZGVd0lCjgtBavBYzELMUA
mNSbZVl2LSMtVXwRvHzKYj2D4ueFjDtChCgGRx9k+U1WLbRn5CwNzbl1gaeABLlb
aXsWCnTn9K1zf+VAGCbGWS7U1819c5Lnnub5+J4dbDuDZLhHQlIf64aQKpYqaYKx
oJbiqbZKZXjjR8i/pZIwCg8iJKk9XPnqnM4/zh0gIvddmnRfmZ3nB58rIZPJOTlV
3mklIEBk/o4UsP5s0iOl2BgZNxgcY51JFuTwW2+uJqjwaJJ2iGcQSLwI7lQDVQVj
WfuWzp8bQCJp5e45qiXwbdOSvf0wQ5RyAnZAp5opyj9Ztf4M6Ho4M4gEsX+pWG7i
jNtCru7hjiEa8C6l6lrjWfTOQR26Ago65V2fO8RFhtULLcvAy5Pu2MdJPIVn63gf
3I2puxuU7iFTyNB75iVzsTfhwSyI7vM3QCP2gYXkhDASgFt7mC27q7D+8lxio95v
Vzapz4tAysZFTMb262qvD7XZNhVT6fO8UJJWqpRLeI/8cvfMToTBYHND/xRnN+yD
vf2Rf5O0QTCW8PkhtZ86lHI/TOKa4UkNm4SI2zEDr/hcD/btN3vQFg6wnNyCFRXJ
aRaHDInnwJu/woNBY6oDGCtmgjibQuMTgsMBDnC898VyhZNmP610cN9FcKjo7APk
C/dzfpCnRQqK7hvB1ohQIH035+XU+eWvO8pVrQiVxsEnnR8H/cLDirh6jy+4Q58K
CIKzjkKpdygtNFCXF0yEPQAWrP5M6FjCKK4ft1FymiWKzi72jqg9fGdDv/7e6pc9
HWCGchUJpKrDQuDwZYP90A8Ybgrgy8GmtbK2VoZdPdWPP9u/HegcIaNzniPpkl+a
yrxc6Y0YOgJ4d98IwFkZm8lhyC2B+PY1bveYIowu1Y0Ao/nZMfNzG1P+LXuLjgSq
INIey5PovybjOi/hDfPA3yVoe6v+LCdPtWi5iHelPEsuszZ45LUoRZn2jg6e1wGe
uZ7JvXhOSCwcnZbZwFfyy+pu54VrkZuhqC/BUyRE/IX1qZUUIbxCzCNOjyGqLsqg
iB6vj3BsO+VpE8EuYM0k59FywtldR2Li/qV6wwtEFxjlXLtUpTQjVGl/fva4o4y6
LmkrmaeIJY67A+JZ4wtVm/3uMRVc0osDXmQzQuSofPBo0JvUEC3XqXwtQQXA38dO
tF89Lv5kjXmHIpU2u84809xvVYI5mxE5WiLUFyxtII/hf+ae8KDtmvZSzHv1RhOl
8jB3O6sMAt2ybUvk2qj2XF20+iG3PpkKNTP1degYgatfQXWvwSgciSRtYjl0lX+/
cb7xlxi2XODmK9/1OfkMVAgZWh0c4ZXo5CFO5GyRSD/jmbrb0DrFZJHDLoJyrE0q
zOsFRFfijWIisLBQLVn2pDU7zZYvKF7A9XcNjrfXm0WRUm052jgvCUithh2x/vzX
WXoRVYDiK8Zn/YA6U0NWJ65d5XWpzUhJykEsC34ylIazwPd7nohqoayI56JW10u/
F5a8S+NiPXkEd0HLDZ0XUN4wkxK3Miy9BrLNy5NCDFUWJ+tqZSno8Jg6e60R1W+l
PjXiqZgGQIvKZ0rYTcH1Ze5EjMdZCyoV8fPZChRb13mg/TmZBCwgVe1/n9ejiYZ/
ftZdIBM7f6a/y1TTvT8bOp5+eoTcOZKoc85GSDx3JvYQKGpPbhozrV4kXoomlwv2
4ZNb+KmLEMCfb6un4QLSo85tY02IFmj0453cmO365+f5V/Q01mekgNihZffiUVRO
QusqyOoI0jfq5Y7KGo4QyXmIevPdQ1s7VjEzO6ztBq1kKzeLZJ08sef9O1m+SoGh
3rIqMwLwbKrg/rX6LBSerRISklghdvN0ZRuP38nVC2f189qVM+MEAyng4si+cZYH
R7ek5jpHO7LUg3YVGIKAIseCRY/8XRTHhORKI2NYNip/wUHwbxHRW93c1n/mUicz
/KzS/7y3aOj7oN3c3Hf5dr/BvPx3JDN4cte0bHILuWj93RFxqlMm/Yeavr6wPgVO
3/ijIypA/XLiq4ym96KTsvm/0ODfieNw9BrXDcZ/696u7RF+xsTZHwLhq136kFOD
OEbd1n89XPG5hmfkPQYmcM6ZO2f5b4/gdz6k+s1WeNlw+gqkVhy6cCIulnw+8AWB
CyAI2usuXPNvWmdkXm6rQMkNSKiPf8VFW59M6NCdmJrIKQ4wcqUCJvwy0lslTJD0
CLbW+XdbKWVbqbCr+c44/ZiohgOSaZCW8llghgpiWsasnzQcf4ulpsITOAtzIWZs
MIsuhiNjqoMFAmjhb5KtaVF1SYGneD3Gp5Fz+gE/FHKa+mw8bRFkYXA+NQ8PcQcy
pa+/LgfG3YVXQYv/wEfi7cwVY+wEdOHcslS2x226sig0WP9QUD9AFUeV3hjHIlMT
uVP+WBVA8/5WYK4COnQIaO2fSN5YkGD2oTC02cXv5IoHnGkDUSVJooTG8nPh1Dj8
p+mYz7AAU1kGcJYwmVmw6Vy+AB9XW7MgR8DuxodaTe2MppS1+t1s3wzAQ0+HmYS1
RGJO65qdBiHwGlItRFAYGIDnT64FbS7SmiG9iNKZcFj/8ormlxt3tvrvyqIS23Vp
Mid2fX7U+4szTa+dDCo6wVWrg6sN/rO7lM0SfUkqahG3AZQPwunf/70BtqPrOCAx
xS9LPpwsiHyLJeukep42EeO0MmPZGhSc9Jhv2HTkSICL/TqkpIsptSYvDSp+Oyum
ANncbNUxstXOvy6wKXMUAaok/REoaxDff6/Eq8uq81+rR303a0UnNSFc3nzwofYK
1ZuJquVancxFTFbrkMG1TmhBJHSMIlcXagXVacrG9Kg0LZ4dsnG+j0OYfLi9zMjZ
eDwBoZApoPputKooI2hrtqrcYairp2avr3Bmoa13ZwaTIOsBB3doXatJsUo+jDcM
jSQiBTwaevQBhnq3Z6OzI3FiVnAJLX3OXwpAPa05gJXWcvlDLODmvXqScoPKlPbh
P31HEC5zvVNDo39/Ja39YpGI3w9PVfUA7Ca4Tok1UrAKuKwR/eT9y8S3ovHgM/RO
phobMW+cMzVBqPrQ9LLDbAcv6GqK8xKZ+ofJoJ3opoX3vE0RLEcREJ1m1tjnO98F
qkoa8KDX8XyVMJjflxWDmuGuZW+FyE+4iR/ULli3JF/Uxbx5sAD/RwmHtsxuY2Vl
I5cN37DWW+17R7y4u/jgN9azyZMu558eAsw+ZnA6iRtrMGmmyHzbVKsIHxN7/GxB
1eh/w3lQYSd0jYjSuAd/585a3RCJRbnT8BBLzzj6pryrwd4OewUx6XLUkjP0Mq6j
X1CoiQg+xgrYuDSPtxiVInR/Bcrg7g4GswbATLPorMp+vjPAOL0WB0ONnZ3vcyGk
11JTRaGwRZ6ACa7Z01P9TYdz37d16J5uVHXIwFzNSj5w3kXTwtN2VTh7eS9jnPxG
kZp475v/5HYAFEy2jB8Amr2Wk37Y+06K2rvKrXCHO3ln0E5iEnywGGHatv4d4gPW
xwMEYukoEqlLbBBDFfx9Qzu5piEyImLTZFkGgin3VdqmwmFhjo/qs/0tquhExQdp
XgHgPg6eGG925ESC9ilg1Z/MmRtIfHMSl9eVEp3peJFvznIbeoJ6oaldyRpbP4wK
NL+txNcWZ101DN/phu8cN7CHDpZUHagRavZ/ec/nf6EteuffUaC3ZJevdLYsxcNW
WFLt2Sms8ozD/Jl1WVw5JC8oeS+f7EmtwRjHoH0ckiO29MoM5SPDN3jklPEWgokI
2pY0qvlBEWuSNQ0v7Tete1mdZUdYVxo7GOR6OIAS6TMHKlmqt2iTnmGAHIdIpBKM
6zo8PzgMqc6jesvRn7FfoGff5LtThpQDL0cOwpeYTL6o8kq+O97X6kr+MSKwN2io
/zwA3JWfuhB2r0AoIuktyAQL8QIo0cW8pm1tduNCho0N7tU2zgqwD//xV+6MTzbG
REtDSo7OxO8lA3lqSouZsN0xTE614ucfL52ueWh4XfKdOPsPsBEkwsKDHnTsSg/V
cbAEmn4Aqq5U70APDaqvvgpdVWA+QkZRWw4j/i0CdIROaEYoNQmnUUqEG3gKF+ZG
med9sFUFDZLAFphJtOC+/1za0dmrGMAxI6TI+y+QeHukKOe+mzzDNAkjiF0BfBfz
R/kS/ES2erDLJzmDClkqT3AS1NFc9o/5dxgHi8kRq0K1aNMlEH5jHgth1ANKdsTI
cce3gmAVgA0qsP3m2Soz3KUgYbQQZj83NTRgJZZQom95V91Zbi8N7ggWkkV4q8zs
jB++ZO9XYGNdWj4e5sMiyv/qlOBALAC+WkRv3BN3HWUJ9jdTKcbyayHMxmMyePEg
2T7ZdKEbLTGdDE2XFzcxpW4L6KQ8BX7sYhlVgfCaynMVAlWkkxsvdzgU+myjT1hu
t57h9GCxHImzbe1CORT2OgCATeOa51mYDwpdxXdzzTiHqy2PWgDyHTPHG9jA5OLR
OemBsq7zjfaX2dVe+nK4O9jHVRAM7hbQhINxxjMVsczJYrwEc6RYGXwLmaux65X4
fr4RNWPxwlX0AW8urZ4CD9mjKb5OhKYpMv19mTXZGq6PeIAeI7cx7pwZDUtLC4Nl
qL6Iw5nszlzSF0Bu3xfh1mCChItIIZmZhMhId0Xdi/bWhx2m2jBdu9zDRLPma5LC
7/w/flzZbzDmZb/vA7B4NutIVvTUk5eU8xRVzioQWVLh1KCOn2e/GybwUxAQxEr1
bavUTavhhl23cAmyqMCNEhvrDHiFc7u2nka0PN3MFLcxii22kX/WYM1ZFTulqkLJ
rRRJ3rEy7jtbPEbk8ccOw2Iiy8yzeeAq+1jjefORCHWBBBSTN/9O7NUQy6Bs6OGA
VCleLFwyZvHhU2IpM8ptRQQMGEa8aV2aJ72wsiwyuIV0gqrl+zL2hFL8fXfEz4Jz
q9e7/hdBTZNvwGsB4FWv8+oZEMv1caNsjCVtNIZKlkeL2af40OmApst548685g2P
GZTVJA3ZCs8g14fDtKxzkahbGlWtZBxGNZKNnfJmCUhvYHFtoIakiQlyiUQ3ryEZ
FgU3Mrnos+MVlNyG5oCRC+PWC1suoIyVjGAFYLjXh3/CULtaSN/BMlmndeXlmD3C
YEU5HUTzNpkhqRncyLHwP5M89PyyQSUcBwD6TVGKEL0rZLusfehuue8Qksn8LAT5
d6rbv418JTlfarsVRYzUgQj4NVgJc1gtw0jsvVxs7Q3/TicEEXkNF+n1hkxbo2tA
LzkcHe43KrwWVIMT4oH39jsO69lLOSkY0TLcRYRSgxkwiXkE2OcYaNcdmbnFh80u
fF4I8NKe7ut8knH4x8+5AZqwLkTx+Zoa/lUHCQzog+Pjz6B4LgdEovlRnEchYBk5
r0ZTLTt9BQf4mvZHlWuqXdQv0mLzjneWMLyS/xarihHPB2QrKcqAQNE15GrHNpfG
bZGZlb6JoKXKpqRbUO3NqJLxp5suTBi7UB8PCC0XpbRN+BBQMVojYqvufsoqlOj9
37vST/mvbg6ZsFJCTjpNUOMHewUigjNQsAUQhPZHyEnFiFG20qkx07+dyySCdhdo
VLu0KAXBC1CSX4oxIjwEivR87J8KieAR5Lik/wRI66BA3iSCr6Kc6ObEwA5tIAgc
TKsKHJfpNS/thaQsbrdO5chr/wfeCBbJBubGltNBbxiCFDIv6aKkzTDuChkL7x17
QOXoFCzBNcUZsw3vaXBELuqzTcfoeqjMfCRi5bIAp+zqS7q/1JCeh+2ewx/c1C/B
x+4ux0v3XINqL7Z/MXMrPrsHOP3xKKNzq4lpHBRd6vbggX5kNIIIEz46F6JQtAGO
AbSNk1RIjuXbqZe4nKY3I0WsnJeY0/e5Ky9fEvJySiYmtmRHMcMuPcVeaNQUQN0X
zyM21jx/imKKhNIdDU/+UWgi8T4hpKUlT91IXy3KgPwY/q0s8tImAxodbNeNsU8r
A4TLUy8Oh+lsiruyDCwxmaFAGiJ3UWbPJq0KTyqEPC2qr/4yprZ0cmGMMTS9sVad
eyogPxhcz80oliXYJXVwi1Uuz5JG6MOQ3SkyssVAklF8ftphW6ec7w/YzcUKFBgb
yU4VNCM1n0cbXQ/WsiyYYT4zxAXU6ppltDM7lpGyq4opxN6l4IibVv5IaJlMV1IQ
r1X/h24NsmSaxdYNH6Yf1K9AJfPFuppV/+JbZuUlWmla+kTfx1u26YW+EQx542aq
yIzwYkyVDFXnYQ9nazDPJNZ9RBUQK77kjpRskSmvRa7miBORmyUj38mw1yFpLi7u
C6xoDudDX2yhiBzoeSHZ7K/6UYxzDW8AKVy8hT3VdUmOvt4INibjmYWFDI0RAQV4
+Rp7f3+k/GiZE/nPhl0+K09igZiKfMa5l2HFJIQNA0TCJ6HaGbiijdKc4tel3cZY
Fzs+vHBGll8iUnDgrLJWtv2/mjicCVrdTzj2AkbYsS5NLamccSD7e7Bp1Cjc93Lu
ENNqnmgm2sG9/FXXTrv8aD1oxR9CKURZwSWsSEE9ZSl2tMi/4lqM5iAPBnFVFC2p
JMYtsXeMBhZItHhBieM2YfWQ0llEV5BygoAwz6RMqdLudAJmFR6eH1GUDbB4D4np
wXbK4HZxKhvbcBURqnW3bwhv2EERxlNWlGHl6BF2d0/HgiNMcXuTkMQcy/gBhMGU
+BzplGiZ1lPKXcRwiIe0WJNGrPaujDTxp3DomW996I/u5xNscyueRPLGxFLNzq9z
ceJKI40tmk0m48fiwtIffvzBazlxm1qJTFXrpABl87yFRHuoRI4ELtvZvYQOdL+c
Ej/1kAYSSaFzy7Adqv16OPh2sDir6Ivuya9sbZi1vmqqy0Y+vODSVwDwYYzVOd+Z
DgKfVi3ytTFZyiKGtmRcgji75fTXx7T799TNn4jLZqgMgKPNK3t1B/FbopZxQRSk
75wHSoRfX4xGFLG2ZQoiVumOjR9Co8tjnKgYktLZxIPKWjonrZaD7oF7NZ0T0a8u
SsNL/uzG1PwnTQWeqBWohYEa7m2usU1IDlM7Y8Z9+M2IR+V/SfKqcm1v9YD01jZo
RZJBnDUX7f74jFoAM5s/BWfIo+aQufihpI1xvGS+34moB3U3C111BodsGFi2UNAj
H+S5K0OfXJO2sCvIa+y1t2FbN+NfEThQNZ2yS3ZqvlXj1a/Zs49s8v71yCRUo1W5
12LdMC9zmXZphlKuU4MPGvPtoqG3HQWGQg2xvOjO+yGJGx97yD0ChMzt52pzitJ8
wAwlXghGVWa/yYJtCqGN4YmWZb3wVaLHjLEbI0EAm1BVHTdfELxOlnk2FnzxWorS
q09/2NuCo8V5yAp5BdAp9YLAGmFZDS35JcEWNqUhhOPaGm+nqePDJsQZU4NRKd8k
uyRZro/p5Lkgg68fjZcig7eCpC4VRX+iOmrtq7y2JL4WZcE8+ZdfHtlAb0632tNs
LWYzaU2yFcd2p3bwftlHmDPNTzV3JP4T1EuxXH5Y9P3Su5vVF84wLLB3UzkFbTwT
IXzfyWfEJWHO3imuKRg5wA8lXv71QrllaKetUMi6ocrHvW7hMtOJIxwxa1gNHDTB
9SOYthhKSxX7DHgzPwXDyvqRd4/nWgYEzAsS3eSmjudtTgEyAzAlZLINSOxIzDOJ
tlVt2L4Xy2uvLb9BJKtVJpbSZ/ra4ke2HeDPqx2HgU7/pJXcg8o9pGOSoiiHHQUl
48h1WWjgTl+NSVXJAPtT3yyqHu3SpA4PlYxKNjOEuVRyNN0520i4ezdROCneMVH1
s9bPQn+jpAU1Ho5+Hgp0ReWzS4qrk6ApJvVeTESx9vsb75ysSt5Hn9fnaQS4SDWY
TtgztzV3nxp7e3S7FfFZTu6yhq+3bMtHMwg1Ve9kdhGPzcJPA3qGpCeoe2jVGif6
u6KhHV29zY7ZBOCST99cv/JU39JMUELq8c/ezDusI/znfqprHSXyIYvLXKGu+rKf
ksuUMY/N6+lvL3Yv1vrSCc5qeurIaIqVg2F1qrBguo/oLdbDRQCynyldS8eW3AjE
i3jT9/gVkdEFpK68h9l2rYaWxO+CpCI4W0PLfOrAF8O/zkyQZOMhsjep/4bEAFoM
zHMlJZK1xxC+skLyuEDX5uNP87c7xLmxVGwR6YUZDKYPxXwp96dExD1D/8q/oL1p
c3yqRW/633huIphbIzm5svOu73acu9Bd8m/VxrTb99oAmsoCLwQmgMMzmleuqK9c
AFzGYYcU+qR1ACDgiCG7wpMpo4GmTE1H57WgRXsj7+YuvTF5ix2Iqzae9OGd677F
9o6JreOylJtFPSbJv2xa8+BFEgnefCc5e7AIzgSM+BALTQIZ4w7xc4j2MRzOvXJT
idLaH1p0jo+oaVfjWrogYc0WS0ZqQn/XERMgQdxuzHbu9BGvzn4bPi4B4d0GJqHA
WPK5UDk8ewVJfX6KEiuWUta8nqAyFJ/hdRGY3i8Z1ydvR+j9aXMzLqKbVTTgx7J+
bkvYan+4dRxWTqq4K4z451kEDfwSjrLOEZwtbVc99U9NpoLpZw9uMyo9f9Je60ZO
VpP9A5tk2vou0e5wEYxo/ScNyWTQnIjtH+oAZW1xTKtSIUTK5k+ohEbICATBVJFJ
CSEkFG8dEEq97og19H1Hv8e4acS7/1WbSeFf+U5+l8CLq4tkBpd2DMjPXS0Q5V4+
c86a7Q7mlTuAmRM3OpFAw5CsIfwQe5MLhYguAGZK018=
`pragma protect end_protected
